��   %��A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING���<�PLC�L* ��ST�A� mTRQ_M<��LINK"2&�SX<*Y<*Z/)I�I*IW*Ie$ �R�V* < $� ENBpV_D�EBU��!PN�U;%� UNEVE~ox  �$��ASS  �S���!����� VIRTUAL�/��!' 1 5� ��� ��R?=?v?a?��?�?�?�?�?�?�:�HE M�!8O&O �������]B�   ^��MO �O�?KL�O�O�O�O�O�OzK1_7R _]_o_Z_�_��d�_�_�_�_���=L���_o?�o��@�3oXojo |o�o�o�o5�o�o�o �o#�$�R)SAw62k���� ���#�5�G��"�  M�s���������͏ߏ����'�9��#�$n% 1521D}U%a{����_ ��}_ԟ������� �R�=�v�a������� ͯ��������<�'� `�K�]���������޿ ſϯ�ӿ8�Ͽ\�G� ��kϤϏϡ������� ��"�	��U��|�� �ߋ��߯�������� 	�B�-�f�M�Wߙ�[� ��W��������,�� )�b�M���q������� ������(L7 p[m����� ���!�H�lW �{�����/ �2//#e/'/�/#/ �/�/�/�/�/�/�/.?�?R?=?v?;g�$R5V[�b�8k?�?Nc?  BFo;gx�? O(O:OLO^OpO�O�O�  h 
�  �:  B`�����������S������������@$���\o�����C���@��@r���C� �O__,_>_P_b_t_ �_�_�_�_�_�?�_�_ o(oOLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����o=o2�� V�1oz�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�C�`�G�Y� ��q���̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|σ��χ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ ��(�:�L�^�p����� ���������� $ 6HZl~��� ������2� Bhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??<?N?5?r?M �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_jQ