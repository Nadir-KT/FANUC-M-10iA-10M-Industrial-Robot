��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �SV �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ڏ1�g H PC�UREQ1 � $SOFT; �T_ID�TOT�AL_EQ� $� � NO�PS_�SPI_INDE���$�X�SC�REEN_NAM�E �SI�GN��� P�K_FIL	$�THKYMPAN�E�  	$D�UMMY12 �� u3|4|�R�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"�SBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�:OF�F_ N�3DELHLOGn25Aa2�?i1@N?�(� -M�H W+0�$=Y $DB� 6�COMW!2MO�� 21\D.	 \vrVE�1$F��A{$O��D�B~�CTMP1_F�E2�G1_�3�B�2��XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�08� �zsaC8hq;�G0 � 
$WARNM�0f�!p,P� �s�pNST� �CORN�"a1FL{TR�uTRAT� �T�p H0ACC�a1���{�OR�I
`"S={RT0_�S�B� CHG,I.1 [ Tp�"3I9�TY�D,P*
2 �`w@� �!R*HD�cJ* C��U2��3��4��5��U6��7��8��94����CO�$ <�� $6xK3 1w`O�_M�@�C t e� E#6NGP�ABA� �c��ZQ���`���@nr��� ¸�P�0����x�p�PzPb26�����"J�_R��BCb�J��3�JVP ��tBS��}Aw��"\��P_*0OFSzR; @� RO_K8����aIT�3��NOM�_�0�1ĥ3��T �� $���2AxP��K}EX�� ��0g0I01��p�
$�TFa��C$MD3&��TO�3�0U� ��/ �Hw2�C%1|�EΡg0wE{`vF�vF�40CPp@��a2 
P$A`PqU�3N)#��dR*�AX�!sDET;AI�3BUFV��p@1 |�p۶�pkPIdT� PP[�EMZ�Mg�Ͱj�F[�SIMQSI�"0�ȪA.�����lw 	Tp|zM��P�B��FACTrbHPE�W7�P1Ӡ��u��M]Cd� �$*1�JB�p<�*1DEC�Hښ�H���b� �� +PNS_E;MP��$GP���B,P_��3�p�@Pܤ��TC��|r��0�s ��b�0�� �B���!
����JR� ��SEGKFR��Iv �aR��TkpN&S,�PVF����� & k�Bv�u�cu��aE�� �!2��+�MQ��E�SI!Z�3����T��P������aRSINF �����kq���������LX�����F�C3RCMu�3CClpG� �p���O}���b�1��������2�V�DxIC��C���r����P��L{� EV �zF�_��F�pNB0��?������A�! �r�Rx����V�lp��2��aR�t�,�g�_�RTx @#�5�5"2��uAR��:�`CX�$LG�p���B�1 `s�P�t�aA�0{�У+0R���t�ME�`!BupCrRA 3tAZ�л�pc�OT�FC�b�`�`�FNp���1��ADI+�a%��b�{�@�p$�pSp�c�`S�P���a,QMP6�`Y��3��M'�CUt��aU  $>�TITO1�S�S�!���$�"0�DBPX�WO��!��$�SK��2�@DBd�"�"@�PR8� 
� ���#� >�q1$��)$��+�L9$?(ӤV�%@?R4C&�_?R4ENE��i'~?�A
�!RE�p�Y2(H �O�S��#$L�3$$@3R��;3�MVOks_D@!V�ROScr�r�w�S���CRIG7GER2FPA�S��>7�ETURN0B�c�MR_��TUː\[��0EWM%���cGN>`��RLA���Eݡ�P�&$�P�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWA�YRMO#�aw!�� CS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�g p�QSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc �@Sp�i�a+ �j�f��ΰAPIx2,��$1F�b�$ѐOT�@A� $DUMMAY��Ft��Ft±� |6U- ` !�HE�|s��~bc�B�@ SUFFI���4PCA�Gs5rCw6dr�!MSWU�. 8!�KEYI��5�TM�1�s�qoA&�vINޱ�D, �/ D��HOST�P!4���<���<�0°<��p<�EM'����Z�� SBL� UL>��0  �	�����DT�01� � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0QSp�����#��SAV� ����c�S< 9�`�f�P$�0E!� YN�_B�#2 0�`D�I�d�pO|�m��#�$F�R_IC� �ENC2_Sd3  ��< 3�9���� cgp����!4�"��2�A��ޖ5���`ǻ�@�Q@K&D-!�a�AV�ER�q����DSP
���PC_�q��"��|�ܣ�VALU�3�HE�(�M�I�P)���OPPm ��TH�*��SH" T�/�Fb�;�d�����d D��16� H(rLL_DU ǀ�a�@��k���֠�OT�"U�/��e��R_NOAUT5O70�$}�x�~�@s��|�C ����C� 2iaz�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|�p�����9 <���z�ΓKI����H猡�BaFEq@{@:� ,��&a? �P_P?��>�����E�@��v�QQ���;fp$TP�$VARI����,�7UP2Q`< W�߃TD��g���`������%���BAC�"=# T2����$)�,+r8³�p IFI��p��� q M�P"�r�l@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� Fa@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(��a�#5T�DG���� �%�r�SS� )�? �P(q1�1�`_(1"811�EC1�3D;5D6�GRA����@�����PW��ON2EBU�G�S�2���gϐ_?E A ��@a �TERM�5yB�5 �ORIw��0C�6 �SM�_-`���0D�5����TA�9EIU}P��F� -Q�ϒA�P�3�@B$gSEGGJ� EL�UwUSEPNFI��pBx��1@��4>DC�$UF�P��$���Q�@C���G�0qT�����SNSTj��PATۡg��APTHJ�A�E*�Z%qB�\`F�{E��F�q�pARxxPY�aSHFT͢�qA�AX_SHOR($�>��6 @$GqP9E���OVR���aRZPI@P@$U?r *a�AYLO���j�I��"��Aؠ��ؠERV��Qi�[Y)��G�@@R��i�e��i�R�!=P�uASYM���uFqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P��֊WOR�@M���k0SMT��G��G1R��3�aPA�@�����5�'�H � :j�A�TOCjA7pyP]Pp$OPd�O��C�%�p�O,!��RE.pR�C�A�O�?��Be5pR��EruIx'QG�e$P�WR) IMdu�RR�_$s��5��B I�z2H8�=�_ADD�RH�H_LENG��B�q�q:�x�R��S�o�J.�SS��SK������� ��-�S�E*���rSN�MN1K	�j�5�@r�֣OL��\�WpW�<Q�>pACRO�p�� �@H ����Q� ��OUPW3�b_>�I��!q�a1������ ��|��������-����:���iIOX2S�=�D�e��]����L $��p�!_O�FF[r_�PRM_���aTTP_��H��M (�pOcBJ�"�pG�$H��LE�C��ٰN � 9�*�AB_�T��
�S�`�S��LV��KRW"duH�ITCOU?BGi�LO�q����`d� Fpk�GpSS� ����HWh�wA��O�.��`INCPU>X2VISIO��!���¢.�á<�á-� ��IOLN)�P �87�R'�[p$S�L�bd PUT_&��$dp�Pz ��� F_AS2Q/�$LD���D�aQ"T U�0]P�A���0��PHYG灱Z����4�UO� 3R ` F���H�Yq�Yx�ɱvpP�Sdp���x��\ٶ���UJ��S��v��NE�WJOG�GN �DIS��&�KĠL��3T |��AV���`_�CTR!S^�FgLAGf2&�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_H��Dq��N?���V��EE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�B�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S S�n���_BUFF�1XY��PT�A$�� �v��f�aL6q1YY��P ���\��pOS1�2��3���_�0Z �  ��aiE�*�.�IDX�dP�RhraO�+��A&ST���R��Yz�<! Y$EK&CK+����Z&m&KF�1[ L ��o�0��]PL�6pwq��t^����w��7�_ \ �`��瀰��7��#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3b�DM�R7��LDR5<4R5ORG.���e2 (`���V�8.��T<�4�d^ �q�<4��-4
R5S�`T00m��0D}FRCLMC!D`�?�?3I@��MIC���d_ d���RQzm�q�DSTB	��  �Fg�HAX�;b �H�LEXC#ESZr�rBMup�a`��B;d��rB`�j�`a��F_A�J���$[�O�H0K�db� \��ӂS�$MB既LIБ}SREQUIR�R>q�\Á�XODEBU��oAL� MP�c�ba��P؃ӂ!BoAND���`�`ad�҆�c�cDC1��IN�����`@�(hB?Nz�@q��o��UwPST8� e�r7LOC�RI�p�EX�fA�p��AoA�ODAQP�f Xf��ON��[rMF�� ���f)�"I��%�e���T���FX�@IGG>� g �q��"�E�0��#���$R�a%;#7y��Gx��VvCP�i�DATAw�pE�:�y��RFЭ�NVh t $MD�qIё)�v+�tń�t�H�`�P�u�|��sANSW}��t�?�u�D�)�b�	@Ði[ �@CU��V��T0�eRR2�j �Dɐ�Qނ�Bd$C'ALI�@F�G�s��2�RIN��v�<N��NTE���kE�`��,��b����_N�l��ڂ��kDׄRmn�DIViFDH�@tـn�$V���'c!$��$Z �����~�[���oH �$BE�LTb��!ACCE�L+��ҡ��IR!C�t����T/!��O$PS�@#2L��q�Ɣ83������� ��PATH������"��3̒Vp�A_�Q��.�4�B�Cᐈ�_{MGh�$DDQ�<��G�$FWh��p`��m�����b�DE���PPABNԗROTSPEED����00J�Я8��@����?$USE_��P��s�SY��c�A- kqYNu@Ag���OFF�q�MOUfN�NGg�K�OL�H�INC*��a��q��Bj�L@�BENCS���q�Bđ���D��IN#"I(���4�\Bݠ�VEO�w�Ͳ23_�UPE�߳LOWL����00����D����BwP��� �1RC<ʀƶMOSIV�JR�MO���@GPERoCH  �OV� �^��i�<!�ZD<!��c��d@�P��V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�(�<�p1Ӣ`0 ��RTI$Qx�0 MO���МB R �0J��D��s�H�����b�DUM2(�S�_BCKLSH_C(���>�=�q�#�U���ԑ���2�t�]ACLALvŲ�1n�P�CHK00'%SD�RTY4�k��y�1�q9_6#2�_UM$Pj�9Cw�_�SCL��Ơ�LMT_J1_LDO��@���q��E������๕�幘SP�C��7������PC�o���H� �PU�m�C�/@�"XT_�c�CN�_��N��e���SFu���V�&#����9��(���=�C�u�SH 6#��c����1�Ѩ�o�`0�͑
��_�PAt�&h�_Ps�W�_10��@4�R�01D�VG�J� 1L�@J�OGW����TORQU��ON *�Mٙ�sRHљ��_W��-�_=��C���I��I�I�II�F�`�JLA.�1[�VC��0�D�BO�1U�@i�B\JR�KU��	@DBL�_SMd�BM%`_sDLC�BGRV�`�C��I��H_8� �*COS+\�(LN�7+X>$C� 9)I�9)u*c,)�1Z2 HƺMY@!�(� "TH&-�)THE{T0�NK23I���"=�A CB6CB=�C�A�B(261C��616SBC�T25GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t��Bȿ6���AQ|r�f$N	E�DpIB U�\B5��$!��!A�%E(G8%(!LPH$U�2׵�2SXpCc%pCr%@�2�&�C�J�&!�VAHQV6H3�YLVhJVuKUV�KV�KV�KV�KV�IHAHZF`RXM��TwXuKH�KH�KH�KUH�KH�IO2LOAH�O�YWNOhJOuKO��KO�KO�KO�KO�&F�2#1ic%�d4G�SPBALANC�E_�!�cLEk0H_�%SP��T&�bc&|�br&PFULC�h`r�grr%Ċ1ky��UTO_?�jT13T2Cy��2N&�v� ϰctw�g�p�0Ӓ~����T��O���� I�NSEGv�!�REqV�v!���DIF�f�1l�w�1m
��OB�q
����MI�ϰ1��LCHWA�R����AB&u�$MECH,1� :�,@�U�AX:�P��Y�8G$�8pn 
Z���|���ROBR�CR�(���N��'�M�SK_�`f�p P+ Np_��R����΄ݡ�1��ҰТ΀�ϳ��΀"�IN�q��MTCOM_C|@j�q  L���p��$NORE�³5���$�r �8� GR�E�SD��0ABF�$XY�Z_DA5A���D�EBU�qI��Q�su �`$�COD��G ��k�F�f��$BUFIND�XР  ��MO�R��t $-�U���)��r�B���S�V���Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��E��{�͐OPWOܭŀv0��SY�SBU�@ʐ$SO!P����#�U"��p�PRUN�I�PA��DH�D����_O�U�=��qn�$^}�IMAG��ˀ��0P�qIM����I�N�q���RGOVCRDȡ:���|�P~���Р�0L_6p���Li��RB���0��M���EDѐF� J��N`M*��ื��˱SL�`ŀw x $OVSL�vwSDI��DEXm�@g�e�9w�����V� ~�N���w����Û�4�ȳ�M�]͐�q|<��� x Hˁ�E�F�ATUS����C�0àǒ��BT�M����If���4p����(�ŀy Dˀ!Ez�g���PE�r��p���
���EXE���V��E�Y�$Ժ ŀz3 @ˁ��UP{�h�3$�p��XN����9�H� �PG�"�{ h $S#UB��c�@_��01�\�MPWAI��PL����LO��<�F�p��$RCVFA�IL_C�f�BW�D"�F���DEFS}Pup | Lˀ�`�D�� U�UN!I��S���R`���_L�pP��̐���ā}��� B�~����|��`ҲN�`KET���y���P� $�~z���0SIZE] �ଠ{���S<�OR~��FORMAT/p` � F���rEMR��y�UX������PLI7�ā � $�P_SW�I���͐�_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W R����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�!O�0\H��6@�@�U�� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�Hӱt��W�UpS���R�M��O㵐.'}q��C�g���@ʣ����S�M��AÂ� � $sPY��$WH`'�NGp���H`��Fb`��Fb��Fb��PLM�@��	� 0h�H�{�X��	O��z�Z�eT�M���G� pS��C���O__0_B_�a��_%�� |S����@	 �v��v �@���w�vr��EM��% [R�fr�B�ː��ftPn��PM��QU� �U�Q��Af�wQTH=�HOL��oQHYS�ES�F,�UE��B��O#��  ��P0�|�gAPQ���ʠu���O��ŀ�ɂv�-�A;ӝGROG��a2D��E�Âv�_�ĀZ�INFO&��+����b�Ȝ�OI킍 ((@SLEQ/�#@������o���S`�c0O�0�01E�Z0NUe�_�AUT<�Ab�COPY���(��{��@M��N������1�P�
� ��RG4I�����X_�Pl�C$�����`�W���P��j@�G���E�XT_CYCtb����p����h�_NA�!$�\�<��RO�`]�� �s m��POR�㸅����SRVt�)l����DI �T_l� ��Ѥ{�ۧ��ۧ �ۧU5٩6٩7٩8��҆AS�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,(@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#q�RQSK;IP�� ĕ�x�-O�`NT!� ��P_x���ǚ@�b�p 1�1�1Ǹ�?� � ?��>��>�&�>�3�z>�9�J2R;n쐖 4��EX� TQ����ށ�Q����[�KFд��@RDCNIf� �U`�X}�R�#%M!*�0�)��$�RGEAR_0I9O�TJBFLG�i&gpERa��TC݃��|����2TH2N���� 1�b��G:q T�0 ����IM���`Ib��w��REF�1�� yl�h��ENAB��lcTPE?@���! (ᭀ����Q�#�~��+2 H�W���2�Қ����"�4�F�X�j�3�қ{��������
j�4�Ҝ��
��.�(@�R�j�5�ҝu������������j�6�Ҟ���(:Lj�7�ҟo�����
j�8�Ҡ��"x4Fj�SMSK������a��E�A~�QREMOTE������@ "1��Q&�IO�5"%I��P���POWi@쐣  �����X�gpi��쐤��Y"$DSB_SIGN4A�Qi��̰C���tRS23�2%�Sb�iDEVICEUS#�R�R�PARIT�!O�PBIT�Q��O?WCONTR��QXⱓ�RCU� M�S�UXTASK�3NxB��0�$TATU�PK��S@@쐦F��6�_�PC}�$F�REEFROMS8]p�ai�GETN@S��UPDl�ARB�S�P%0���� !>m$USA���a8z9�L�ERI�0f�&�pRY�5~"_�@f�qP�1�!�6WRK�D9�F9ХFR�IEND�Q4bUFx��&�A@TOOLHF�MY5�$LEN�GTH_VT��FCIR�pqC�@�E� �IUFIN�R����RGI�1�AITI:�xGX��I�FG2�7G1a����3��B�GPRR�DA��Oa_� o0e�I1RER�0đ�3&���TC���AQJV �G|�.2���F��1�!d�9Z�8 +5K�+5��E�y�L0�4��X �0m�L
N�T�3Hz��89��%��4�3G��W�0�W�RdD�Z��Tܳ���K�a3d��$cV �2���1��I1TH�02K2sk3K3Jci�aI�i�a�0L��SL��R$Vؠ�B�V�EVk�]V*R��� �,6Lc���9V2�F{/P:B��PS_�E���$rr�C�ѳ3$A0��wPR���v�U�cSk�� {��8��G� 0���VX`�!�tX`��0P�Ё��
�5SK!� �"-qR��!0���z�MNJ AX�!h�A�@�LlA��A�THIC��1�������1TF�E���q>�IF_C	H�3A�I0�����G1�x������9��Ɇ_JF҇PR|(���RVAT�� �-p��7@�����DO�E��COU�(��AXIg��O�FFSE+�TRIG�SK��c���Ѽ�e��[�K�Hk���8�IG#MAo0�A-��ҙ��ORG_UNEV���� �S�쐮�d �$�������GROU��ݓTqO2��!ݓDSP���JOG'��#	�_P'�2OR���>P67KEPl�IR�0�2PM�RQ�AP�Q���E�0q�e���SYS�G��"��PG��BRAK*Rd�r�3�-���0����ߒ<pAD�ݓ�J�BSOC� N��DUMMY14��p\@SV�PDE_�OP3SFSPD�_OVR��ٰC�O��"�OR-��Nı0.�Fr�.��OV��SFc�2�f��F���!4�S��RA�"L�CHDL�REC�OV��0�W�@M�յ�RO3��9_�0� @�ҹ@�VERE�$OF�S�@CV� 0BWD�G�ѴC��2j�
�T�R�!��E_F�DOj�MB_CM4��U�B �BL=r0�w�=q�tVfQ��x0spd��_�Gxǋ�AM��`k�J0������_M���2{�#�8$CA��{Й���8$HB�K|1c��IO��8.�:!aPPA"�N��3�^�F���:"�DVC_DB�C��d�w"����!��1���ç�y3����ATIO� �q0�UC�&CAB�BS�PⳐ�P�Ȗ��_0c�S�UBCPUq��S �Pa aá�}0�Sb��c���r"ơ$HW_AC���:c��IcA�A~-�l$UNIT��l��ATN�f�����CYCLųNEC�A��[�FLTR_2_FI���(��}&Ɩ�LP&�����_S[CT@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb��r�: _T��PROX��O�� EM�_�r��8u�q u��q��DI�0e�RAOILAC��}RMƐCLOԠdC��:anq���wq����PR��S�LQkfC�ѷ 	���FUNCŢ�rRINkP+a�0 ��!3RA� >R 
Я8�ԯWAR�#BLFQ��A�����DA�����LDm0�aB9�2�nqBTIvrb8ؑ���PRIAQ1�"AFS�P�!���𰠓�`%b���M�I1U�DF_j@��y1�°LME�FA�@H�RDY�4��Pn@R�S@Q�0"�MUL�SEj@f�b�q ��X��ȑ���m$.A$�1$c1�Ó���� x~�EGvpݓ�q!cAR����09>B��%��AXE��RKOB��W�A4�_�-�֣SY���!6��&S&�'WR���-1����STR��5�9�E�� 	5B��=Q�B90�@6������O�T�0o 	$�A�RY8�w20���	�%�FI��;�$LGINK�H��1�aI_63�5�q�2XYZ"��;�q�3@�R�1�2�8{0B�{D��� CFI��6G��
�{��_J��6��3aO�P_O4Y;5�QT�BmA"�BC
�z�D�U"�66CTURN3�vr�E�1�9���GFL�`���~ �@��5<:7�� 1��?0K�Mc�68�Cb�vrb�4�ORQ ��X�>8�#op�������wq�Uf�����TOVE�Q��M;�E# �UK#�UQ"�VW�ZQ �W���Tυ� ;��� �QH�!`�ҽ��U�Q�W`keK#kecXER�
�	GE	0��S�dAWaǢ:D���7!�!AX�rB!{q ��1uy-!y�p z�@z�@z6Pz\P z� z1v�y� y�+y�;y�Ky� [y�ky�{y��y�qޜyDEBU��$ ����L�!º2WG` � AB!�,��SV���� 
w���m� ��w����1���1���A ���A��6Q��\Q���!��m@��2CLAB�3B�U�����S 7 ÐER����� � $�@� A6ؑ!p�PO���Z�q0w�^�_MRA�ȑ� d  T�-�ERR��STYz�B�I�V3@��cΑTOQ�d:`L � �d2ᕴP��˰[!_ � p�`T}0i��_V1�r�a'�4�2-�2<�����@P�����F�$W���g��V_!�l�$�P����c��q"��	�SFZN_wCFG_!� 4�� ?º�|�ų����@�Ȳ�W W]���\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(�����!�s�Q�g�P{RV H�ELLĥ� }56�B_BAS!�GRSR��ԣo �#QS��[��1r�%��U2ݺ3ݺ4ݺ5ݺ�6ݺ7ݺ8ݷ��R�OOI䰝0�0NL�K!�CAB� ��A[CK��IN��T:��1�@�@ z�m�_P�U!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KcARӑ�@��RE~���P��(��QUE������P
��CST?OPI_AL������0&���㰑�0SE�Ml�b�|�M��d�T�Y|�SOK�}�DI������(���_T}M\�MANRQ���0E+�|�$KEYSWITCH&�	���HE
�BE�AT����E� LE(Ғ���U��FO���|��O_HOM��O�REF�PPR�z��!&0��C+�OA�ECO��B�rIOCM�D8׵��]���8�` � �D�1����U��&�M�H�»P�CFORC<��� �'�����OM�  � @�V��|�U,3P� 1(-�`� 3-�4���NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F��V ��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7s�VP�U�PD��  ���|�԰��YSLO>Ǣ� � z��� ����o�E��`>�^t���АALUץ����C�U���wFOqID_YL�ӿuHI�zI�?$FILE_���tf��$`�JvSA���� h���E_B�LCK�#�C,�D_CPU<�{�<�o�����tJr��R ;��
PW O�[ ��LA��S��8������RUNF�Ɂ ��Ɂ����F�ꁡ�ꁾ�� �TBCu�C�� �X -$�LENi��v������I��G�LOWo_AXI�F1�
�t2X�M����D�
 ���I�� ��}�T#OR����Dh��� L=��⇒�s���#�_MA`�ޕ���ޑTCV����T ���&��ݡ����J�$����J����Mo����J�Ǜ �������2��� v�����F�JK��VKi�ΡvњΡ3��J0�ңJ�JڣJJ�AAL�ң�ڣ��4�5z�&�N1-�9����J��L~�_Vj�Z����� ` �GGROU�pD��B�NFLIC��R�EQUIREa�E�BUA��p����2�¯�����c��� \��APPR���C���
�EN��CLOe��S_!M v�,ɣ�
���o� ��MC�8&���g�_MG�q��C� �{�9���|�B;RKz�NOL��|�:� R��_LI|���$��k�J����P
��� ڣ�����&���/���Q6��6��8��r�>��� ��8��%�W�2�e�PATHa�z�p�z�=�vӥ��ϰ�x�CN=�CA������p�IN�U�C��bq��CO�UMB��YZ������qE%����2������PAYwLOA��J2L3pOR_AN��<�L���F�B�6�R�{�R_F�2LSHR��|�L�OG��р��ӎ���ACRL_u��������.���H�p�$H�{���FLEX
���J�� : �/����6�2�����;�M�_�F16�����n���������ȟ��E ҟ�����,�>�P� b���d�{������ ������5�T��X��v���Eťm Fѯ�������@&�/�A�S�e�D�Jx�� � �������j�4pAT����n�EML  �%øJ����ʰJE��CTR,�Ѭ�TN��F&��HAND_VB[q
�pK�� $�F2{�6� �rSW�i�D�U��� '$$Mt�h�R��08@��@<b 35��^6A�p 3�k��q{9t�A�̈p
��A��A�ˆ0��U����D��D��P��G��IST��$A��$AN��DYˀ�{�g4 �5D���v�6�v��5� ���^�@��P��� ��#�,�5�>�+p�K�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������$uN���
D�찙H������"CqE�N� a�DI��>�OpbtC�Dpx�� �
�2IxQA�q��q���-��s �� �����{ ��OMME���rr/�TVpP�T�P ���qe�i� ���P�x ��yT�Pj�� $DUMM�Y9�$PS_6��RFq�  ��:�� ���!~q�c X����K�STs��ʰSBR��M2�1_Vt�8$SV_ERt�O��z���WCLRx�A  O�r�?p? Oր � �D $GLOB���#LO��Յ$�po��P�!SYS�ADR�!?p�pTC}HM0 � ,�����W_NA���/�e�$%SR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T>D�XSCRE�ƀ5�� ��STF���#}�pТ6�C�] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��uD�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRI# �m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$���VSHI9F��|s�P�p��6�s���R���OS�URW�pRADIz��2�_�q�h�`g! �q)�LUza�$OUTPUTg_BM��IML��oR6(`)�@TILN<SCO�@Ce� ;��9��F��T�� a��o�>�3���$��w�2u�<qV�zu9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+��t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2$��2���5��`�? ��ZAB�CS��  $��2��J�
���$$�CLAS������AB���'@@V�IRT��O.@AB�S�$�1 <E�� < *AtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v�����M@[�AXLր`�&A��dC  ���IN8��ā��PRE������LARM�RECOV �<I䂥�NG�� �\K	 =#�
�J�\�M@PPLIC��?<E�E��HandlingTool ��� 
V7.50�P/28 *A��b��
�_S�W�� UP*A�� ��F0ڑ����A����� 20���*A���:�����m(B �7DA5�� �~'@	b@�𞝓None������� ��Tg}�*A4�`x��P_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ�:�i�n�����#B)B ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��&��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���o&�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� ��PB�Z?����5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`ϖ�S:�(����Yp0�_)o�S`�BBia�P�_mo8j�(�aKoo�o9i�(Ѕ�og�o�o�oLnf��oGq:I�ZDEFg f8��)�R�6pbuf.txt m�]n�@����# �	`(Ж�A=L�m��zMC�21�=���9���4�=��n׾�Cz  BH�BCCPUeB���CF�;.�<C���C5�rSZE@D�nyD�Q��D��>���D�;D�����F��>�F�$G}RB�Gzր���SY��!�vqGR���Em�(�.��(�(��<�q�G�Sx2��Ң �� &a�D�j���E�e���EX�EQ��EJP F�E��F� G��ǎ^F E�� �FB� H,- �Ge��H3Y����  >�33� ���xV  in2xQ@��5Y���8B� A�AST<#�
� �_'�%��w�RSMOFS��،~2�yT1�0DE' �O c
�(�;;�"�  <�6��z�R���?�j�C�4��SZm� W�(�{�m�C��B-G��C�`@$�q��T�{�FPROG !%i����c�I��� ��Ɯ�f�KEY_TOBL  �vM�u�� �	
��� !"#$%&'�()*+,-./�01c�:;<=>�?@ABC�pGH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������p���͓���������������������������������耇����������������������!j�LCK�.�j���STAT����_AUTO_�DO���W/�IN?DT_ENB߿21R��9�+�T2w�X�STOP\߿2TR�Ll�LETE�����_SCREEN� ikc�sc��U��MME�NU 1 i  <g\��L�SU +�U��p3g����� ��������2�	��A� z�Q�c����������� ����.d;M �q����� �N%7]�m ���/��/ J/!/3/�/W/i/�/�/ �/�/�/�/�/4??? j?A?S?y?�?�?�?�? �?�?O�?O-OfO=O OO�OsO�O�O�O�O�O�_�O_P_Sy�_M�ANUAL��n�DwBCOU�RIG��>�DBNUM�p���<���
�QPXW�ORK 1!R� ү�_oO.o@oRk�Q__AWAY�S��/GCP ��=��df�_AL�P�db�RYв������X_�p 1}"�� , 
�^@���o xvf`MT��I^�rl@�:sON�TIM�����ɼZv�i
õ�cMO�TNEND���dR�ECORD 1(�R�a��ua�O� �q��sb�.�@�R� �xZ�������ɏۏ 폄���#���G���k� }�����<�ş4��X� ��1�C���g�֟�� ������ӯ�T�	�x� -���Q�c�u������� ���>����)Ϙ� Mϼ�F�࿕ϧϹ��� :�������%�s`Pn&� ]�o��ϓ�~ߌ���8� J�����5� ��k� ���ߡ��J�����X� �|��C�U������ ����0�����	���dbTOLEREN�CqdBȺb`L��͐PCS_CFG� )�k)wd�MC:\O L%0?4d.CSV
�P�c�)sA �CH
� z�P)~����hMRC_OUT *�[�`+P ?SGN +�e�r���#�10-M�AY-20 10�:38*V27-J{ANj21:4r�v P;����)~�`pa��m��PJP�ѬVERSI�ON S�V2.0.�6tE�FLOGIC 1�,�[ 	DX��P7)�PF."PROG_ENB�o�rj ULSew �T�"_WRSTJNEp��V�r`dEMO_O�PT_SL ?	��es
 	R575)s7)�/??�*?<?'�$TO  a�-��?&V_@p�EX�Wd�u�3P�ATH ASA�\�?�?O/{IC�T�aFo`-�g|dsegM%�&ASTBF_TTS�x�Y^C��SqqF�PMAU� t/Xr�MSWR.�i6(.|S/�Z!D_N �O0__T_C_x_g_�_��tSBL_FAU�L"0�[3wTDI�AU 16M6p���A1234567890gFP?BoTofoxo�o�o �o�o�o�o�o,�>Pb�S�pP�_ ���_s�� 0` �����)�;�M� _�q���������ˏݏ8��|)UMP�!�3 �^�TR�B�#�+�=�PMEfEI�Y�_TEMP9 ÈÓ3@�3A v�UN�I�.(YN_BR�K 2Y)EMGDI_STA�%�WЕNC2_SC/R 3��1o"� 4�F�X�fv�������0��#��ޑ14�����)�;�����ݤ5�����x�f	 u�ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/߭P� b�t�� ��xߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N���r� �������������� &8J\n�� ������" `�FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/4?,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O?�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�O�O �o�o�o
.@R dv������ ���*�<�N�`�r� ���o����̏ޏ��� �&�8�J�\�n����� ����ȟڟ����H��ETMODE 1�6��� 
��ƨ
R�d�v�נ�RROR_PROoG %A�%�:����  ��TABL/E  A�������#�L�RRSEV_NUM  ��Q��K�S����_AUTO_EN�B  ��I�Ϥ_;NOh� 7A�{�}R�  *�������������^�+રĿֿ迄�HIS�O�͡I�}�_ALMw 18A� �;�����+�e�w� �ϛϭϿ��_H���  A���|���4�TCP_VER� !A�!����$�EXTLOG_R�EQ��{�V�S�IZ_�Q�TOL � ͡Dz���=#׍�XT_B�WD����r���n�_�DI�� 9���}�z�͡m���ST�EP����4��OP�_DO���ѠF�ACTORY_T�UN�dG�EAT?URE :�����l�Han�dlingToo�l ��  - C�Englis�h Dictio�nary��ORD�EAA Vi�s�� Masteyr���96 H���nalog I/yO���H551���uto Soft�ware Upd_ate  ��J���matic Ba�ckup��Par�t&�ground Edit���  8\ap�Camera��F���t\j6R�elyl���LOADR�7omm��shq��oTI" ��co��
! o���p�ane�� 
!���tyle s�elect��H5�9��nD���oni7tor��48�����tr��Relia�b���adin�Diagnos�"����2�2 ual� Check S�afety UI�F lg\a��h�anced Ro�b Serv q� ct\��lUs�er FrU��D�IF��Ext. oDIO ��fiAs d��endr �Err L@��I%F�r��  �П��90��FCTN /MenuZ v'���74� TP In���fac  S�U (G=�p���k Excn g��3��High-wSper Ski+�  sO�H9 � m�munic!�on5sg�teur� �����V����c�onn��2��ENމ�Incrst�ru���5.fd�KAREL �Cmd. L?u�aA� O�Runw-Ti� Env��R��K� ��+%�s#�S/W��74��L?icenseT��  (Au* ogBook(Sy���m)��"
MACROs,V�/Offse��a�p��MH� ����p�fa5�MechS�top ProtL��� d�b i��Shif���j545�!xr ��#���,pb ode Switch��m\e�!o4.�& pro�4���g��Multi�-T7G��net�.Pos RGegi��z�P���t Fun���3s Rz1��Numx ������9m�1�  �Adjuj��1 J7�7�* ����6�tatuq1EIK�RDMtot���scove�� ���@By- }uest1�$Go� � U5�\SNPX �b"���YA�"Li�br����#�� �$~@h�pd]0�J�ts in VCCCM�����0�  �u!��2 R�0�/�I�08��TMI�LIB�M J92:�@P�Acc>�F�{97�TPTX�+6�BRSQelZ0�M�8 Rm��q%��6�92��Unexc�eptr motn>T  CVV�P���KC����+-��~K  II)�VS�P CSXC�&.ac�� e�"�� t�@�Wew�AD� Q�8bvr nm�en�@�iP� a�0y�0�pfGri�dAplay !�� nh�@*�3R�1M-�10iA(B20k1 �`2V"  F����scii�lo{ad��83 M��yl����Guar�dO J85�0�mP'��L`���stuaPa9t�&]$Cyc����|0ori_ x%Da�ta'Pqu���cAh�1��g`� j� RLJam�5���IMI De-B(�\A�cP" #^0C~  etkc^0�asswo%q�)6�50�ApU�Xn�t��Pven�CT�qH�5�0YELLOW BO?Y���� Arc�0vi�s��Ch�Wel=dQcial4Izt�Op� ��gs�`k 2@�a��poG3 yRjT1 NEf�#HT� xyWbF��! �p�`gd`����p\� =P��JP�N ARCP*P�R�A�� OL��pSup̂fil��p��J�� ��cro�670�1C~E�d���SS�pe�tex��$ �P� So7 t^� ssagN5 <Q"�BP:� �9 "0�Q#rtQC��P�l0dpn�笔�rpf�q��e�ppmas�cbin4psy=n�' ptx]08��HELNCL �VIS PKGS9 �Z@MB &���B J8@IPE� GET_VAR� FI?S (Un�i� LU�OOL:� ADD�@29.KFD�TCm���E�@�DVp���`A�ТN�O WTWTEST �� �!��c��FOR ��ECT� �a!� ALSE� ALA`�CPMO-130��� b �D: HANG FROMg��2���R709 DRA�M AVAILC�HECKS 54�9��m�VPCS �SU֐LIMCH�K��P�0x�FF WPOS� F�� q�8-12 C�HARS�ER6�O�GRA ��Z@AV�EH�AME��.SV��Вאn$��9�wm "y�TRCv�� SHADP�UP�DAT k�0��S�TATI��� M�UCH ���TI�MQ MOTN-�003��@OB�OGUIDE DAUGH���b��@�$tou� �@C� <�0��PATH�_��MOVET�� R�64��VMXPA�CK MAY A�SSERTjS��C�YCL`�TA��B�E COR 71��1-�AN��RC �OPTIONS � �`��APSH-�1�`fix��2�S�O��B��XO򝡞�_�T��	�i��0j��d�u�byz p wa��y�٠HI�������U�pb XSPD �TB/�F� \hcehΤB0���END�[CE�06\Q�p{ }smay n@��pk��L ��tr'aff#�	� ���~1from sy�svar scr��0R� ��d�DJUD���H�!A��/��SET ERR��D�P7����NDA�NT SCREE�N UNREA �VM �PD�D��P�A���R�IO gJNN�0�FI��}B��GROUNנD Y�Т٠�h�SVIP 53 Q�S��DIGIT �VERS��ká�N{EW�� P06�@=C�1IMAG�ͱ4���8� DI`����pSSUE�5��EPLAN JON�� DEL���157�QאD��CALL�I���Q��m���IP�ND}�IMG N�9 PZ�19��MwNT/��ES ���`LocR Hol�߀=��2�Pn� PG�:��=�M��can�����С: 3D� mE2view gd X��ea1 ��0b�pof Ǡ"�HCɰ�ANNO�T ACCESS? M cpie$E�t.Qs a� lo^MdFlex)a:���w$qmo G�sA�9�-'p~0��h0pa���eJ AUTO1-�0��!ipu@Т|<ᡠIABLE+�� 7�a FPLN:9 L�pl m� �MD<�VI�и�W�IT HOC�Jo~1Qui��"���N��USB�@�Pt� & remov����D�vAxis �FT_7�PGɰC�P:�OS-14�4 � h s 2968QՐOST�p � CRASH D�U��$P��WOR�D.$�LOGI�N�P��P:	�0�0�46 issue�E�H�: Slo[w st�c�`�6����໰IF�I�MPR��SPOT�:Wh4���N1STyY��0VMGR�\b�N�CAT��4oR�RE�� � 5�8�1��:%�RTU�!Pe -M a�SE:B�@pp���AGpL��r�m@all���*0a�OCB WA����"3 CNT0� T9DWroO0a�larm�ˀm0d� t�M�"0�2|� 9o�Z@OME<�� ���E%  #1-�S�RE��M�st}0g�     5K�ANJI5no �MNS@�INISITALIZ'�3 E�f�we��6@�� dr�@ fp �"��SCII L��afails w|��SYSTE[��i��  � Mq��1QGro8�m �n�@vA����&��nx�0q��RWRI �OF Lk��� \gref"�
�up� de-rela�Q_d 03.�0SS�chőbetwe�4�IND ex 6ɰTPa�DO� �l� �ɰGigE��soperabi]l`p l,��Hc�B��@]�le�Q0c�flxz�Ð���O�S {����v4pfigi GLA�$�c2z�7H� lap�0�ASB� If��g�2 l\c�0��/�E�� EXCE	 㰁�P���i��� o0��Gd`]Ц�f<q�l lxt��EFal��#0�i�O�Y�n�CLOS��S[RNq1NT^�F��U��FqKP�ANIO' V7/ॠ1�{����DB �0���v��ED��DET|��'� �bF�NLI;NEb�BUG�T�:��C"RLIB��A���ABC JAR�KY@��� rkeMy�`IL���PR���N��ITGAR� D$�R �Er *�T��a�U�0��h�[��ZE V� TASK p.vr��P2" .�XfJ�srqn�S谥dIBP	c����B/��BUS.��UNN� j0-��{��cR'���LO�E�DIVS�CUL`s$cb����BW!���R~�W`P�����I�T(঱tʠ�OF��UNEXڠ+����p�FtE��SVE�MG3`NML 5�05� D*�CC_SAFE�P*� ���� PET��'P�`��F  !���IR(����c i S>� �K��K�H GU�NCHG��S�M�ECH��M��T�*�%p6u��tPOR�Y LEAK�J���SPEgD��2�V 74\GRI���Q�g��CTLN��TRe @�_�p ��6�EN'�IN���`���$���r��T3)�.i�STO�A�s�	L��͐X	���q��1Y� ��TO2�J �m��0F<�K����D)U�S��O��3	 9�J F�&���S?SVGN-1#I�N��RSRwQDAU�C@ޱ� �T6�g��� 3��]���BRKCTR8/"� �q\j5��_��Q�S�qINVJ0D ZO�Pݲ���s���г�Ui ɰ̒�a�D�UAL� J50�e�x�RVO117 AW�TH!Hr%�nN�247%�52��|�&aol ���R��(�at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���M�d�Rǰt� \fosB�A�0Np�c�����{�U��ROP �2�b�pB��ITP�4M��b !AU�t c0< � plet9e�N@� z1^q�R635 (Ac�cuCal2kA���I) "�ǰ�1
a\�Ps��ǐ� b���0P򶲊���ig�\cbacul "A3p_ �1��ն����etaca��AT���PC�`�����;_p�.pc!Ɗ�<�:�circB����5�tl��Bɵ�:�f!m+�Ί�V�b�ɦ�~r�upfrm.����ⴊ�xed��Ί�N~�pedA�D �}b>�ptlibB�� �_�rt��	Ċ�a_\׊ۊ�6�fm�� ��oޢ�e��̆Ϙ���c�Ӳ�5�j>�����#tcȐ��	�r���ʸ�mm 1��T�sl�^0��T�mѡ�#�r�m3��ub Y�q�s3td}��pl;�&�cckv�=�r�vf������9�vi����Cul�`�0fp�q ��.f��� daq�; i Data A�cquisi��nB�
��T`��1��89��22 D�MCM RRS2�Z�75��9 3 �R710�o59�p5\?��T "��1 (D�T� nk@��������E Ƒ�ȵ��Ӹ�etdm�m ��ER����gxE��1�q\mo? ۳�=(G���[0(

�2�` ! �@�JMACRO��S�kip/Offs�e:�a��V�4o9<� &qR662����s�H�
 6Bq8�����9Z�43 �J77� 6�J783�o ��n�"vv�R5IKCBq?2 PTLC�Z�g R�3 (�s�, �������0�3�	зJԷ\sf�mnmc "MN�MC����ҹ�%mnf�FMC"Ѻ0�>� etmcr� ��8���� ,�pDp �  874\p'rdq>,jF0�ޢ�axisHPr�ocess Axwes e�rol^�PRA
�Dp� 56o J81j�59� 56o6� ���0w��690 98� [!I#DV�1��2(x2��2ont�0�
�����m2���?C��e�tis "ISD���9�� Fprax�RAM�P� D��d�efB�,�G�is_basicHB�@p޲{6�� 708�6��(�Acw:�������D
�/,��AMOX �� ��DvE��?;T��2>Pi� RAFM';�]�!PAM�V�W�Ee`�U�Q'
bU�75��.�ceNe� nt?erface^�1' 5&!54�K��b(Devam±�/�#����/<�Tane`"�DNEWE���btp_dnui �AI�_�s2�d_rsono���bAsfjN��bdv_arFvf�x0hpz�}w��hkH9x�stc��gApon1lGzv{�ff� �r���z�3{q'�Td>pchamp�r;e�p� ^597@7��	܀�4}0��mɁ��/�����lf�!�pcochmp]aMP&xB�� �mpev��8����pcs��Ye�S�� Macro�OD��16Q!)*��:$�2U"_,��Y�(PC ��$_;�������o��J�gegemQ@GEMSW�~ZG�gesndy��OD��ndda��S��s1yT�Kɓ�su^Ҋ�ĩ�n�m���L��  ���9:p'ѳ޲���spotplusp���`-�W�l�J��s��t[�׷p�key�ɰ�$��s�-Ѩ��m���\featu� 0FEAWD�o;olo�srn'!�2 p���a�As3��t�T.� (N. A.)��!e!�J#
 (j�,��oBIB��oD -�.�n��k9�"K��u[-�_����p� "PSE�qW����wop "sEЅ�&�:�J��� ���y�|��O8��5� �Rɺ���ɰ[��X� ������%�(
ҭ�q HL�0k�
�z�@a!�B�Q�"(g� Q�����]�'�.��� ��&���<�!ҝ_�#��tpJ�H�~Z��j��� ��y������2��e� �����Z����V��! %���=�]�͂��^2�@�iRV� on�Q$Yq͋JF0� 8ހ�`�	(^�dQueue���X\1�ʖ`�+~F1tpvtsn��YN&��ftpJ0v �RDV�	f��J1 iQ���v�en�^�kvstk��mp���btkclrq8���get�����r��`kacqk�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�m	c�N+v3�_� �����.v�/\jF��� �`Q�΋�ܒ�N50 (FR�A��+��͢fraparm��Ҁ�} =6�J643p:V��ELSE
#�V�AR $SGSY�SCFG.$�`_UNITS 2�D`G~°@�4Jgfr��4A�@FRL-��0ͅ �3ې���L�0NE�: �=�?@�8�v�9~Q�x304��;�BPR�SM~QA�5TX.�$VNUM_OLp��5��DJ507��~l� Functʂ�"qwAP��琉�3 �H�ƞ�kP9jQ�Q5 ձ� ��@jLJzBJ[ �6N�kAP����S>��"TPPR��\�QA�prnaSV��ZS��AS8Dj510U�-�`cr�`8 ���ʇ�DJR`jYȑH_  �Q �P�J6�a21��48�AAVM 5̕Q�b0 lB�`TU�P xbJ54s5 `b�`616����0VCAM ~9�CLIO b71�5 ���`gMSC8�
rP R`�\sSTYL� MNIN�`J6�28Q  �`NR�Ed�;@�`SCH ���9pDCSU M�ete�`ORSR� Ԃ�a04 kR�EIOC �a5.�`542�b9vpP@<�nP�a�`�R�`7�`��MASK 3Ho�.r7 �2�`OOCO :��r3� �p�b�p���r0X��a��`13\mn�a3?9 HRM"�q�q~��LCHK�u�OPLG B��a0�3 �q.�pHCR� Ob�pCpPosyi�`fP6 is[r�J554�òpDS�W�bM�D�pqR�a337 }Rjr0 �1�s�4 �R6�7��52�r5 �2�r7 1� P6���Regi��@T�uFRD�M�uSaq%�4�`9{30�uSNBA�u�SHLB̀\sf�"pM�NPI�S�PVC�J520v��TC�`"MNрoTMIL�IFV��PAC W�pTP�TXp6.%�TELN N Me��09m3UEC9K�b�`UFR�`���VCOR��VIPuLpq89qSXC�S��`VVF�J�TPy �q��R626l��u S�`Gސ�2�IGUI�C��P�GSt�\ŀH86�3�S�q�����q34:sŁ684���a��@b>�3 :B��1� T��96 .�+�E�51 y�q53̀3�b1 ���b1 �n�jr9 ���`VAsT ߲�q75 s�xF��`�sAWSMӞ�`TOP u�ŀRq52p���a80 
��ށXY q���0 \,b�`885�QXр�OLp}�"pE࠱t�p�`LCMD��EgTSS���6 �>V�CPE oZ1�gVRCd3
�NLH�h��001m2Ep���3 f��p��4 //165C��6l����7PR��008 �tB��9 -200��`U0�pF�1޲1	 ��޲2L"���p���޲4��5 \h�mp޲6 RBCF`�`ళ�fs�8 ������~�J�7 rbcfA�L�8\PC����"�32m0u�n�K��Rٰn�5 5EW�
n�9 z��4�0 kB��3 ��6|ݲ�`00iB/��I6�u��7�u��8 �0�������sU0�`�t� �1 05\rb��2 E���K���dj���5˰��60��a�HУ`:�63�jAF�_���F�7 ڱ݀H�a8�eHЋ��cU0���7�p��1u��8<u��9 73����&��D7� ��5t�W97 ��8U�1���2��1�1:���h���1np�"��8(�U=1��\pyl��,�p��v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6C B���цp��1��r��1�`͵155ض�157 �2��62 �S����1b��2$����1Π"�2����B6`�1<c�4� 7B�5 DR��8�_�B/��187 �uJ�8 06�9s0 rBn�1 (���202 0EW,�ѱ2^��2��90�U12�p�2��2 b��u4��2�a"RB����9\�U2�`w�l����4 60Mp��7�������b�s
5 ¿�3����pB"9 �3 ����`ڰR,:7 �2��V�2���5���2^��a^9����qr����n�5 ����5᥁"�8a�Ɂ}�5B���5����`!UA���� ��86 �+6 S�0��5�p�2<�#�529 �2^��b1P�5~�2�`���&P5��8"��5��u�!�5��ٵW544��5��R��P nB^z�c (4�����U5J�V�5��1�1^���%�����5 b2a1��gA��58W[82� rb��5N��E�5890r� 1�95 �"������ c8"a��|�L ���!�J"5|6��^!��6��B�"8�`#��+�58%�6B�AME�"�1 iC��622D�Bu�6V��d� 4��{84�`ANRSP�e/S� C�5 � �6� ��� \� �6�� �V� 3t��� �T20CA�R��8�� Hf� 1DH�� A�OE� �� ,|�� �0\�� �!64K��ԓrA� ��1 (M-7�!/50T�[PM��P�Th:1�C�#Pe� ��3�0� 5`M75cT"� �D8p� �0�Gc� u�4��i1-7'10i�1� Skd�7�j�?6�:-HS, � �RN�@�UB�f<�X�=m75sA*A�6an���!/CB�B2.6A �0;A�CIB�A��2�QF1�UB2�21� /70�S� �4��A��Aj1�3p���8r#0 B2\m*A@�C��;bi"i1K�u"A�~AAU� imm7c�7��ZA@I�@�Df��A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5�*A�EA�5B�4>\77
B7=Q�D�2�Q$BR�E7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E
"l7�@7�A
1�E�V$~`�W2%Q�R9ї@0L_�#����"Aȉ��b��H3s=rA/2�R5nR4�74rNUpQ1ZU�A�s\m9
1M92L2�!F!^Y�ps� 2ci��-?�qhimQ�t  w043�C��p2�mQ�r�H_ �H2�0�Evr�QHsXBSt62�q`s����� �<�Pxq350_*A3#I)�2�d�u0�@� �'4TX�0�pa3i1A3sQ25�c��st�r�VR1%e�q0
��j1��O2  �A�UEiy�.�‐ �0dCh20$CXB79#A��ᓄM Q1]�~�� 9�Q��?PQ��qA!P vs� 5	15aU����?PŅ���ဝQ9A6�zS*�7�qb5�1p����Q��00P(��V7]u�aitE1���À�p?7� !?�z��r=bUQRB1PM=�Q�a9��H��QQ�25L��������Q��@L���8ܰ��y00\}ry�"R2BL�t�N  ��� �1Dp�2�qeR�5���_b�3�X^]1m1lcqP1�a��E�Q� 5F����!5<���@M-16Q��  f���r��Q�e� ��8� PN�LT_�1��i1��9453��@�e�|�b1l>F1u *AY2�
��R8�Q����RJ�J3�D}T� 85
Qg�/0��*A!P@�*A�Ð𫿽�2ǿپ6t�6=Q���P�ȓ��� AQ�  g�*ASt]1^u�ajrI� B����~�|I�b��y&I�\m�Qb�I�uz��A�c3Apa9q� B6�S��S��m���}�8�5`N�N�  �(M���f1���6�����161��5�s`�SC��U��A�����5\set06c�����10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��� �5�B��B��h`�F� ��X0���A:���C�M�B��AZ��@��4�6i� ���� e�O�-	�� �f1��F �ᱦ�1pF�Y	���T6HL3���U66~`���U�dU�9D20Lf0��Qv � ��fjq��N���� ��0v
� ��i	�	.��72lqQ2�������� \chng�move.V��d����@2l_ar f	�f~��6��� ���9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�A]�,�V�1\�Qn�BJ�2W�EM!5�0��)�#:�64��F��e50S�\��0� =�PV���e�������E�����m7;shqQSH"U��)@��9�!A��(����� ,p�ॲTR1!��,�60e=�4F�����2��	 R-����� ������Ж��4���LSR�)"�!l�OA��Q�) %!� 16�
U/��2�"2��E�9p���2X� SA�/i��'�
7F�H �@!B�0��D���5V ��@2cVE��p��T�2�pt갖�1L~E�#ȚF�Q��9E�#De/��RT��59���	�A��EiR������9\7m20�20��+�-u�19r4�`�E1�= `O9`�1"ae��O2��_$W}am4�1�4�3�/d1c_std��1)�!�`_T��r�_ 4\jdg�a�q�PJ%! ~`-�r�+bgB��#Nc300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W�"Ps A��e���� t�i�P�W.��c�@FX.�e�kE14��44�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2a���2A;_2��QW2��bF�(�V11�23`�`��X5�Ra21�!J*9�a:88J99X�l5�m1a첚��*���(85�&��� ����P6���R,!52&A����,fA9INfI50\u�z�OV
 �v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&� �P1��vB)e�m������1p� �1D�p�27�F�KA�REL Use =S��FCTN��� J97�FA+�� (�Q޵�p%�)?�V�j9F?(�j�Rtk?208 "Km�6Q��y�j��iæPr�9��s#��v�krcfp�RCFt3���Q�¿kcctme�!M�E�g����6�mai�n�dV�� ��ru��kDº�c���o��L��J�dt�F ����.vrT�f������E%�!��5�FRj7%3B�K���UER�H�J�O  J�� (ڳF���F�q�Y�&T���p�F�z��19�tk vBr���V�h�9p�E�y�<�k������;�v���"CT��f�� ��)�
І��)�V	� 6���!��qFF��1 q���=�����O�?�$"����$��je���T?CP Aut�r�<�520 H5�J[53E193��9��+96�!8��9��	 n�B574��52�uJe�(�� Se%!�Y�����u��ma�Pqtool�ԕ��������conrel��Ftrol Re?liable�Rmv9CU!��H51���p�� a551e"<�CNRE¹�I�c�&��it�l\�sfutst "�UTա��"X�\u@��g@�i�6Q]V0�B$,Eѝ6A� �Q� )C���X��Yf�I�1�|6s@6i��T6AIU��vR�d�
$e%1��2�C58�E6���8�Pv�iV4OFH58�SOeJ� mvBM6E~O58�I�0�E�#+@ �&�F�0���F�P6a����)/++�</N)0�\tr1�����P �,pɶ�rmaski�msk�aA���Iky'd�h	A	�P�s�DisplayI�m�`v����J88G7 ("A��+Heůצprds��IϩǪ��h�0pl�2�R2Ƚ�:�Gt�@��PRD�TɈ�r�C�@Fm�8�D�Q�AscaҦ�� V<Q&��bVvbrl�eې@��^S��&5�Uf�j8710�yAl	��Uq���7�&��p�p��P^@�P�firmQ����Pp�2�=bk�6�r�3��6��otppl��PL���O�p<b�ac�q	��g 1J�U�d�J��gait_9e��Y�&��Qx���	�Shap��eration�0<��R67451j9:(`sGen�ms�42-f��r�p�5����2�rsgl�E��pp�G���qF�205p��5S���Ձ�retsdap�BP�O�\s�� "GCR�ö? ^�qngda�G��V��st2axU��A1a]��bad�_�>btputl/�&�|e���tplibB_��=�2.����5���gcird�v�slp���x�hex��v�rqe?�Ɵx�key��v�pm��x�us$�6�gcr��F���p���[�q27j92��v�ollismqS�k�9O�ݝ� (p#l.���t��p!o��A29$Fo8��cg7no~@�tptcls` �CLS�o�b�\�km�ai_
�s>�v�o�	�t�b���ӿ�E��H��6�1enu�501�[m��ut�ia|$calma�UR��CalMat�eT;R51%�i=1 ]@-��/V� ��Z��� �fq1�9 "K9�E�L����2m�C�LMTq�S#��et �LM3!} �F�c�nspQ�c���Oc_moq��� ��cc_e�����su���ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ���N�sve��C�clm��&Ao# �|$find�e�0STD� ter Fi�LANG���R���
��n3��z0C3en���r,���� ��J����� ���K ��Ú�=���_Ӛ���r� "FNDRК� 3��f��tguid�䙃N�."��J�tq�� �������@������J����_�� ����c��	m�Z�~�\fndr.��n#>
B2p��Z�C�P Ma�����3�8A��� c��6� ( ���N�B�������� 2�$�81��m_���"ex�z5 �.Ӛ��c��bS���efQ��	���RBT;�OPTN �+#Q�*$�r *$��*$r*$%/s#C��d/.,P�/0*ʲDPN��$���$*��Gr�$k Exc��'IF�$MASK��%93 H5�%H�558�$548 H�$4-1�$��#1(�$�0 E�$��$�-b�$���!UPDT �B�4�b�4�2�49��0�4a�3�9j0"Mx�49�4  ��4<�4tpsh���4<�P�4- DQ� �3 �Q�4�R�4�pR%0�2�r�4.b
E\���5�Ax�4��3adq\�5K979":E�ajO? l "DQ^E^�3i�Dq ��4ҲO) ?R�? ��q�5��T��3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F蠠�4��.�5y N|� �2il(in�4��31 JH1�2Q4�251ݠ�4rma	l� �3)�REo�Z_ �æOx����4��^F�?onorTf��7_ja��UZҒ4l�5rms�AU�Kkg���4�$HCd\�fͲ�eڱ�4�RE	M���4yݱ"u@�RE�R5932fO��47|Z��5lity,�Up��e"Dil\�5���o ��7987p�?�25 �3hk910 �3��FE�0=0P_>�Hl\mhm�5 ��qe�=$�^�
E�x�u�IAymptm�U0��BU��vste�y\ �3��me�b�DvI�[� Qu�:F�Ub�*_�
EL,�su��_ �Er��ox���4hGuse�E-�?�sn��������FE��,�box�����c݌,"� ������z��M��<g��pdspw)�	� �9���b���(��1���c��Y�R� � �>�P���W��������'�0ɵ�[���͂���  �� ,@� ��A�bump�šf��B*�Box%��7Aǰ60�BBw�\��MC� (6�,f��t I�s� ST ��*��}B�����=w��"BBF
�>��`���)��\bb?k968 "�4��ω�bb�9va699����etbŠ��1X�����ed	�F�b�u�f� �sea""������'�\��,� ���b�ѽ�o6�H�
�x�$�f���!y�����Q[�! tpe�rr�fd� TP�l0o� Recov�,��3D��R64�2 � 0��C@}s�� N@��(U�rroč��yu2r��  �
  �����$$CLe� ��������������$z�_DI�GIT��������.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$j���+c:PROD�UCTM�0\PG/STKD��V&oho�zf99��D����$FEAT_�INDEX��xd���  �
�`ILECOM�P ;���#���`�cSETUPo2 <�e�b?�  N �a�c�_AP2BCK �1=�i  �)wh0?{%&c����Q�xe%�I �m���8��\� n����!���ȏW�� {��"���F�Տj��� w���/�ğS������ ���B�T��x���� ��=�үa������,� ��P�߯t������9� ο�o�ϓ�(�:�ɿ ^���Ϗϸ�G��� k� �ߡ�6���Z�l� �ϐ�ߴ���U���y� ���D���h��ߌ� ��-���Q������� ��@�R���v����)� ����_�����*�� N��r��7� �m�&�3\t�i
pP 2#p*.VRc�*��� /�ƗPC/1/F'R6:/].��/+T�`�/�/F%�/�,�`r/?�*.F��8?	H#&?e<x�/�?;STM �2��?�.K �?�=�iPendant? Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OpoO�O_:JPG _�J_�56_�O_�_�	�PANEL1.D	T�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�W�I��
TP�EINS.XML��0\���q�Custom T?oolbar	���PASSWOR�DyFRS:�\L�� %Pa�ssword Config���֏ e�Ϗ�B0���T�f� ���������O��s� �����>�͟b��[� ��'���K��򯁯� ��:�L�ۯp�����#� 5�ʿY��}��$ϳ� H�׿l�~�Ϣ�1��� ��g��ϋ� ߯���V� ��z�	�s߰�?���c� ��
��.��R�d��� ����;�M���q�� ����<���`������ %���I�������� 8����n���!� �W�{"�F �j|�/�S e��/�/T/� x//�/�/=/�/a/�/ ?�/,?�/P?�/�/�? ?�?9?�?�?o?O�? (O:O�?^O�?�O�O#O �OGO�OkO}O_�O6_ �O/_l_�O�__�_�_ U_�_y_o o�_Do�_ ho�_	o�o-o�oQo�o �o�o�o@R�ov ��;�_�� �*��N��G���� ��7�̏ޏm����&� 8�Ǐ\�돀��!��� E�ڟi�ӟ���4�ß X�j��������įS���w������B�#���$FILE_DG�BCK 1=���/���� ( �)
S�UMMARY.DyGL���MD:������Diag� Summary���Ϊ
CONSLOG�������D�ӱ�ConsoleO logE�ͫ���MEMCHECK�:�!ϯ���X�Me�mory Dat�a��ѧ�{)>��HADOW�ϣ����J���Shad�ow Chang�esM�'�-��)	FTP7Ϥ�3������Z�mmen�t TBD��ѧ0�=4)ETHERNET��������T�ӱEther�net \�figurationU��ؠ��DCSVRF��߽߫�����%��� verify� all��'�1P{Y���DIFF��p����[���%��diff]�������1R�9�K��� ����X��CH�GD������c��r����2ZAS�� ��GAD���k��z��FY3bI[�� �/"GAD���s/�����/*&UPDAT�ES.� �/��FORS:\�/�-Ա�Updates �List�/��PS�RBWLD.CM�(?���"<?�/Y�P�S_ROBOWEL��̯�?�?��?&� O-O�?QO�?uOOnO �O:O�O^O�O_�O)_ �OM___�O�__�_�_ H_�_l_o�_�_7o�_ [o�_lo�o o�oDo�o �ozo�o3E�oi �o���R�v ���A��e�w�� ��*���я`������ ���O�ޏs������ 8�͟\�����'��� K�]�쟁����4��� ۯj������5�įY� �}������B�׿� x�Ϝ�1���*�g��� ��Ϝ���P���t�	� ߪ�?���c�u�ߙ� (߽�L߶��߂��� (�M���q� ���6� ��Z������%���I� ��B�����2������h����$FIL�E_� PR� ���������MDONL�Y 1=.�� 
 ���q��� �������~% �I�m�2 ��h��!/�./ W/�{/
/�/�/@/�/ d/�/?�//?�/S?e? �/�??�?<?�?�?r? O�?+O=O�?aO�?�O �O&O�OJO�O�O�O_��O9_�OF_o_
VI�SBCKL6[�*.VDv_�_.POFR:\�_�^.P�Vision VD file�_ �O4oFo\_joT_�oo �o�oSo�owo�o B�of�o�+� ������+�P� �t������9�Ώ]� 򏁏��(���L�^�� �����5���ܟk� � ��$�6�şZ��~������
MR_GR�P 1>.L~��C4  B����	 W������*u����RHB ��2 ���� ��� ���B�����Z�l� ��C���D�������Ŀ���J8�L��~%J�tF�{5U��R�S����ֿ Gn��E��.E88��-���:u�{�@ ����@A��A� f�?h�!A��r��E�� F@ �������ھ��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<,6\b�π+�&�(�a�L߅�p�A��A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�PJ��P��T���ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�O�гߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������s[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U��0
//./A�#��� �~/����/�/�/ �/� ?2?D?V?h?�/ ?�?�?�?�?�?�?� ��@O?dO�/�O�O �O�O�?�O�O__*_ MON_�Or_�_�_�_�_ 	OO-O�_A_&ouOJo \ono�o�o=o�o�o�o �oo�o4FXj |�_�_�_o�7o ��0�B�T�#x��� �������e����� ,�>�����ŏ�� �Ο������:� L�^�p�����'���ʯ ܯ� �O�a�s����� l���������ƿؿ�� ��� �2�D�g��z� �Ϟϰ����#�5�G� I��}�R�d�v߈ߚ� iϾ��������)߫��<�N�`�r��XST_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������O�C�R.RDzVT=#��K@9�BOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ�{
�Å��ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A��W�@<�P�R�
h�B�b�A��j���a��:��Dzۀ���߹�����j���( �� -��C���'�7��&���q�Y������ �?�ff ���gy ������q:a��
>N+�  PƱj�(�� ��7	���|�/?����xZ�p�<
6b<߈�;܍�<�ê�<� <�&Jσ�AI�ɳ+����?fff?I�?y&�k�@�.��J<?�`� q�.�˴fɺ�/�� 5/����j/U/�/y/ �/�/�/�/�/?�/0?q��F�?l??��?/�?+)�?�?�E��� E�I�G+� F��?)O�?�9O_OJO�OnO�Of�BL޳B�?_h�.��O �O��%_�OL_�?m_�?��__�_�_�_�_�
��h�Îg>��_Co�_goRodo�oF�GA�ds�q�C�op�o�o|�����$]Hq���D��fpC���pCHm�ZZ7t���6q�q�����N'�3A�A��AR1AO�^?�$�?�K��0±
=ç>�����3�W
�=�#�W��e���9�����{����<���(�B�u�����=B0�������	L��H��F�G���G���H�U`E���C�+����I#�I���HD�F���E��RC�j=���
I��@�H�!H�( E<YD0q �$��H�3�l�W��� {��������՟��� 2��V�A�z���w��� ��ԯ�������� R�=�v�a��������� ���߿��<�'�`� Kτ�oρϺϥ����� ���&��J�\�G߀� kߤߏ��߳������� "��F�1�j�U��y� ������������0�@�T�?�Q����(�1g��3/E�����5������q�3�8�����q4�Mgs&IB�+2D�a���{�^^	���P���uP2P7Q4_A��M0bt��R����X��/   �/ �b/P/�/t/�/ *a@)_3/�/�/�%1a�?�/?;?M?_?q?  �?�/�?�?�?�?�O 2 F�$N�vGb�/�A��@X�a�`�qC��C@�o��O2���OF� �DzH@�� F�P D���O�O�ys<O!_3_E_W_i_~s?���@@pZ�.t22!:2~
 p_�_ �_�_	oo-o?oQoco�uo�o�o�o�o��Q ���+��1���$MSKCFMA�P  �5� �6�Q�Q"~��cONREL  �
q3�bE�XCFENB?w
8s1uXqFNC_Qt�JOGOVLIM�?wdIpMrd�bKE�Y?w�u�bRU�N�|�u�bSFSPDTY�avJu�3sSIGN?QtTO1MOT�Nq�b�_CE_GRP [1p�5s\r� ��j�����T��⏙� �����<��`��U� ��M���̟��🧟� &�ݟJ��C���7��� ����گ�������4��V�`TCOM_C_FG 1q}�V�p�����
P�_AR�C_\r
jyUA�P_CPL��ntN�OCHECK ?={ 	r ��1�C�U�g�yϋ� �ϯ���������	���({NO_WAITc_L�	uM�NTX��r{�[m�_E�RRY�2sy3�� &�������r��c� ��T_MO���t��,  *A�$�k�3�PARAM:��u{��V[ﰽ�!�u?�� =9@3�45678901 ��&���E�W�3�c������{������� �����=�UM_RSPACE ��Vv��$ODR�DSP���jxOF�FSET_CAR9Tܿ�DIS���PEN_FILE�� �q��c֮�OPT?ION_IO���PWORK v_�ms �P(��R�Q
�j.j	 ���Hj&6$� R�G_DSBL  ��5Js�\��R�IENTTO>p�9!C��Pq=#��UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	�lmb�`�x7J�`������a�< ���`� ��b, H(���H3k7HS�M5G�22G�?��Gp
��
��!��'|, CR�>�>q�GsuaT��3���  �4spBpyr  ]o��*SB_����=j]��t�q� ��rna �,��~�6  ��UPQ�|N��M�,k�!�	'�� � ��I�� �  ��%�=��ͭ����ba	���I  �n @��~����p����� �N	 U�[�'!o�:q�pC\�C�@@sBq��|��� m�
�AT\��h@ߐ�n��$��Z�B\��A����p� �-�qbz �P��t�_�������( �� -��恊�n�ڥD[A]Ѻ�b4�'!��~(p �?�ff� ��
����OZ�R���8��z���>΁  Pia��(�ವ@����ک�a�c�dF#?˙���x����<
�6b<߈;����<�ê<�? <�&�o&ς)�A�lcΐI�*�?offf?�?&c�ޒ�@�.uJ<?�`��Yђ ^�nd��]e��[g��G� �d<����1��U�@� y�dߝ߯ߚ����߼� 	���-������&��~"�E�� E��?G+� Fþ��� ��������&��J�(5��bB��AT�8� ђ��0�6���>���J� n�7��[m��0��h��1��>�M�I
�@��A�[���C-�)��?Ƀ��� /�Y���Jp��vav`CH�/������}!@�I�Y�'�3A��A�AR1A�O�^?�$�?�����±
=�ç>����3�W
=�#�����+e��ܒ������{����<���.(�B��u��=B0�������	��*H�F�G����G��H��U`E���C��+�-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�? O�?3OOWOBOTO�O xO�O�O�O�O�O�O_ /__S_>_w_b_�_�_ �_�_�_�_�_oo=o (oaoLo�o�o�o�o�o �o�o�o'$] H�l����� ��#��G�2�k�V� ��z���ŏ���ԏ� ��1��U�g�R���v� ����ӟ�������-�:�(���������a����xQ�c�,!3�8�}�<��,!4Mgs�����ɢIB+կ篴a?���{����A�/�e�S���w��P!�P�������7�`�ӯ�ϑ�R9��Kτ�oχϓϥ�  ���χ����)�� M����������{߉�����ߒߤ�������  )�G�q��_���2 wF�$�&Gb����n�[ZjM!C��s�@j/�A�S���F�� Dz���� F�P D��W����)������������x?��ͫ@@
9�E��E��E��
 v����� ��*<N`ܷ*P ���˨��1��$PARA�M_MENU ?�-�� � DEF�PULSEl	�WAITTMOU�T�RCV� �SHELL_�WRK.$CUR�_STYL��,OPT�/PT�B./("C�R_DECSN���,y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?��USE_PROG %�%�?�?�3CCR�����7�_HOST !F�!�44O�:T̰�?PCO)ARC�O�;_TIME�XB��  �GDEB�UGV@��3GINP_FLMSK�O��IT`��O�EPGA�P �L��#[CH��O�HTYPE����?�?�_�_�_�_ �_oo'o9obo]ooo �o�o�o�o�o�o�o�o :5GY�}� ���������1�Z��EWORD �?	7]	RS�`�	PNS��$��JOE!>�T�Es@WVTRACE�CTL 1x-�]� ��Ӱ���ɆDT Q�y-���D 7� ��,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�T�(� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ j��_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�_����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v��������//"#�$PGT�RACELEN � #!  ���" �8&_�UP z��e�g!o S!h �8!_CFG {Fg%Q#"!x!�$�J �#|"DEFSP/D |�,!!J ��8 IN TR�L }�-" 8��%�!PE_CON�FI� ~g%��g!�$�%�$L�ID�#�-74G�RP 1�7Q!��#!A ����&ff"!A+33�D�� D]� ?CÀ A@+6�!�" d�$�9�9*1*0?� 	 +9�(8�&�"�? ´	C�?�;B@3AO�?OIO�3OmO"!>�T?��
5�O�O�N�O �=��=#�
 �O_�O_J_5_n_Y_��O}_�_y_�_�_�_ G Dzco" 
o Bo�_Roxoco�o�o�o �o�o�o�o>)�bM��;
V7�.10beta1��$  A��E�rӻ�A �" �p?!G��q>����r��0�q{�ͻqBQ��q�A\�p�q�4�q�p
�"�BȔ2�D�V��h�w��p�?�?)2 {ȏw�׏���4� �1�j�U���y����� ֟������0��T� ?�x�c�������ү�� ��!o�,�ۯP�;�M� ��q�����ο���ݿ �(��L�7�p�+9��sF@ �ɣͷ� ��g%������+�!6 I�[߆������ߵߠ� ��������!��E�0� B�{�f�������� �����A�,�e�P� ��t���������� ��=(aL^� ������' 9$]�Ϛ��ϖ� ������/<�5/`� r߄ߖߏ/>�/�/�/ �/�/?�/1??U?@? R?�?v?�?�?�?�?�? �?O-OOQO<OuO`O �O�O�O�O���O_�O )__M_8_q_\_n_�_ �_�_�_�_�_o�_7o Iot���o�o�� �o�o�o(/!L/^/p/ �/{*o����� ����A�,�e�P� b����������Ώ� �+�=�(�a�L���p� �����Oߟ񟠟� � 9�$�]�H���l�~��� ��ۯƯ���#�No`o ro�on��o�o�o�oԿ ���8J\ng� ���vϯϚ������� 	���-��Q�<�u�`� r߫ߖ��ߺ������ �;�M�8�q�\���� ����z������%�� I�4�m�X���|����� ������:�L�^��� Z���������� �$�6�H�Sw b������� //=/(/a/L/�/p/ �/�/�/�/�/?�/'? ?K?]?H?�?��?�? f?�?�?�?O�?5O O YODO}OhO�O�O�O�O �O�O&8J4_F_� ���_�_��_�_ "4-o�O*ocoNo�o ro�o�o�o�o�o�o )M8q\�� �������7� "�[�m��?����R�Ǐ ���֏�!��E�0� i�T���x�������� _$_V_ �2�l_~_�_������R�$PLI�D_KNOW_M�  �T������SV ��U͠�U��
��.�ǟR��=�O�����mӣM_?GRP 1��!`U0u��T@ٰo�
ҵ�
���Pзj� �`���!�J�_�W� i�{ύϟϱ�������X��߱�MR�����1T��s�w� s��� �޴߯߅��ߩ߻��� ��A���'���� �����������=� ��#���������}�������S��ST��1W 1��U# ���;0�_ A .�� ,>Pb���� ����3(i L^p������2*���	<-/3/)/;/M/�4f/x/�/�/5 �/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?M_AD  d#�`PARNUM  w�%OWSCH?J ME
�Gp`A�Iͣ�EUPD`O�rE
a�OT_CM�P_��B@�P@'�˥TER_CHK'U��˪?R$_6[�RSl�¯��_MO�A@�_�U_�_RE_R/ES_G �� >�oo8o+o\oOo�o so�o�o�o�o�o�o�o�W �\�_%�U e Baf�S� �� ��S0����SR0 ��#��S�0>�]�b���S�0}������RV �1�����rB@c]���t�(@c\�����D@c[��$���RTHR_�INRl�DA��˥d�,�MASS9� Z�M�MN8�k�MON�_QUEUE a���˦��x� RDNPUbQN{�P[���END���_ڙEX1E�ڕ�@BE�ʟ>��OPTIOǗ�[���PROGRAM7 %��%��ۏ��O��TASK_I�AD0�OCFG ኞ�tO��ŠDATuA���Ϋ@��27�>�P�b�t���,� ����ɿۿ�����#�x5�G���INFOU���������ϭϿ� ��������+�=�O� a�s߅ߗߩ߻���������^�jč� �yġ?PDIT �ίc���WERF�L
��
RGADoJ �n�A��¹�?����@���IOORITY{�QV���MPDSPH������Uz����OTO�Ey�1�R� (/!AF4�E�P]�~��!tcph�>��!ud��!icm��ݏ6�XY_ȡ�R�=�ۡ)� *+/ ۠�W:F �j����� �%7[B�=*��PORT#�BC�۠����_C?ARTREP
�R�> SKSTAz��Z�SSAV���n�	�2500H86A3���r�$!�R����q�n�}/x�/�'� URGE��B��rYWF� DO{�rUVWV��$�A��WRUP_DEL�AY �R��$RO_HOTk��%O�]?�$R_NORM�ALk�L?�?p6SE�MI?�?�?3AQS�KIP!�n�l#x 	1/+O+ O ROdOvO9Hn��O�G�O �O�O�O�O_�O_D_ V_h_._�_z_�_�_�_ �_�_
o�_.o@oRoo vodo�o�o�o�o�o�o �o*<Lr`���n��$RCgVTM�����p�DCR!�L���qC`N�C����C�Q?���>r��<|��{4M�g�&����/��Z��t�����l4�{�4Oi��O <�
6b<߈;�܍�>u.�?!<�&{� b�ˏݏ��8����� ,�>�P�b�t������� ��Ο���ݟ��:� %�7�p�S������ʯ ܯ� ��$�6�H�Z� l�~�������ƿ��� տ���2�D�'�h�z� ���ϰ���������
� �.�@�R�d�Oψߚ� �߾ߩ��������� <�N��r����� ��������&�8�#� \�G�����}������� ����S�4FXj |������� ��0T?x� u����'// ,/>/P/b/t/�/�/�/ �/�/�/�?�/(?? L?7?p?�?e?�?�?� �?�? OO$O6OHOZO lO~O�O�O�?�?�O�O �O�O __D_V_9_z_ �_�?�_�_�_�_�_
o o.o@oRodovo�X�q�GN_ATC 1��� AT&FV0E0�k�ATDP/6�/9/2/9�h�ATA�n,�AT%G1%B9�60�i+++��o,�aH,�qI�O_TYPE  ��u�sn_�oRE�FPOS1 1�>P{ x�o�Xh_�d_���� �K�6�o�
���.����R����{{2 1�P{���؏V�ԏz�<���q3 1��$��6�p��ٟ���S4 1�����˟����n���%�S5 1� <�N�`�����<���S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB�-�|f��S8 1������Y�������y�SMASK 1�P�  
9�G��XN	OM���a~߈Ӂq?MOTE  h�~t���_CFG ������рrPL_R�ANG�ћQ��PO�WER ��e���SM_DRY�PRG %i�%���J��TART ��
�X�UME_�PRO'�9��~t_�EXEC_ENB�  �e��GSP�D������c��TD�B���RM��MKT_!�T���`�OBOT_NAM/E i���i�OB_ORD_N_UM ?
�\q�H863 � �T���������bPC_TIME�OUT�� x�`S�232��1��k� LTEAC�H PENDAN �ǅ�}���`�Mainten�ance Con�s�R}�m
"{�dKCL/Cg��Z ��n� No Use}�	��*NPO��х����(CH�_L�������	��mMAVAI�L��{��ՙ�S�PACE1 2��| d��(>���&���p��M,8�?�ep/e T/�/�/�/�/�W// ,/>/�/b/�/v?�?Z? �/�?�9�e�a�=?? ,?>?�?b?�?vO�OZO@�?�O�O�Os�2�/O*O<O�O`O�O �_�_u_�_�_�_�_[3_#_5_G_Y_o}_ �_�o�o�o�o�o[4.o@oRodovo$ �o�o����"�	�7�[5K]o�� A����	�̏�?�&�T�[6h�z����� ��^�ԏ���&��;�\�C�q�[7������ ��͟{���"�C�� X�y�`���[8���� Ưدꯘ��0�?�`��#�uϖ�}ϫ�[G ;�i� �ϋ
G� ����$� 6�H�Z�l�~ߐ��8 ǀ������߈��d (���M�_�q��� ���������?��� 2�%�7�e�w������� �������������!� RE�W������ ����?Qw `�� @0���ߖrz	�V _�����
/L/ ^/|/2/d/�/�/�/�/ �/�/?�/�/�/*?l? ~?�?R?�?�?�?�?�? �?�?2O�?
��O�[_MODE  y�˝IS ���vO,*ϲ�O�-_��	M_v_#dCW�ORK_AD�M{,�$bR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/D���d;2BaR��WY��^����^R^	r  P���� �  �8�P�	�D��GYk}� �������Qp/@/R//<)P;�o\T���Qpg-�t��_DiKT��[  � lv%����� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OWW�# �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_olO ~Od+No`oro�o�o�o �o�o�o�o&8 J\n������u�  0�"0g�/ �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q�����$o�� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E����� Do��������ҿ��� ��,�>�P�b�tφ� �Ϫϼ���������w
�  58�J�\�n� �ߒߜկ��������� 	��-�?�Q�c�u��8���� ��- ����� �2�D�V�h� z�������������������& ���%	1234�5678�" 	��/� `r�������� (:L^p� ������ // $/6/H/Z/l/~/��/ �/�/�/�/�/? ?2? D?V?h?�/�?�?�?�? �?�?�?
OO.O@Oo? dOvO�O�O�O�O�O�O �O__*_YON_`_r_ �_�_�_�_�_�_�_o oC_8oJo\ono�o�o �o�o�o�o�oo" 4FXj|���������	��s�3�E�W�{�Cz�  Bp��   ���2���z�$�SCR_GRP �1�(�U8(ӿ\x^ �@  �	!�	 ׃��� "�$� ��-��+���R�w����D~�����#����O����M-10iAo 8909905 �Ŗ5 M61C �>4��Jׁ
� ���0�����#�1�	"�z�����h��¯Ҭ ��� c���O�8�J�� �����!�����ֿ.��B�y����������A��$�  @��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ�� ��������%��I�4� m��<�l߃ߕߧ���B���\����1� �U�@�R��v��� ��������;���*<=�
F���?�d��<�>HE����@��:��� B����ЗЙ���EL_�DEFAULT � �����B�MIPO�WERFL  ��$1 WFDO� $��ERV�ENT 1������"�pL!DUM_EIP���8��j!AF_�INE �=�!�FT���!���4 ��[!�RPC_MAI�N\>�J�nV�ISw=���!7TP�PU��	�d�?/!
PMON_PROXY@/��e./�/"Y/�f�z/�/!RDM_'SRV�/�	g�/#?G!R C?�h?�o?!
pM�/�i�^?�?!RLSY3NC�?8�8�?O�!ROS�.L�4�?SO"wO�#DOVO �O�O�O�O�O_�O1_ �OU__._@_�_d_v_ �_�_�_�_o�_?oo�coiICE_KL� ?%y (%�SVCPRG1@ho8��e���o�m3�oD�o�`4 �`5(D-�`6PU�`7x }�`���l9��{�d:?��a�o��a �oE��a�om��a�� �aB���aj叟a� ��a�5��a�]��a ����a3����a[�՟ �a�����a��%��aӏ M��a��u��a#����a K�ů�as���a��mo b�`�o�`8�}�w��� ����ɿ���ؿ��� 5�G�2�k�VϏ�zϳ� �����������1�� U�@�y�dߝ߯ߚ��� ��������?�*�Q� u�`��������� ���;�&�_�J��� n�����������sj_DEV y	��MC:Lw!`OUT"�,REC �1�Z� d   	 	�������

 �Z�{0H6l Z�~����� � //D/2/h/z/\/ �/�/�/�/�/�/�/? �/,?R?@?v?d?�?�? �?�?�?�?�?OO(O NO<OrOTOfO�O�O�O �O�O�O_&__J_8_ Z_\_n_�_�_�_�_�_ �_�_"ooFo4oVo|o ^o�o�o�o�o�o�o�o 0TBxf� ���(���,� �P�>�`���h����� ����Ώ��(�:�� ^�L���p�������ܟ ���� �6�$�Z�H� ~���r�����دƯ� ���2��&�h�V��� z�����Կ�ȿ
��� ��.�d�RψϚ�|� �Ϭ���������<� �`�N�pߖ߄ߺߨ� ��������8�&�\��J�l��jV 1��w Pl�	}� � �F��
TYPEVF�ZN_CFG ��x�d�7�GRP 1��A�c ,B� A�� D;� B����  B4�RB21HEKLL:�(
� X����%RSR����E0i T�x�������/Sew_�  ��%w������#������A�2�#�d����HK 1��� ���m/ h/z/�/�/�/�/�/�/ �/
??E?@?R?d?�?��?�?�?��OMM �����?��FTOV_ENB ���+��HOW_REG_�UIO��IMWA�ITB�JKOU�T;F��LITIM�;E���OVAL|[OMC_UNITC��F+�MON_AL�IAS ?e�9 ( he�s_(_ :_L_^_��_�_�_�_ �_j_�_�_oo+o�_ Ooaoso�o�oBo�o�o �o�o�o'9K] n����t� ��#�5��Y�k�}� ����L�ŏ׏���� ��1�C�U�g������ ����ӟ~���	��-� ?��c�u�������V� ϯ������;�M� _�q��������˿ݿ ����%�7�I���m� ϑϣϵ�`������� ߺ�3�E�W�i�{�&� �߱������ߒ��� /�A�S���w���� X����������=� O�a�s���0������� ������'9K] ����b�� �#�GYk} �:������ /1/C/U/ /f/�/�/ �/�/l/�/�/	??-? �/Q?c?u?�?�?D?�? �?�?�?O�?)O;OMO _O
O�O�O�O�O�OvO��O__%_7_�C�$�SMON_DEF�PRO ����`Q �*SYSTEM*  d=OU�RECALL ?�}`Y ( �}�4xcopy f�r:\*.* v�irt:\tmp�back�Q=>1�92.168.4��P46:8736� �R�_�_�_�K}5�Ua�_�_�V�_goyo��o}9�Ts:or�derfil.dat.l@oVo�o�o{}0�Rmdb:+o �o�Q�obt�c�_ 2o?U��
�o� �Sod�v����o�o6 Q���+ƏO `�r����*�<��ޟ ���'���K�\�n�����
xyzra?te 61 +�=� O���������504 *�үc�u� ������5�6�ٿ��� �"���5�ѿb�tφ�r�6����emp:�2164 W�����:��.��*.d����`��`�r߄ߗ�1 +� =�O�������)��� ����c�u���5� ���������"Ͻ��� ��b�t���������Q� U�����
�����N� ��hz���:��� ��
��A��d v���.;���� /��O`/r/�/ ��2��/�/? '�/K\?n?�?�� 8/��?�?�?/#/�? G/OjO|O�ߡ�3OEO�WO�O�O�O�Ɨ1356?��Ob_t_�_�/ �/4?5X�_�_�_?"? �_5X�_boto�o�ϫ_|��͐6088 Wo �o�o�o߹o�i�o` r��O��;M�� �_'_�t��c�u� ���_�_5o�gُ��� o"o���hяb�t�������$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1����?���% ֟��&�	��\�?� f���u��������ϯ ��"��F�)�;�|�_� ������ֿ��˿�� �B�%�f�I�[Ϝ�� ���ϵ�������,�� 6�b�E߆�i�{߼ߟ� ����������L�/� V��e������� �����6��+�l�O� v��������������� 2V9K�o ������� &R5vYk�� ���/��<// F/r/U/�/y/�/�/�/ �/?�/&?	??\??? f?�?u?�?�?�?�?�? �?"OOFO)O;O|O_O �O�O�O�O�O�O_�O _B_%_f_I_[_�__ �_�_�_�_�_�_,oo 6oboEo�oio{o�o�o �o�o�o�oL/ V�e����� ���6��+�l�O��v�������PARAoM �����_ �	��P�����OFT_�KB_CFG  �ヱ���PIN_�SIM  ����C�U�g�����RV�QSTP_DSB�,�򂣟����SR� �/�� & � ULTIROBOTTASK������TOP_O�N_ERR  ����PTN �/�@��A	�RING_P�RM� ��VD�T_GRP 1�<ˉ�  	���� ��������Я���� �*�Q�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߣߠ߲����� ������0�B�i�f� x������������ �/�,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZ�~���� ���/ /G/D/V/ h/z/�/�/�/�/�/�/ ?
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_�8___\_��VPRG�_COUNT�q�@���RENBU��UM�S��__UP�D 1�/�8  
s_�oo*oSo No`oro�o�o�o�o�o �o�o+&8Js n������� ��"�K�F�X�j��� ������ۏ֏���#� �0�B�k�f�x����� ����ҟ������C� >�P�b���������ӯ�ί�����UYS�DEBUG�P�P��)�d�YH�SP_PwASS�UB?Z��LOG ��U��S)�#�0� � ��Q)�
MC�:\��6���_MPAC���U���Qñ�8� �Q�SAV ������ǲ&��ηSV;�TEM�_TIME 1���[ (m��&�����}YT1SVGgUNS�P�U'�U����ASK_OPTION�P�U�Q�Q���BCCFG 3��[u� n�A�a�`a�gZo��� �ߕ��߹������� :�%�^�p�[���� ������ �����6�!� Z�E�~�i���������&�������&8�� nY�}�?�� ԫ ��(L :p^����� ��/ /6/$/F/l/ Z/�/~/�/�/�/�/�/ �/�/2?8 F?X?v? �?�??�?�?�?�?�? O*O<O
O`ONO�OrO �O�O�O�O�O_�O&_ _J_8_n_\_~_�_�_ �_�_�_�_o�_ o"o 4ojoXo�oD?�o�o�o �o�oxo.TB x��j���� ����,�b�P��� t�����Ώ��ޏ�� (��L�:�p�^����� ��ʟ��o��6� H�Z�؟~�l������� د���ʯ ��D�2� h�V�x�z���¿��� Կ
���.��>�d�R� ��vϬϚ��Ͼ����� ��*��N��f�xߖ� �ߺ�8��������� 8�J�\�*��n��� ���������"��F� 4�j�X���|������� ������0@B T�x�d���� �>,Ntb ������/� (//8/:/L/�/p/�/ �/�/�/�/�/�/$?? H?6?l?Z?�?~?�?�? �?�?�?O�&O8OVO hOzO�?�O�O�O�O�O �O
__�O@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<o^o�oro �o�o�o�o�o�o  J8n$O��� ��X���4�"��X�B�v��$TBC�SG_GRP 2��B�� � �v� 
 ?�  ������׏ �������1��U�g��z���ƈ�d,� ���?v�	 H�C��d�>�����e�CL  B�p��Пܘ������\)��Y  A��ܟ$�B�g�B�Bl�i�X�ɼ���X��  D	J���r�����C����үܬ	���D�@v�=�W�j� }�H�Z���ſ���������v�	�V3.00��	�m61c�	*`X�P�u�g�p�>���2v�(:�� ��p���  O�����p�����z�JCFG� �B��� �����������=��=�c�q� K�qߗ߂߻ߦ����� ���'��$�]�H�� l������������ #��G�2�k�V���z� ������������ �p*<N���l� ������#5 GY}h��� �v�b��>�// / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?d? R?t?v?�?�?�?�?�? O�?*OO:O`ONO�O rO�O�O��O�O�O_ &__J_8_n_\_�_�_ �_�_�_�_�_�_�_o Fo4ojo|o�o�oZo�o �o�o�o�o�oB0 fT�x���� ���,��P�>�`� b�t�����Ώ����� ��&�L��Od�v��� 2�����ȟʟܟ� � 6�$�Z�l�~���N��� ��دƯ�� �2�� B�h�V���z�����Կ ¿����.��R�@� v�dϚψϪ��Ͼ��� ����<�*�L�N�`� �߄ߺߨ����ߚ�� �����\�J��n�� ���������"��� 2�X�F�|�j������� ��������.T Bxf����� ��>,bP �t�����/ �(//8/:/L/�/�� �/�/�/h/�/�/�/$? ?H?6?l?Z?�?�?�? �?�?�?�?O�?ODO VOhO"O4O�O�O�O�O �O�O
_�O_@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<oro`o �o�o�o�o�o�o�o &�/>P�/�� �������4� F�X��(���|����� ֏����Ə0��@� B�T���x�����ҟ�� ����,��P�>�t� b������������� ��:�(�^�L�n��� ����2d�����̿ �$�Z�H�~�lϢϐ� �������Ϻ� ��0� 2�D�zߌߞ߰�j��� �������
�,�.�@� v�d��������� ����<�*�`�N��� r������������� &J\�t�� B������ F4j|��^����/�  2 6# 6&J/6"��$TBJOP_�GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� ƞ6$ @2 �"	� �C�� �&b�  Cق'�!�!>ǌ��
559>��0+1�33=��CL� fff?>+0?�ffB� J1��%Y?d7�.��/>;��2\)?0��5���;��h{CY� �  @� ~�!B�  A�P?��?�3EC�  D��!�,�0*BO���?�3JB��
:�/��Bl�0��0�$��1�?O6!Aə�3AДC�1D�G6Ǌ=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__<�O�O>B�\JU�O�HH�1ts�A@g33@?1� C�� ��@�_�_&_8_>��D�UV_0�LP�Q30O<{�zR� @�0 �V�P!o3o�_<oRifo Po^o�o�o�oRo�o�o �o�oM(�ol��p~��p4�6&��q5	V3.0}0�#m61c�$�*(��$1!6�A�� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�IR�CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;S@;Q�U�|8�`rz@/&�8�6&<��1��w�^$ESTPAR�S  *({ _#H�R��ABLE 1%�p+Z�6#|�Q�Q � 1�|�|�|��5'=!|�	|�
|��|�˕6!|�|�:|���RDI��z!ʟܟ� ��$���O������¯ԯ�����S��x# V���˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���U-����ĜP�9� K�]�o��-�?�Q�c��u���6�NUM  ��z!� �>  Ȑ����_CF�G �����!@�b IMEBF_T�T����x#��a�VE�R��b�w�a�R {1�p+
 (3�6"1 ��  6!�� �������� �9�$�:� H�Z�l�~���������@������^$��_���@x�
b MI_�CHANm� x� >kDBGLV;0o��x�a!n ETHE�RAD ?�
� �y�$"�\&�n ROUT��!�p*!*�SN�MASK�x#�255.h�fx�^$OOLOFS_�DI��[ՠ	OR�QCTRL � p+;/���/+/=/ O/a/s/�/�/�/�/�/���/�/�/!?��PE?_DETAI���PON_SVOF�F�33P_MON� �H�v�2-9S�TRTCHK ����42VTCOMPATa8�24�:0FPROG �%�%MULTIROBOTTOx!O06�PLAY���L:_INST_M�P GL7YDUS8���?�2LCK�LPKQUICKMEt ��O�2SCRE�@}�
tps�@�2�A�@�I��@_Y����9�	SR_GR�P 1�� ���\�l_zZg_@�_�_�_�_�_�^�^� oj�Q'ODo/ohoSe ��oo�o�o�o�o�o �o!WE{i�������	1234567�h�!���X�E1�V[�
 �}ipn�l/a�gen.htmno��������ȏ�~�Panel� setup̌}��?��0�B�T�f� ��񏞟��ԟ� ��o����@�R�d�v� �����#�Я���� �*���ϯůr����� ����̿C��g��&� 8�J�\�n�����϶� ��������uϣϙ�F� X�j�|ߎߠ����;� ������0�B��*N�UALRMb@G ?�� [��� ���������� ��%� C�I�z�m�������v�SEV  �����t�ECFG CՁ=]/BaA$�   B�/D
 ��/C�Wi{� ������4 PRց; �To�\o�I�6?K0(%����0���� �//;/&/L/q/\/`�/�/�/l�D ��Q�/I_�@HIS�T 1ׁ9  �(  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1 Ec0p?�?�?�?/C�� >?P=962 n?�?
OO.O�?�?�136c?|O�O�O�OAO SO�?�O__0_�O�O _Lu_�_�_�_:_�/�_ �_oo)o;o�__oqo �o�o�o�oHo�o�o%7I~��a81�o u������o� ��)�;�M��q��� ������ˏZ�l��� %�7�I�[������� ��ǟٟh����!�3� E�W����������ï կ�v���/�A�S� e�Pb������ѿ� �����+�=�O�a�s� ϗϩϻ�������� ��'�9�K�]�o߁�� �߷��������ߎ�#� 5�G�Y�k�}���� �����������1�C� U�g�y���v������� ����	�?Qc u��(���� )�M_q� ��6���// %/�I/[/m//�/�/ �/D/�/�/�/?!?3? �/W?i?{?�?�?�?�� ���?�?OO/OAOD? eOwO�O�O�O�ONO`O �O__+_=_O_�Os_ �_�_�_�_�_\_�_o o'o9oKo�_�_�o�o �o�o�o�ojo�o# 5GY�o}�������?��$UI�_PANEDAT�A 1������  	�}�0�B�T�f�x��� )����mt� ۏ����#�5���Y� @�}���v�����ן�� �����1��U�g�N�\����� �1�� Ïȯگ����"�u� F���X�|�������Ŀ ֿ=������0�T� ;�x�_ϜϮϕ��Ϲ� �����,ߟ�M�� j�o߁ߓߥ߷���� ��`��#�5�G�Y�k� �ߏ���������� ����C�*�g�y�`� ��������F�X�	 -?Qc����߫ ����~; "_F��|�� ���/�7/I/0/ m/�����/�/�/�/�/ �/P/!?3?�W?i?{? �?�?�??�?�?�?O �?/OOSOeOLO�OpO �O�O�O�O�O_z/�/ J?O_a_s_�_�_�_�O �_@?�_oo'o9oKo �_oo�oho�o�o�o�o �o�o�o#
GY@ }d��&_8_�� ��1�C��g��_�� ������ӏ���^�� �?�&�c�u�\����� ��ϟ���ڟ�)�� M�����������˯ ݯ0�����7�I�[� m����������ٿ� ҿ���3�E�,�i�P� �ϟφ��Ϫ���Z�l�}���1�C�U�g�y���)߰�#�������  ��$�6��Z�A�~� e�w��������� ��2��V�h�O������v�p��$UI_P�ANELINK �1�v� � �  ���}1234567890����	 -?G ���o�� ���a��#5G�	����p&���  R��� ��Z��$/6/H/ Z/l/~//�/�/�/�/ �/�/�/
?2?D?V?h? z??$?�?�?�?�?�? 
O�?.O@OROdOvO�O  O�O�O�O�O�O_�O �O<_N_`_r_�_�_�0,���_�X�_�_�_  o2ooVohoKo�ooo �o�o�o�o�o�o� �,>r}����� �������/� A�S�e�w�������� я���tv�z��� �=�O�a�s������� 0S��ӟ���	��-� ��Q�c�u�������:� ϯ����)���M� _�q���������H�ݿ ���%�7�ƿ[�m� ϑϣϵ�D������� �!�3�Eߴ_i�{�
 �߂����߸������ /��S�e�H���~� ��R~'�'�a��:� L�^�p����������� ���� ��6HZ l~���#�5�� � 2D��hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?�/�?�?�?�? �?�?m?OO&O8OJO \O�?�O�O�O�O�O�O �O[�_��4_F_)_j_ |___�_�_�_�_�_�_ o�_0ooTofo��o ��o��o�o�o ,>1bt��� �K����(�:� ���{O������ʏ ܏�uO�$�6�H�Z� l���������Ɵ؟� ���� �2�D�V�h�z� 	�����¯ԯ����� �.�@�R�d�v���� ����п���ϕ�*� <�N�`�rτ��O�Ϻ� Io���������8�J� -�n߀�cߤ߇����� �����o1�oX��o |����������� ��0�B�T�f���� ����������S�e�w� ,>Pbt��' �����: L^p��#�� �� //$/�H/Z/ l/~/�/�/1/�/�/�/ �/? ?�/D?V?h?z? �?�?�???�?�?�?
O O.O��ROdO�߈OkO �O�O�O�O�O�O_�O <_N_1_r_�_g_�_7O�M�m�$UI�_QUICKME�N  ���_AobRESTORE 1��  ��|��Rto�o�im �o�o�o�o�o: L^p�%��� ���o����Z� l�~�����E�Ə؏� ��� �ÏD�V�h�z� ��7�������/���
� �.�@��d�v����� ��O�Я�����ß ͯ7�I���m������� ̿޿����&�8�J� �nπϒϤ϶�a��� ����Y�"�4�F�X�j� ߎߠ߲������ߋ����0�B�T�gSC�RE`?#m�u1sco`uU2��3��4��5��6��7��8��bUGSERq�v��Tp঑�ks����4��5*��6��7��8��`�NDO_CFG ��#k  n` �`PDATE ����Non�ebSEUFRA_ME  �TA��n�RTOL_AB�RTy�l��ENB�����GRP 1��ci/aCz  A�����Q�� $�6HRd��`U������MSK  ������Nv�%��U�%���bVI�SCAND_MA�X�I��FAIL_IMG� ��PݗP#��IM�REGNUM�
�,[SIZ�n`��A�,VONT�MOU��@����2��a���a����F�R:\ � �MC:\�\wLOG�B@F� !�'/!+/O/�U�z MCV��8#UD1r&E�X{+�S�PPO�64_��0'f�n6PO��LI�b�*�#V���,�f@�'�/� =	��(SZV�.�����'WAI�/ST�AT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_�JMPERR 1��#k
  �23�45678901 dF�ψO{O�O�O�O�O �O_�O*__N_A_S_x�_
� MLOWc>8
 �_TI�=��'MPHASOE  ��F��P�SHIFT�15 9�]@<�\� Do�U#oIo�oYoko�o �o�o�o�o�o�o6 lCU�y�� ��� ��	�V�-��e2����	VSwFT1�2	V�M�� �5�1G� ����%A�  BU8̀̀�@ pك�Ӂ˂�у��z�ME�@�?�{��!c>&+%�aM1��k�0��{ �$`0TDI�NEND��\�O � �z����S��w���P���ϜRELE�Q��Y���\�?_ACTIV��<:�R�A ��e���e�:�RD� ���YBOX �9��د�6��02����190.0m.�83���254��QF�	� �X�j��1�robot����   px�૿�5pc�� ̿�����7�����-�^f�ZABC�����,]@U��2ʿ�eϢ� �ϛϭϿ����� �� �V�=�z�a�s߰�E�	Z��1�Ѧ