��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8GW�+0�$Y $DB\� 6COMW!2�MO� H.	 �\rVE�1$F8�RA{$O�UD�cB]CTMP1_FtE2}G1_�3�B�2ոGXD�#
� d $CARD_EXIST4�$FSSB_T�YP!AHKBD�_SNB�1AGN G�n $SLO�T_NUM�AP�REV4DEBU�� g1G ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�U0LEToE_OK�BUS�oP_CR�A$;4xAV� 0LACIw�1�R�@k �1$@M{EN�@$D�V��Q`PvVA{QLv� OU&R ,AЧ0�!� B� LM�_O�
eR�"CAsM_;1 xr~$ATTR4��@� ANNN@5I�MG_HEIGH|�AXcWIDTH4�VT� �UU0F_�ASPEC�A$�M�0EXP�.@A�X�f�CF�D ?X $GR� � �S�!.@B�PNFL�I�`�d� UIREx 3T!GITCH+Cj�`N� S�d_LZ`2AC�"�`EDp�dL� J�4S�0� <zNa%q;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_�S~BG CHG,I.1 [ T�`�"3I�pTYD�@*
2 3`#@� �!�B*HDDcJ* Cd�U2_�3_�4_�5_�U6_�7_�8_�9�;CO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"�P_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0��1p�34 >��DC �� Ќ@��hPV���mEX�p� �0g0xۤ�p�r
$TF��2C$MD3i�TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F�"F��40CP@�a2 6�@$�PPU�3N�)ύRևA�X�!DU��AI�3BUF�F=�@1� |pp���pPIZT� PP�M��M�y��F�SIMQSI�"ܢVAڤrT�=�w T�`�(zM��P�B�qFAkCTb�@EW�`P1�BTu>�MC�� �$*1JB8`p�*1DEC��F����Q��� ��H0CHNS_EMP1�$G��8��@!_4�3�p|@P��3�TCc�(r/�0-sx� �ܐ� MBi��!�����JR� i�SEGF�R��Iv �aR�TrpN�C��PVF4|>�bx &� �f{uJc!�Ja��� !2�8�ץ�AJ���SIZ�3S�c�B�TM���g�|��JaRSINFȑ b���q�۽�н�����L�3�B���CRC�e�3CCp��� �c��mcҞb�1J�c�P��.����D$ICb�Cq�5r�ե��@v�'����EV���zF��_J��F,pN��ܫ��?�4�0A�! � r���h�Ϩ��p�2��͕a�� �دp�R>�Dx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�IM��UR��QUA1w  $@TITO1�/S@S�!����"0�?DBPXWO��B0=!5�$SK���2M	@DBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z���LB�)$�/���� %�/��$C�!&?�$ENE�q.'*?�Ú �RE�p2(H ���O�0#$L|3$$�#�B[�;�К�FO_D��ROSr�#������3�RIGGER�6P�ApS����ETUR�N�2�cMR_8�T�Uw��0EWM��M�GN�P���B#LAH�<E���P��O&$P� �'P@D�Q3�CkD{��DQฑ�4�11��FGO_oAWAY�BMO��t�Q#!� CS_�o)  �PIS�  I gb {s�C��A��[ �B$�S��AbP�@�EW-�TNTVճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_S}V�bEXCLU�:�nONL2��S1Y�*a&�OT�a'�HI_V�4��B���_ *P0� 9�9_z��p ���A;SG�� +nrr� @6Acc*b��G�#@E��V.iHb?fANNU�N$0.$fdID�U�2�SC@�`�i�a�p�j�fb�pOGI$2,O�$FibW$}��OT9@�1 $DUMMYT��da���dn�� � �E- 7` ͑HE4(s�g�*b�SAB��SUF�FIW��@CA*=�c5�g6�a��DMSW�E. 8�Q�KEYI5���T�M�10s�qA�vIN䊱��D��/ Dބ�HOST_P! �rT��ta��tn��tsp��pEMӰV��� S�BLc ULI�0  8	=ȳ�ј �Tk0�!1 � �$S��ESAMPL���j�۰f璱f���I��0��[ $SUB �k�#0�C��T�r#a�SAVʅ��c����C��P�fP$n0E��w YN_B#2� 0Q�DI{dlpO�(��9#$�R_�I�� �ENC�2_S� 3  5�C߰�f�- �SpU����!4�"g�޲r�1T���5X� j`ȷg��0�0K�4�<AaŔAVER�qĕ�9g�DSP�v��PC��r"��(���ƓoVALUߗHE��ԕM+�IPճ��OkPP ��TH���֤��P�S� �۰F���df�J� �q��%T�ET+6� H�bLL_DU s�~a3@{��3:���OTX"���s��0�NOAUTO�!7��p$)�$�*��cT4�(�Cy�8�C, ұ"�q&�L�� _8H *8�LH  <6����c"�`, `� ��kª�q��q��sq���~q��7��8��9R��0����1��1̺U1ٺ1�1�1 �U1�1�2(�2�����2̺2ٺ2�2��2 �2�2�3J(�3��3��̺3ٺU3�3�3 �3�3�4(¸#�T�?��!9 <�9�&�z���I��1���M��QFqE@'@� : ,6���Q? �@P?Q9��5�9�E�@�A��a�A� ;p�$TP�$VA�RI:�Z���UP2f�P< ���TDe�@��K`Q�����wBAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�H  ��P�!�F@`�!>t ;E��sC�ST�D�  D���c�<� 	C�� {��_���l���R  ����FORCEUyP?b��FLUS�`�H�N>�F ���RD_CM�@E������� ��@vMP��REMr F�Q��1k@����7Q
K4	NJ�5EcFFۓ:�@IN2Q��OVO�OVA��	TROV���DyTՀ�DTMX�  ��@�
ے_PHX"p��CL��_Tp�E�@�pK	_(�Y_QT��v(��@A;Q	D� ������!0�tܑ0RQ���_��a����M�7�CL�dρRIV'�{���EARۑIOHP�C�@����B�B��C�M9@���R �GgCLF�e!DYk(�M�ap#5TuDG��� �%�qFSSD �s? P�a�!�1����P_�!�(�!1R��E�3�!3�+5�&O�GRA��7�@��i;�PW��ONn��EBUG_SD2H��P{�_E A�`�=��TER�M`5Bi5Q���ORI#e0C�9S�M_�P��e0D�9T�A�9E�9UP\�F�� -�A{�A�dPw3S@B$SEG��:� EL{UUSE.�@NFIJ�B$��;1젎4�4C$UFlP=�$,�|QR@"��_G90Tk�D��~SNST�PATx����APTHJ3Q�E�p%B`�'EC���AR$P�I�aSHFTy�A�A�H_SHORР꣦6% �0$�7PE��E�GOVR=��aPI�@��U�b �QAYLOW���IE"�r�A8��?���ERV��XQ �Y��mG>@�BN��U\��R2!P.uA�SYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC����EP;�uP;�6WOR�>@M`�0SM5T6�G3�GR��13�aPAL@���`�q�u_H � ���'TOCA�`P	P�`$OP����pѡ�`0O��R%E�`R4C�AO�p��Be�`R�Eu�h|�A��e$PWR�3IMu�RR_�cN�\�q=B I&2H���p_ADDR��H_LENG�B�q�qT�q$�R��S�JڢSS��SKN��u\�0�u̳�uٳSE�A��jrS��MN�!K������b����O�LX��p����`ACRO3pJ�@��X��+��Q��6�OUP3�b_�IX��a�a1��}򚃳���(�� H��D��ٰ��氋�VIO2S�D������	�7�L $xl��`Y!_OFFr^�PRM_��/�_HTTP_+�H:�wM (|pOBJ]"l�p��$��LE~C�d���N � \��֑AB_�Tq�b��S�`H�LVh��KR"uHITC�OU��BG�LO�q���h�����`���`SS� ���HQW�#A:�Oڠ<`�INCPU2VISIOW�͑��n��t�o��to�ٲ �IO�LN��P 8��R���p$SLob� PUT_n�$�p��P& ¢��Y F�_AS�"Q��$AL������Q  U�0�	P4A��^���ZPH�Y��-��y��U9OI �#R `�K�����$�u�"pP pk���$�����Y��UJ5�S-���NE�6WJOGKG̲DI=S�� �Kp���&�#T (�uAVF�+`��CTR�C
�FL�AG2��LG�dU� ���؜�13LG_SIZ����b�4�Xa��a�FDl�I`� w� m�_�{0a�^��c g���4�����Ǝ���x{0��� SCH_���a7�N�d�VW����E�"����4��U�M�Aљ`LJ�@�DAUf�EAU�p��d|��r�GH�b/���BO}O��WL ?��6 IT��y0�R;EC��SCR ܓ��D
�\���MARGm�!��զ ��d%�$����S����W����U� �JGM[�MN�CHJ���FNKEuY\�K��PRG���UF��7P��FWDv��HL��STP���V��=@��А�RS"��HO`����C9T�� b ��7�[�UL���@6�(RD� ����Gt��@PO��������M�D�FOCU��RG�EX��TUI��I��4�@�L� ����P����`��Pr��NE��CANA���Bj�VAILI�C�L !�UDCS_H!II4��s�O�(!"�S���S�缳!��BUFF�!Xj�?PTH$m�@��v`��D���AtrY�?P��j�3��`WOS1Z2Z3Z�8�� Z � ���[aEȤ��ȤID%X�dPSRrO��ԬzA�STL�R}�Y�&�� Y$E�C���K�&&y�� [ LQ��+0 0�	P���`#qdt
�U��dw<���_ \ �`4Г�\��Ѩ#\0�C4�] ��CL�DPL��UTRQL�I��dڰ�)�$FLAG&�� 1�#�D����'B�LD�%�$�%ORGڰ5�2�PVŇV�Y8�s�T�r�$}d^ A���$6��$�%S�`�T� �B0�4�6RCLMC�4]?o?�9�세�MI�p}d_ Yd=њRQ���DSTB�p� �;F�HHAX�R |JHdLEXCESr�8BM!p�a`�D/B�T�E��`a�p=F_A7Ji��KbOttH� K�db \Q����v$MBC�LI�|�)SREQUIR�R�a.\o�AXDEB�UZ�ALt M��c@�b�{P����2A#NDRѧ`�`d;�2��ȺSDC��N�IN@l�K�x`��X� N&���aZ���UPST�� ezrLOCf�RIrp�EX<f�A�p�9AAODA�Q��f XY�OND�rMF,Łf��s"��}%�e/� ���F�X3@IGG�� g ��t"��ܓs#4N�s$R�a%��i�L��hL�v�@�DATA#?pE�%�tR���Y�Nh t �$MD`qI}�) nv� ytq�ytHP`�P�xu��(�zsANSW�)�yt@��yuD+�)p\b���0o�i �@�CUw�V�p 0XeR;R2��j Du�{Q���7Bd$CALI�A@��G��2��R�IN��"�<E�NT	E��Ck�r^�آXb,]���_N�qlk����9�D���Bm��DI�VFDH�@���qn�I$V,��S�$��$Z�X�o�*����oH �$BELTʾu!ACCEL�8.�~�=�IRC�� �䰠D�T�8�$P)S�@�"L���r���#^�S�Eы T�PACTH3���I���3x�p�A_W��ڐ���2rnC��4�_MG�$DD��T���$FW�Rp9��I��4��DE7�PPA�BN��ROTSPCEE�[g�� J���[�C@4���$U'SE_+�VPi�ƣSYY���1 �aY�N!@A�ǦOFFܐqǡMOU��NG����OL����INC�tMa6��HB��0HBENCS+�8q9B�p�4�FDm�IN�I`x�]��B��VE��|#�y�23_UP�^��LOWL����p� B���Du�9B#P�`�x ���BCv�r�MgOSI��BMOU���@�7PERCH  ȳOV��â
ǝ ����D�ScF�@MP����� Vݡ�@y��j�LUk��Gj�p�U�P=ó���ĶTRK|��AYLOA�Q e��A��Ԓ����N`��F�RTI�A$��MOUІ�HB�BS0�p7D�5���ë�Z�D�UM2ԓS_BC?KLSH_CԒk� ���ϣ���=���xޡ �	ACLAL"�q��1м@��CHKt� �S�RTY�� ^�%E1Qq_�޴'_UM�@�C#���SCL0�r�LMT�_J1_L��9@H�qU�EO�p�b�_�8e�k�e�SPC�㡘u���N�PC�N�H�z \P��C�0~"X�T��CN_:�N�9��I�SF!�?�V ���U�/���ԒT���CB!�SH�:�� E�E1T�T����y����T��PA ��_P��_� =������!(����J6 L�@��晰OG�G�TORQU��ONֹ��E�`R��H�E�g_W2���_郅���UI�I�I��Ff`�xJ�1�~1�VC"3�0BD:B�1�@8SBJRKF�9�0DBL_SMt��2M�P_DL��2GRV����fH_��d����COS���LN H������� �!*,�aZ����fMY�_(�TH|��)THET0��NK23���"��[CB�&CB�CAA��B�"��!��!�&SqB� 2�%GTS�Ar�CIMa�����,4x#97#$DU�� �H\1� �:Bk62�:A9Q(rSf$NE�D�`AI��B+5��$̀�!A�%�5�7����LPH�E�2���2S C%C%�2-&FC(0JM&̀V�8V�8߀�LVJV!KV/KV�=KVKKVYKVgIH��8FRM��#X!KH�/KH=KHKKHYKH*gIO�<O�8O�YNUOJO!KO/KO=KUOKKOYKOM&F�2��!+i%0d�7SPBALANCE_o!�[cLE0H_�%S�Pc� &�b&�b&PFULC�h�b�g�b�%p�1k%�UTOy_��T1T2�i/�2N��"�{�t#�@Ѱ`�0�*�.�T���OÀ<�v INSE9G"�ͱREV4vͰ�l�DIF�ŕ�1llzw��1m�0OBpq�я?�MI{���n?LCHWARY�_��AB��!�$ME�CH�!o ��q�AX��P����7Ђ�`�n 
�d(�U�ROB��CRԒH���=���MSK_f`�_p P �`_��AR/�k�z�����1S�~�|�z�{���z��qI�NUq�MTCO�M_C� �q � ���pO�$N'OREn����pЂor 8p GRe��uSDZ�AB�$XYZ_DA�1<a���DEBUUq�������s z`$��C;OD�� L����p�$BUF/INDX|�c�=��MORm�t $فUA��֐����y��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p} =�C�}pt�@b�D��FRIrӚ�T��RO@ \�E�}���c�OPWO�Yq�v0Y�SY�SBU/@v�$SO!Pġd���ϪUΫ}p�PRUN����PA�D���rɡL�_O�Uo顢q�$^)�IMAG��w���0P_qIM��L�I�Nv�K�RGOVCRDt��X�(�P*�J�|��0L_�`]�L�0�RB1�����M��ED}��p 
��N�PMֲ�஑w��SL�`q�w x �$OVSL4vS;DI��DEX�� ��#���-�V} *�N4�\#�B�2�G�B�
_�M���q�E� x Hw��p�ЯATUSW���Cp�0o�s���BTM��*��I�k�4��x�\԰q�y Dw�E&���@E�r��7����З�EXE��ἱ������f q�z @�w���UP'��$�pQ�XN������ļ��� �PG΅{� h $SUB�����0_���!�M/PWAIv�P7ãՓLOR�٠F\p˕�$RCVFAILs_C��٠BWD΁|�v�DEFSP!p | Lw����p��\���UNI+������H�R�+�}_%L\pP��t�P��p�}H�> �*�j�(�s`:~�N�`KETB�%��J�PE Ѓ~��J0SIZE	 ��X��'���S�OR��FORMAT�`��c X��WrEM�t���%�UX��G�G�LI���p�  $>ˀP_SWI�p{�	 �J_PL��A�L_ �����AR��B��� C��D��$E��.�C�_�U�� � �� ���*�J3xK0����TIA4��u5��6��MOM��@������ˀB�ЃAD����������PU� NR���������m��� A$PI�6q��	�� ���K4�)6�U���w`��SPEEDgPG��������� ��4T�� � @��SAMr`��\8�]��MOV_�_$��npt5��5���1���2��������d'�S�Hp�IN� '�@�+����4(x$4+T+GAMMWf|�1'�$GET`��p���Da���

pL�IBR>�II2�$HI=�_g�t��2�&�E;��(A�.� �&LW�-6<�)56�&]���v�p��V��$PDCK���q��_?�����q�&���7��4���9+� ��$IM_SR�pD�s�rF��r�rLE���Om0H]���0���pq���PJqUR_SCR�N�FA���S_SA�VE_D��dE@�NOa�CAA�b�d@�$ q�Z�Iǡs	�I� �J �K� ����H�L�� >�"hq������ ɢ�� bW^US�A���M4���a�� )q`��3�WW�I@v�_��q���MUAo�� �� $PY+�3$W�P�vNG�{� �P:��RA��RH��RO�PL�����q� ��sJ'�X;�OI�&�Zxe8 ���m�� p��ˀ�3s�O�O�O�O�Ot�aa�_т� |�� q�d@��.v��.v��d@��[wFv��E���%��r;B�w�|�tPn���PMA�QUa ��Q8��1٠wQTH�HOLW�oQHYS��ES�F�qUE�pZB��Oτ�  ـPܐ(�AP����v�!�t�O`�q��u�"���FA��IGROG�����Q2����o�"��p��INFOҁ�׃V����R��H�OI��� (�0SLEQ����@��Y�3����Á��P�0Ow0���!E�0NU��AUT<�A�COPY�=�(/�'��@Mg�N��=��}1������ ��RG4��Á���X_�P�C$;ख�`��W���P��@�������E�XT_CYC b�HᝡRpÁ�r��_NAe!А����ROv`	�� �s ���POR_�1�E2�SRV �)l_�I�DI��T_� k�}�'���dЇ�����U5��6��7��8i��H�SdB���2�$R��F�p��GPLeAdA
�TAR�Б@�0��P�楔d7� ,�0FL`Ѧo@YN��K�M��Ck��PWR+�9ᘐ=��DELA}�d�Y�pAD�a�RQSwKIP4� �A�Z$�OB`NT����P_$�M�ƷF@\b Ipݷ�ݷ�ݷd�� ��빸��Š�Ҡ��ߠ�9��J2R�� ��� 4V�EX� TQQ����TQ������� ��`�#�RD�C�V� �`��X)�R�p�����r��~m$RGEAR_� sIOBT�2FLG��LfipER�DTC����Ԍ���2TH2N<S}� 1���uG T\0 ���u�M\Ѫ`I�d"��REF�1Á� yl�h��ENAB��cTPE�04�]�� ��Y�]��ъQn#��*���"�������2�Қ��߼���������3�қ'�9�K�]�o���P��4�Ҝ�����P�������5�ҝ!�@3�E�W�i�{��6����������������7�ҟ-?Qcu�8�Ҡ��������SMSKJÁ�l��a��EkA~�rREMOTE6�����@�݂TQ&�IO}5�IS�t�R�W@��� ��pJ����p�����E�"$DSB_S�IGN�1UQ�x�Cx\�TP��S232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+�TQ��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�PHE#�0�����p_XP�C)�$FREEFROMS	pna��GET�0��UPD��A�2�%�SP|� :��� !$USAN�na&����ERI�0�Rp�RYq5*"_j@�P8m1�!�6WRK9K�D���6��QFRIgEND�Q�RUFg��҃�0TOOL�6M�Y�t$LENG�TH_VT\�FI!R�pC�@ˀE> +IOUFIN-RM���RGI�1ÐAIT�I�$GXñ3IvFG2v7G1���p3�BơGPR�p�1F�O_0n 0��!RE��p�53҅U�TC��3A�A��FU�G(��":���e1n!��J�8�%����%]��%�� 74�OX O0�L��T�3H&��8���%b4J53GE�W�0�WsR�TD����T��M�����Q�T]�$V C2����1�а91�8��02�;2k3�;3 �:ifa�9-i�aQ���NS��ZR$V��2BVwEV�2A Q�B;�����&�S�`��F`�"�k�@�2a�PS�E��$r1C��_g$Aܠ6wPR��7vMU�cS�t '��529�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx_�����BSOC����N��DUMMY�14�p@SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW_C��U��S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}����_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�SQ�pC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EG� �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G + AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC  o�ER|f�5� � $�@�_ A��!�PO���à�0#�
�_M�RAt�� d r� T��ٔERR��L=�;TY&���I��qV�0�cz�TOQ�dB�PL[ �d�"��	���C! � p�p`T)0���_V1�Vr�aӔ����2ٛ2�E����@�H�E���G$W�����V!��$�P��o�c�I��aΣ	 HEL�L_CFG!�� 5��B_BA�Sq�SR3���� a#Sb���1��%��2��3��4���5��6��7��8���RO����I0�03NL�\CAB+�����ACK4�����,��\@2@�&�?�_PUf�CO. U�OUG�P~ ����m�������{TPհ_KAR�Ll�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h�8�]�l0SEM�4Ĳ(�M4�6�TYN�SO���DIZ�~�AӸ����m_TM�MOANRQ��k0E�����$KEYSWITCH���m���{HE��BEAT��E- LE~����ȅU��F!Ĳ���B�O�_HOM=OGREFUPPR&��y!�� [�C��O��-E�COC��Ԯ0_IO#CMWD
�a��m��� � Dh1���	UX���M�βgPgC�FORC��� 챒m�OM.  �� @�5(�U�#P�, 1��, 3��4�5��NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�� �� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E�VP���UPDs� � �`NЦ�5�YS�LOt�� � �L��d���A�aTAp�0d��|�ALU:eLd�~�CUѰjgF!a�ID_L�ÑeHI��jI��$FILE1_���d��$2�f;SA>�� hO��`?E_BLCK��b|$��hD_CPUy@M�yA��c�o�da�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA�i�J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP��_(�g�����pr��� `�`GROU�w`��B��NFL�IC��f�REQUwIRE3�EBU�0�qB���w�2����p����q5�p�� \^��APPR��C}��Y�
ްEN٨CL9O7��S_M��H����u�
�qu�� ���MC�����9�'_MG��C�Co��`pM�в�N�BRKL�GNOL|�N�[�R���_LINђ�|�=�J����Pܔ�������� ���������6ɵ��̲8k����q���G� ��
��q)�<�7�PATH3�L�@B�L��H�wࡠ�J�CN�CA�Ғ�ڢ6B�IN�rUCV�4aZ��C!�UM��Y,���aE�p����������PAYLOAJ2L`R_A	N�q�Lpp����$�M�R_F2LS3HR��N�LOԡ��Rׯ�`ׯ�ACRL�_G�ŒЛ� ��H�j`߂$HM���FWLEXܣ�qJ�u� :���� ���������1�F1�V�j�@�R�d�v�������E����ȏ ڏ����"�4�q��� 6�M���~��U�g�y�$ယT��o�X��H� �����藕?����� ǟِݕ�ԕ�����%�7��JJ�� �� V�h�z���`A�T�採@�EL�� �S��J|�Ŝ�J�Ey�CTR��~�T�N��FQ��HAN/D_VB-���v`n�� $��F2M����ebSW?��'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)�F�AW�Z`i�Aw�A���X X�'pi�Dw�Dʆ�Pf�G�p�)ST�k��!x��!N��DY �pנM�9$`%Ц�H� �H�c�׎���0� ��Pѵڵ������p������ ����1��R�6��QAS�YMvř���v��pJ���cі�_SH>� �ǺĤ�ED����������J�İ%��C�I\Dِ�_VI�!X|�2PV_UNIX�FThP�J��_R�5_R c�cTz�pT�V��@��� İ�߷��U ����_ �T��Hqpfˢ��aEN�&3�DI����O4d`J�� x g"IJAAȱz�aabp�coc��`a�pdq�a� �^�OMME��� h�b�RqAT(`PT�@ � S��a7�;�Ƞ�@ȷh�a�iT�@<� �$DUMMY9�Q�$PS_��R�FC�  S�v ��p���Pa� XXƠ���STE����SBRY�M21_�VF�8$SV_E�RF�O��LsdsCLRJtA��Odb`�O�p � D ?$GLOBj�_LO���u�q�cAp�rܛ@aSYS�qADqR``�`TCH  � ,��ɩb�oW_NA����7��SR���l ���
*?�& Q�0"?�;'?�I)?�Y) ��X���h���x����� �)��Ռ�Ӷ�;��Í�v�?��O�O�O�D�XOSCRE栘p�����ST��s}�y`����%��/_HA�q� TơgpTYP�b����G�aG���Od0IS_䓀d�;UEMd� ����p�pS�qaRSM_��q*eUNEXCE1P)fW�`S_}pMрx���g�z�����ӑC�OU��S�Ԕ 1-�!�UE&��Ubwr���PROGM�F�L@$CUgpP�O�Q��5�I_�`H>� � 8�� �_HE�PS�#��`?RY ?�qp�b���dp�OUS>�� � @6p�v�$BUTTp�R|pR�COLUMq�<e��SERV5��PANEH�q� w� �@GEU��Fy��)$HE�LPõ)BETERv�)ෆ���A  � ��0��0��0�ҰIN簪c�@N(��IH�1��_�o ֪�LN�r'� �qpձ_ò=��$H��TEX8l����FLA@��/RELV��D`���������M��?,@�ű�m����"�USRVIEW�q�� <6p�`U�`��NFI@;�FOsCU��;�PRI@�m�`�QY�TRI}P�qm�UN<`�Md� #@p�*eW�ARN)e6�SRT+OL%��g��ᴰ�ONCORN��RA�U����T���w�V�IN�Le� =$גPATH9�ג�CACH��LOG�!�LIMKR���x�v���HOST��!�b�R��OgBOT�d�IM>�	 �� ���Zq��Zq;�VCPU_�AVAIL�!�EX	�!AN���q�`�1r��1r��1 ��\��p�  #`C�����@$TOOLz�$��_JMP�� ���e$S�S����VSHI9F��Nc�P�`ג��E�ȐR����OS�UR��Wk`RADILѮ��_�a��:�`9a��`a�r��LULQ�$OUTPUTg_BM����IM��AB �@�rTILNSCO��C7� ������&�� 3��A���q���m�I�2G��o�y@Md9�}��yDJU��N��WAIT֖�h}��{�%! NE�u��YBO�� �� $`�t��SB@TPE��NECp�J^FY�nB_T��R�І�a�$�[YĭcB��dM ���F� �p�$�pvb�OP?�MAS�W_DO�!QT�p�D��ˑ#%��p!"D�ELAY�:`7"JOY�@(�nCE$���3@ �xm��d�pY_ [�!"�`�"��[���P�? EaZAB�C%��  $��"R��
E`�$$�CLAS�������!pE`� � V�IRT]��/ 0AB�S����1 5�� < �!F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZi{0-�AXL�p��"��63  �{tIN8��qztPRE�����v�p�uLARM�RECOV �9�rwtNG�� �.;	 =#�
��.�0PPLIC���?5�p��HandlingTool o�� 
V7.50�P/23 �!�P�B��
��_S�Wt� UP�!�� x�F0��t���A�0v� 86-4�� �it�y�� N2 �7DA5�� j�� QB@<��o�Noneisͅ�˰ ��T��]�!LAAx-yrP_l�V�uT�:�s9�UTO�"����t�y��HGAPO�N
0g�1��Uh�D� 1581�����̟ޟry����Q 1���p� ,�蘦���;�@��q�_��"2 �3c�.�H����D�HTTHKY X��"�-�?�Q���ɯ ۯ5����#�A�G�Y� k�}�������ſ׿1� ����=�C�U�g�y� �ϝϯ�����-���	� �9�?�Q�c�u߇ߙ� �߽���)�����5� ;�M�_�q����� ��%�����1�7�I� [�m����������! ����-3EWi {������ )/ASew� ���/��/%/ +/=/O/a/s/�/�/�/ �/?�/�/?!?'?9? K?]?o?�?�?�?�?O��?�?�?O#O]���T�O�E�W�DO_C�LEAN��7��CN�M  � ��__/_A_S_�D?SPDRYR�O��HIc��M@�O�_�_ �_�_oo+o=oOoao�so�o�o���pB��v �u���aX�t����|��9�PLUGG����G��U�PRCvPB��@��_�orOxr_7�SEGF}�K[mwxq�O�O������?rqLAP �_�~q�[�m������ ��Ǐُ����!�3�>x�TOTAL�f y�x�USENU�p©� �H���B��RG�_STRING �1u�
��Mn�S5�
ȑ_�ITEM1Җ  n5�� ��$�6�H� Z�l�~�������Ưد����� �2�D��I/O SIGN�AL̕Try�out Mode�ӕInp��Simulatedב�Out��O�VERR�P = �100֒In �cycl��בP�rog Abor���ב��Stat�usՓ	Hear�tbeatїM?H Faul��Aler'�W�E�W� i�{ύϟϱ������� �CΛ�A���� 8�J�\�n߀ߒߤ߶� ���������"�4�F�pX�j�|���WOR{p Λ��(ߎ����� �� $�6�H�Z�l�~����� ���������� 2PƠ�X ��A {������� /ASew������SDEV [�o�#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y?PALTݠ1�� z?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O��O�O�O_�?GRI �`ΛDQ�?_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|�� �������0�xB�T��oPREG�> �� f���Ə؏��� � �2�D�V�h�z��������ԟ���Z���$ARG_��D �?	���;���  w	$Z�	[O��]O��Z�p�.�SB�N_CONFIG� ;��������CII_SAV/E  Z������.�TCELLSE�TUP ;�%�HOME_IO�Z�Z�%MOV_8��
�REP�lU��(�UTOBACK�ܠ��F�RA:\z� X\�z�Ǡ'`�z����ǡi�INI�0�z���n�MESSAG���ǡC���ODE_D�������%�O�4�n�PAU�SX!�;� ((O>��ϞˈϾ� �����������*� `�N߄�rߨ߶�g�l ?TSK  wͥ�<_�q�UPDT+���d!�A�WSM_kCF��;���|'�-�GRP 2:�V?� N�BŰA�߾%�XSCRD1�1�
7� �ĥĢ ����������*��� ����r����������� 7���[�&8J\�n��*�t�GRO�UN�UϩUP_kNA�:�	t�n�_ED�17��
 �%-BCKEDT-�2�'LK�`���-t��z�q�q�z���2t1������q�k�(/��ED3/��/�.a/8�/;/M/ED4�/t/�)?�/.?p?�/�/ED5`??�?<?.�?8O�?�?ED6O�?�qO�?.MO�O'O9OED7�O`O_�O.�O8\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o�_�	-9o�oo%oCR _ 9]�oF�o��k� � NO_DE�L��GE_UN�USE��LAL_OUT �����WD_ABO�Rﰨ~��pITR�_RTN��|N'ONSk���˥�CAM_PARA�M 1;�!�
 �8
SONY �XC-56 234567890� ਡ@����?��( АP\�
���{����^��HR5q�̹��ŏR�57ڏ�Aff���KOWA S_C310M
�x�}̆�d @<� 
���e�^��П\ ����*�<��`�r��g�CE_RIA_UI�!�=�F��}�z� ��_�LIU�]���ꋐ<��FB�GP ]1��Ǯ��M�_�q�0�C*  �����C1��9��@Ҩ�G���CR�C]���d��l��s��R������[Դm��vꨰ������� +C����(������=�HE�`ONFI�ǰ�B�G_PRI 1�{V���� �ϨϺ����������CHKPAUS��w 1K� ,!u D�V�@�z�dߞ߈ߚ� �߾������.��R��<�b���O��x������_MOR��� ���!C4<<��� 	 ��� ��*��N�<����䡑��?��q?;�;�����K��9�P��|�ça�-:���	�

��M��@�pU�ð��<��,~���DB���튒)�
mc:cpmi�dbg�f�:�JI�I�¥�p��/�  � W �M�� ��s>�  �ݕ�U�?U��p�pUg��/� ���PWf��M/w�O/�
DEFg l��s)��< buf.txt s/�t/��ާ�)��	`�����=L�m��*MC��1��a��?43��1����t�īCz  B�HH�CPUeB��$�B^O�:���
C���B��bY
K�D�ny�D��C�|@�>s��D�� �C�g�=F�&��E�CeE�d��Bn"�F��E�_Y	��!,�&w�1���s�e��.�p ��1�BDw�M@x8��1eҨ����g@D�p@�0EYK�EX��EQ�EJP� F�E�F�� G��>^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE ���F 
Q��;��(P  B_<_��R¯���	op6��A�Y
s@ ]AQ�2s@�C�0B3�MaC{@@�*cw��UT�pFP?ROG %�z�o�oigI�q���v��ld�KEY_TBL � �&S�#� �	
��� !"�#$%&'()*+,-./01i��:;<=>?@A�BC� GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������vq���͓���������������������������������耇����������������������p`LCK�l4�p`��`STAT ��S_AUTO_DO����5�INDT_'ENB!���R�Q?��1�T2}�^�STO�Pb���TRLr`L�ETE��Ċ_S�CREEN ~�Zkcsc���U��MMENU �1 �Y  <�l�oR�Y1�[��� v�m���̟�����ٟ �8��!�G���W�i� �������ïկ��4� ��j�A�S���w��� ��迿�ѿ����T� +�=�cϜ�sυ��ϩ� ��������P�'�9� ��]�o߼ߓߥ���� ����:��#�p�G�Y� ����������$� ���3�l�C�U���y� ���������� ��	�VY)�_MANU�AL��t�DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�mg�(&/~&lMZ�IdPx�@P@#ONTIM6ه� d�`&��
�e�MOTNE�ND�o�RECO_RD 1(�[g2�/{�O��!�/k y"?4?F?X?�(`?�? �/�??�?�?�?�?�? )O�?MO�?qO�O�O�O BO�O:O�O^O_%_7_ I_�Om_�O�_ _�_�_ �_�_Z_o~_3o�_Wo io{o�o�_�o o�oDo �o/�oS�oL �o����@�� �+�yV,�c�u�� ������Ϗ>�P��� ��;�&���q���򏧟 ��P�ȟ�^������ I�[����� ���$��6�������jTO�LERENCwB����L�͖ C�S_CFG )��/'dMC:�\U�L%04d.'CSV�� c��/#[A ��CH��z� �//.ɿ��(S�R�C_OUT *���1/V�SGN� +��"��#��10-FEB-�20 17:32~027-JANp��21:48+ P;��ɞ�/.���f�pa�m�?�PJPѲ���VERSION �Y�V2.�0.�ƲEFLO�GIC 1,� 	:ޠ=�ޠ�L��PROG_E�NB��"p�ULS�k' ����_WRSTJNK ��"f�EMO_OPT_�SL ?	�#
� 	R575 /#=�����0�B��>��TO  �ݵ�l���V_F EX��d�%��PATHw AY�A\�����5+ICT�F�u-�j�#�egS�,�ST?BF_TTS�(�	�d���l#!w�� M�AU��z�^"MSWX�.�<�4,#�Y�/�
!J�6%�ZI~m��$SB�L_FAUL(�0��9'TDIA[�1�<�<� ����12345678#90
��P��H Zl~����� ��/ /2/D/V/h/��� P� ѩ �yƽ/��6�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�,/�gUMP���� ��ATR���1OC@P�MEl�OOY_TE{MP?�È�3F�8��G�|DUNI��.��YN_BRK �2_�/�EMGDI_STA��]�'�@�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�Q�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��QDzr�=#�דQXT_BWD��p��xf́t�_DIn�� 9�5�d��T�QsRֆSTEP���:P�OP_D�Ov�f�PFAC�TORY_TUN�wdM�EATUROE :�5̀rQ�Handl�ingTool ��� \sfm�English �Dictiona�ry��roduAA Vis�� Master��ީ�
EN̐nalog I/O��ީ�g.fd̐ut�o Softwa�re Update  F OR��matic Ba�ckup��H59�6,�ground Editޒ�  1 H5�Camera�F���OPLGX�elyl𜩐II) X�7ommՐshw���7com��co����\tp���pan}e��  opl���tyle sel�ect��al C�nJ�Ցonit;or��RDE���tr��Relia�b𠧒6U�Dia�gnos(�푥�5�528�u��he�ck Safet�y UIF��En�hanced Rob Serv%��q ) "S�r�U?ser Fr[������a��xt. D�IO �fiG� �sŢ��endx�Ekrr�LF� pȐ�ĳr됮� ���� � !��FCTN /Menu`�v-�ݡ|���TP Inې�fac�  ER_ JGC�pב_k Exct�g���H558��igh�-Spex�Ski~1�  2
P���?���mmunic�'�ons��&�l�uqr�ې��ST Ǡ���conn��2ި�TXPL��nc=r�stru�����"FATKA�REL Cmd.� LE�uaG�54�5\��Run-T�i��Env��d�
!���ؠ++�s�)�S/W��[�LicenseZ��� 4T�0�ogB�ook(Syڐm�)��H54O�MA�CROs,\�/O�ffse��Loa��MH������r,� k�MechStop Prot����� lic/�MiвShif����ɒ�Mixx��)���x�SPS�Mode �Switch�� �R5W�Mo�:�.�� 74 ����g��K�2h�ult�i-T=�M���LN (Pos�Regiڑ������|d�ݐt Fun��⩐.�����Numx~����� lne�|�ᝰ Adjup������  - W���tatuw᧒T��RDMz�o}t��scove U�9���3Ѓ�uest 492�b*�o�����62;�?SNPX b ����8 J7`���Li3br��J�48����"�� �Ԅ�
�6O��� Parts i�n VCCMt�3�2���	�{Ѥ�J9�90��/I� 2� P��TMILI�B��H���P�A�ccD�L�
TE�$TX�ۨ�ap1�S�Te����pke�y��wգ�d���Unexcep=tx�motnZ���������є�� qO���� 90J��єSP CSXC`<�f��Ҟ� Py�sWe}���PRI��>vr�t�menz�� ��iPɰ�a�����vGri=d�play��v���0�)�H1�M-�10iA(B20�1 �2\� 0\}k/�Ascii��l�Т�ɐ/�Col���ԑGuar� �
�� /P-�ޠ"Kv��st{Pat �:�!S�Cyc��΂�orie��IFn8�ata- quҐ��� ƶ��mH57m4��RL��am����Pb�HMI D�e3�(b����PC�Ϻ�Passwo�+!��"PE? Sp�$�[���tp��� vKen��Tw�N�p��YELLOW B�OE	k$Arc��v�is��3*�n0W�eldW�cialh�7�V#t�Op�����1y� 2F�a�portN�(�p�T1�T� �� �ѳxy]�&TX��t�w�igj�1� b� �ct\�JPN �ARCPSU P�R��oݲOL� S;up�2fil� &�PAɰאcro�� �"PM(����O$SuS� eвtex�ԣ r���=�t�s'sagT��P���P@�Ȱ�锱�rt�W��H'>r�dpn��n1
t�!�� z ��ascbi?n4psyn��+A}j�M HEL��NCL VIS �PKGS PLOA`�MB �,�4�VW�RIPE �GET_VAR {FIE 3\t���FL[�OOL: �ADD R729.FD \j8'�iCsQ�QE��DVvQ��sQNO WTW�TE��}PD  ��^��biRFOR ���ECTn�`��ALSE ALAfP�CPMO-130�  M" #h�D�: HANG F�ROMmP�AQfr���R709 DR�AM AVAIL?CHECKSO!���sQVPCS SU��@LIMCHK �Q +P~dFF PO�S��F�Q R59�38-12 �CHARY�0�PR�OGRA W�SwAVEN`AME�P�.SV��7��$E�n*��p?FU�{�TR}C|� SHADV0�UPDAT KC|JўRSTATI�`~�P MUCH y��1��IMQ MO?TN-003��}��ROBOGUIDE DAUGH�a8���*�tou�����I� Šhd�ATH|�PepMOVET��ǔVMXPACK� MAY ASS�ERT�D��YCL�fqTA�rBE C�OR vr*Q3rA�N�pRC OPToIONSJ1vr̐PSH-171Z@-x�tcǠSU1�1`Hp^9R!�Q�`_T�P���'�j�d{tb�y app wac 5I�~d�PHI����p�aTEL�MX?SPD TB5bLu� 1��UB6@�qEN�J`CE2�61��p���s	�may n��0� R6{�R� >�Rtraff)��� 40*�p��fr���sysvar ?scr J7��cNj`DJU��bH �V��Q/�PSET �ERR`J` 68���PNDANT �SCREEN U�NREA��'�J`D��pPA���pR`IgO 1���PFI�p}B�pGROUN�P�D��G��R�P�QnRS�VIP !p�a�PD�IGIT VER�S�r}BLo�UEW~ϕ P06  �!��MAGp�abZV��DI�`� SS�UE�ܰ�EPL�AN JOT` D�EL�pݡ#Z�@D�͐CALLOb�Q �ph��R�QIPN�D��IMG�R7{19��MNT/�PWES �pVL�c���Hol�0Cq���tP�G:�`C�M�caynΠ��pg.v�S�: 3D mK�v_iew d�` �p���ea7У�b� o�f �Py���ANN�OT ACCESGS M��Ɓ*�t47s a��lok��Flex/:�Rw�!mo?�PA?�-�����`n�pa S�NBPJ AUTO-�06f����TB���PIABLE1q �636��PLN:Y RG$�pl;pNW7FMDB�VI���t�WIT 9x�0@o���Qui#0�ҺPN� RRS?pUSB��� t & remov�@ )�_��&�AxEPFT_=� �7<`�pP:�OS�-144 ��h qs�g��@OST� �� CRASH �DU 9��$�P�pW� .$��L/OGIN��8&�J���6b046 issue 6 Jg���: Slow ��st��c (HCos`�c���`IL`�IMPRWtSPO�T:Wh:0�T�S�TYW ./�VMGqR�h�T0CAT��hos��E�q���� �O�S:+pRSTU' k�-S� ����E:��pv@�2�N� t\hߐ��m ���all��0�  �$�H� WA͐��3 CNT0 T��� WroU�alacrm���0s�d � @�0SE1���r R{�OMEBp���K� �55��REàSEs�t��g    } �KANJI��no���INIS?ITALIZ-p�d�n1weρ<��dr�� lx`�SCI�I L�fail�s w�� ��`�YSTEa���o��PvЧ IIH���1W�G�ro>Pm ol\�wpSh@�P��Ϡn� cflxL@АW{RI �OF Lq���p?�F�up��d�e-rela�d� "APo SY�c}h�Abetwe:0IND t0$gb#DO���r� `��GigE�#ope�rabilf  P�AbHi�H`��c�le{ad�\etf�P8s�r�OS 030��&: fig��GL�A )P ��i��7�Np tpswx�B��If�g�������5aE�a EXC�E#dU�_�tPCLO�S��"rob�NTdpFaU�c�!����PNIO V750�Q1��Qa��'DB ��P M�+Pv�QED�DET���-� \rk��ON�LINEhSBUG�IQ ߔĠi`Z�IB�S apABC �JARKYFq� ����0MIL�`� R��pNД �p0GAR��D*pR��P�"'! jK�0cT�P��Hl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P��`WIBPK05��!FȐB/��BUSY RUNN��C "�򁐈��R-p��LO�N�DIV�Y�CUL��fsfoaBW�p����30	V��ˠIT�`�a505.�@O=F�UNEX�P1bҬaf�@�E��SVwEMG� NMLq�� D0pCC_SA�FEX 0c�08"qD. �PET�`N@�#'J87����RsP�TA'�M�K�`K��H GUNCHG^۔MECH�pMcz� T�  y, g@��$ ORY LE�AKA�;�ޢSP�Em�Ja��V�tGR�Iܱ�@�CTLN�TRk�FpepR��j50�EN-`IN�����p �`�Ǒ�k!��T3/dqo�SKTO�0A�#�L�pA �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`D	U��aO�supk�t4� � P�F� Bnf��Q�PSVGN-18��V�SRSR)J�UP�a2�Q�#D�q� l O��QBRKCTR5Ұ�|"-��r�<pc�j!INVP�D ZO� ��T`�h#�Q�cHset,x|D��"DUAL� �w�2*BRVO117 A]�TNѫt�+bTa2473��q.?���sAUz�i�B�complete���604.� -^�`hanc�U�� F��e8��  ��npJtPd!q��`��w� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP��R�R(}\xPe� aʰ�I���E��1��p�� j  �� xSP�^P �A�AxP�q �5 sig��a��"AC;a��
�bCe�xPb_p��.pc�]l<bHbcb_cicrc~h<n�`tl1� ~`xP`o�dxP�b]o2�� �cb�c�ixP�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`�cptlibxzxP�l�cr�xrxP\�blpsazEdxP_fm�} gcxP�x���o|sp�or�mc(��ob_jzo"p�u6�wf��t���wms�1q��sld�)��jmc�o\�n�b�nuhЕ��|st�e���>�pl�qp�iwc1k���uvf0uߒ<��lvisn�CgoaculwQ
E �F  ! Fc.f9d�Qv�� qw����Data Acq/uisi��nF�|1��RR631`��TR��QDMCM �2֝P75H�1�P58�3xP1��71��559`�5�P57<PxP�Q����(���Q���o pxP!daq�\�oA��@�� �ge/�etdms�"�DMER"؟,�p#gdD���.�m���-��qaq.<᡾xP#mo��h���f{�u��`13��MACRO�s, SksaffP�@z����03�SR�QT(��Q6��1�Q9ӡ��R�ZSh��PxPJ6+43�@7ؠ6�P�@�PRS�@���e �Q��UС PIK�Q5?2 PTLC�W���xP3 (��p/O ��!�Pn �xP5���03\sfmn�mc "MNMCPq�<��Q��\$AcX�FM���ci,Ҥ�X�����cdpq+�
�sk��SK�xP�SH5�60,P��,�y�r�efp "REF�p�d�A�jxP	�of��OFc�<gy�to��TO_����ٺ����+je�u��caxis2�xPE�\�}e�q"ISDTc�|�]�prax ���MN��u�b�is�de܃h�\�w�xP!� isbasic���B� P]��QA7xes�R6�������.�(Ba�Q�ess��xP���2�pD�@�z�atis�� ��(�{�����~��m��FMc�u�{�
���MNIS��ݝ�� ��x����ٺ��x�� j75��Dev�ic�� Inte�rfac�RȔQJ�754��� xP�Ne`��xP�ϐ2��б����dn� "�DNE���
tpodnui5UI��ݝ	bd�bP�q_rsofOb
?dv_aro��u�����stchkc��z	 �(}�onl��G!ff L+H�J(��"l"/��n�b��z�haSmp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!2���xpc_2pcch=m��CHMP_�|8бpevws��2�ΌpcsF��#C �SenxPacro0�U·�-�R6�Pd�@xPk�����p��gT�L��1d M�2`��8��1c4ԡ�3 qem��GEM,\i(��Dgesnd�5���H0{�}Ha�@sy���c��Isu�xD��Fmd ��I��7�4���u���AccuCal�P��4� ��ɢ7ޠB0���6+6f�6��9!9\aFF q�S(�U��2�
X�p�!Bd�ѳcb_�SaUL�� � �� ?�ܖto���otplus\tsrnغ�qb�W�p��t���1��To�ol (N. A�.)�[K�7�Z�(P��m����bfclls� k94�"K4p���qtpap� �"PS9H�stpswo��p�L7��t\�q����D�yt5� 4�q��w�q��� �Mz�uk��rkey�����s��}t�sfe7atu6�EA��� cf)t\Xq�����df�h5���LRC0�md�!�587���a�R�(����2V��8lc?u3l\�pa3}@H�&r-�Xu���t,�� �q "�q�Ot��~ ,���{�/��1c�}����y�p�r��5����S�XAg�-�y���Wj�874�- iR�Vis���Queu�� Ƒ�-�6�1$���(����u����tӑ����
�tpv�tsn "VTS�N�3C�+�� v\pR�DV����*�prd�q\�Q�&�vst�k=P������nmx&_�դ�clrqν���get�TX��Bd���aoQϿ�0q�str�D[� ��t0�p'Z����npv��@�enlIP0��D!0x�'�|���sc ߸��tvo/��2�q���vb����q����!���h]��(� Control�PRAX�P5��5�56�A@59�P5-6.@56@5A��J69$@982 �J552 IDVR7�hqA���16�Hx���La�� ���Xe�frlparwm.f�FRL��am��C9�@(F �����w6{���A���QJ643�� 5}0�0LSE
_p�VAR $SGS�YSC��RS_UNITS �P�2�4�tA�TX.$VN�UM_OLD 5`�1�xP{�50+��"�` Funct ���5tA� }��`#@�`E3�a0�cڂ��9����@H5נ� �P���(�A����۶}�����ֻ}��bPR�b�߶~ppr4�TP�SPI�3�}�r�10�#;A� t�
`���1���96�����%C�� Aف��J�bIncr�	����\�`��1o5qni4�MNINp	xP�`����!��Hour_  � 2�21 �A�AVM���0 ���TUP ��?J545 ���6162�VC�AM  (��CLIO ���R6�N2�MSC� "P ��STYL�C�28�~ 13\�NRE� "FHRM S�CH^�DCS}U%ORSR {b��04 �E�IOC�1 j 5742 � os| �? egist��Ի��7�1�oMASK�934"�7 ��OCO ���"3�8��2���� 0 HB��ڢ 4�"39N� R�e�� �LCHK�
%OPLG%��3�"%MHCR.%MCd  ; 4? ��6 d�PI�54�s� D[SW%MD� pQ�K!637�0�0p"�Y1�Р"4 �6<2?7 CTN K � +5 ���"7��<2�5�%/�T�%FRD�M� �Sg!��9�30 FB( NBA��P� ( HLB  7Men�SM$@jB�( PVC ��290v��2HTC�C?TMIL��\@?PAC 16U�hA�J`SAI \@ELN���<29s�UE�CK �b�@FRM� �b�OR���I�PL��Rk0CSXsC ���VVFna}Tg@HTTP �N!26 ��G�@~obIGUI"%�IPGS�r� H863 qb�!�07r�!�34 �r�84 �\so`! Qx`CC3� Fb�21�!969 rb!51 ���!S53R% 1!s3!���~�.p"9js V{ATFUJ775"���pLR6^RP�WS�MjUCTO�@xT5�8 F!80���1X�Y ta3!770 ���885�UOL�  GTSo
�{` L�CM �r| TSS��EfP6 W�\@CPgE `��0VR� �l�QNL"��@00�1 imrb�c3� =�b�0���0�`6� w�b-P- R-��b8n@5EW�b9 �Ґa� ���b�`ׁ~�b2 2000���`3��`4*5�`5 !�c�#$�`7.%�`�8 h605? U�0�@B6E"aRp76� !Pr8 t�a�@�tr2 iB/d�1vp3�vp5 ȂRtr9Σ�a4@-pN�r3 F��r5&0�re`u��r7 ��r�8�U�p9 \h7�38�a�R2D7�"�1f��2&�7<� �3 7iC���4>w5Ip�Or60� C�L�1bEN�4 I�pyL�uP��@N�&-PJ8�N�8NeN�C9 H�r`�E�b7]�|���8�ВࠂG9 2��a`0�q�Ђ5�%U097 �0��@1�0���1� (�q�3 5R ���0���mpU���0�0�7*�H@(q��\P"RB6�q124�b;��@���@�06� x�3 pB�/x�u ��x�6 H606�a1� ��7 6 ���p��b155 ����7>jUU162 ��3 g��4*�65 2e "_��P�4#U1`���B1���`=0'�174 �q���P�E186 R L��P�7 ��P�8&��3 (�90 B�/�s191����@2s02��6 3���A�RU2� d��O2 b2h`��4��b��2�4���19v RQ�2��u2d�Tpt)2� ��H�a2hP�$2�5���!U2�p�p"
�2�p��@5�0-�@��8 @�9��T�X@�� �e5�`rb	26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0@�gqGA���a�52ѐ�Ḳ6�6�0ہ5� ׁ2��84�E��9�EU5@ٰE\�q5hQ`S�2ޖ5�p\w�۲�pJ �4-P��5�p1\t�H�-4��PCH�7j��phiw�@��P�x��?559 ldu� P �D���Q�@�������A �`.��P>��8�g581�"�q58�!�AM۲T�A iC�a589��@�x���F�5 �a��12׀ 0.�1���,�2�����,�!P\h8��Lp ���,�7��6�084�0\��ANRS 0C}A��p��{��sran��FRA�� �Д�е���A%�� �ѹ�Ҍ�����(�� ��Ќ���З���������ь����$�G��1��ը��������� xS�`�q�  �����`6�4��M��iC/50T-H������*��)p46��� C��xN����m75s֐�� Sp��b46���v����ГM-7�1?�7�З����4A2������C��-��F��70�r�E��/h����O$��rlD���c7c7C� q��Ѕ���L��/���2\imm7c7�g������`���(��e�����"� �������a r��&c�T,�Ѿ�"��,��� ��x�Ex�m7�7t����k���5������)�iC��-HS-� B
_� >���+�Т�7U�]P���Mh7�s��a7������-9?�?/260L_������Q�������]�9pA/@���q�S�х��^�h621��c��92������.�)92c0�g$�@������)$��5$���pcylH"O"
�21�8��t?�350� ���p��$�
�� F�350!���0�x�9�U/0\m9��M9A3��4%�� s��3M$��X%u<���"him98J3����� i d�"m4~��103p�� ����h�794̂�&R���H �0����\���g�5A U��՜��0���*2� �00��#06�а�Ճ�է!07{r  ��������kЙ@�����EP�#�������?��#!�;&0s7\;!�B1P��@�A��/ЁCBׂ2�!��:/��?�ҽCD25�L����0�"l�2BL
#��B��\20�2_�r�re� ��X��1��N����A@��z��`C�pU��`��04��Dy	A�\�`fQ��s�U���\�5  ��� p�^P��<$85���+P=�ab1l��1LT��lA8�!uDnE(�.20T��J�1 e�bH85���b�Ռ�5[�16Bs��������d2��x��m6t!`Q����b�ˀ���b#�(�6iB ;S�p�!��3� ���b�s��-`�_�W80�_����6I	$�X5�1�U85��R�p6S����/�/+q�!@�q��`�6o��5m[o)�m6sW��Q�|�?��set06p h��3%H�5��10p$@����g/�JrH��?  ��A��856����F�� ���p/2��h�܅�✐)�5��̑v�𘜐(��m6��Y�H�ѝ̑m�6�Ҝ��ae6�DM����-S�+��H2�����Ҽ� � �r̑��✐��l���p1���F����2�\t6h T6H����Ҝ�'Vl ���ᜐ�V7ᜐ/�(���;3A7��p ~S��������4�`堜��V���!3��2��PM[��%ܖO�chn��vel5���8�Vq���_arp#���̑�.���2l_h�emq$�.�'�6415���5���?����F�����5g�L�ј�[���1��𙋹1<����M7NU�Р���eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h������ u���㜐��ZS0�!ܑ4���M-����S�$̑�ք �� 0���<�����07shJ�H�v�À�sF� �S*󜐳���̑���vl�3�A�T�#��Q�0��Te��q�pr����T@75j�5�dd�̑ 1�(UL�&�(�,���0��\�?���̑�a�� xSP���a�eD�w�2��(�	�2�C��A/���\�+p�<����21 (ܱ�CL S����B̺@��7F���?�<�lơ1L����c� ���u19�0����e/q���O���9�K��r9 (��,�Rs�ז�5�<G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O���M1!41w���2T@� _std��G�y�� �ң�H� jdgm����w0\� �1L� ��	�P�~�W*�b���t 5������3�,���E{���d���L��5\L��3�L�|#~���~!���4�#��O����h�L6A�������a2璥���44������[6\j4s ��·���#��ol�E"w�8Pk�����?0x j�H1�1Rr�>��]�2a�2Aw�P ��	2��|41�8��ˡ��@{� �%�A<��� +� ?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R�� ˑb�W���Fs���) �ѐ�!���a�1�����5��16�16C���C����0\imBQ��d����b��\Be5�-���DiL����O�_�<ѠPEtL �E�RH�ZǠPgω�am1l��u���̑�b@�<����<�$�T� ̑�F����Ȋ�DpbĜ�X"��hr��pĻ ���^P��9��0\� j971\�kckrcfJ�F�s�����c��e "CTME�r���ɛ�|�a�`main.[�8�g�`run}�_vc�#0�w�1Oܕ�_u����bctme���Ӧ�`ܑ�j73�5�- KARE�L Use {�U���J��1���p� Ȗ�9�B@���L�9��7j[�atk208 "K��(Kя��\��9��a���̹����cKRC4�a�o ��kc�qJ� &s�����Grſ�fs�D��:y��s�ˑ1X\�j|хrdtB�, L��`.v�q�� �spǑIf�Wfj52��TKQuto Seut��J� H5K7536(�932���-91�58(�9�BA��1(�74O,A$�(TCP Ak���/�)Y� �\tpqtool.v���v���! con�re;a#�Cont�rol Re�b{le��CNRE(� T�<�4�2���D�)���NS�552��q(g�� (򭂯4X�cOux~�\sfuts�UTS`�i�栜���At�棂��? 6�T�!�SA OO+D6���������,!��6c+� igt�t6i��I0�T�W8 ���la��vo58�o�bFå򬡯i��Xh��!Xk�0Y!8�\m6e�!6EC���v��6���������<16�A���A�6s����U�g�T|�,����r1�qR����Z4�T�����,#�eZp)g����<ONO0���uJ��tCR;��F<�a� xSP�f���prdsuchk� �1��2&&?���t��*D%$�r(�✑ �娟:r��'�s�qO��<scrc�C�\At�trldJ"o��\�V����Pay�lo�nfirm�l�!�87��7��A�3ad�! �?@ވI�?plQ��3���3"�q��x pl��`���d7��l�calC�uDu���;���mov�����initX�:s8O��a8�r4 ��r67A4|��e Genera#tiڲ���7g2q$g R� (S�h��c ,|�bE��$Ԓ\�:�"���4��4�4�. sg��5�F$d6"�e;Qp "SHA�P�TQ ngcr pGC�a(�&"� ���"GDA¶��r�6�"aW�/�$d�ataX:s�"tp�ad��[q�%tput;a__O7;a�o8�1�yl+s�r�?�:�#$�?�5x�?�:c O�:Ay O�:�IO�s`O%g�qǒ�?�@0\ۜ�"o�j92;!�Pp�l.Collis�QSkip#��@5� �@J��D��@\ވ�C(@X�7��7�|s}2��ptcls�#LS�DU�k?�\_� ets�`�< �\�Q��@���`dcKLqQ�FC;��J,όn��` (��4eN����T�{���' j(�c�����/IӸaȁ<��̠H������зa�e\mcc�lmt "CLM��/��� mate\v��lmpALM�?>p7qmc?�����2vm�q��%�3s��_�sv90�_x_msu�2L^v_� K�o��{in�8(3r<�c_logr��r�trcW� �v_3�~yc��d�<�ste��der$c;Ce� Fiρ��R��Q�?�l�enter߄|��(�Sd��1�TX�+fZK�r�a99sQ9+��5�r\tq\� _"FNDR����STDn$�LANG�Pgui��D⠓�S������csp�!ğ֙uf䟀ҝ�s����$�����e +�=����������������w�H�r\fn�_�ϣ��$`x�tcp�ma��- TCP������R638 aR�Ҡ��38��M7p,���Ӡ�$Ӡ��8p0Р�VS,�>�tk��99�a��B3���P�զԠ��D�2�����UI��t���hqB���8���������p���re8�ȿ��exe@4π��B���e38�ԡG�r�mpWXφ�var @�φ�3N�����v�x�!ҡ��q�R�BT $cOP�TN ask E�0��1�R MAS�0�H593/�96g H50�i�480ԅ5�H0��m�Q�K(��7�0�g�Pl�h�0ԧ�2�ORDP���@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`am��b��7�.f���u�d��r��splayD�E���1wПUPDT Ub��8o87 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60�q��B����qs�can��B���aAd@�������q`� �䗣�#��К�`2�� vlv��Ù�$�0>�b���! S���Easy/К�Ut�il��룙�511# J�����R7 ���Nor֠��inc�),<6Q�� �`c��"4�[���986(FVRx So����q�nd6����P��4� a\ (��
  ������"�d��K�bdZ����men7���- Me`tyFњ�Fb��0�TUa�577?i3R��\�5�au?��!� n����f������l\m�h�Ц�űE|h#mn�	��<\O�$��e�1�� l!���y��Ù�\|p�����B���Ћmh �@��:.aG!�� �/�t�55�6�!X��l�.us��Y/k)eOnsubL���eK�h�� �B\1;5g?�y?�?�?D��?*rmx�p�?Ktbox O�2K|?�G��C?A%das���?1ӛ#� � TR��/��P�4B�`�U@�P�V�P"�Q�P0�U �PO��P�"�T3�U�P �f�Pk"�2}�4�T�P �f�P2�"�Q5�S�Q@���R?Ă�Q3t.�PF׀al��P+O�n�P517��IN0a���Q(}g��PES	Tf3ua�PB�l�i�g�h�6�aq��P �� xS��` � n�0mbump�P�Q969g�69�Qq��P0�baAp�@>Q� BOX��,�>vche�s�>ve�tu㒣=wffse�3���]�;u`aW��:zol�sm<u�b�a-��]D�K�ib�Q�c����Q<twaǂ �tp�Q҄Taror Recov�br�O�P�642�����a�q��a⁠QErǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>��pjot��PXc��C��1�adb -�ail���nag���b�QR629�a�Q��b�P�  �
 � �P��$$CL~[q ����������$�PS?_DIGIT���"�!�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��������*璬1:P�RODUCT�Q0�\PGSTK�bV�,n�99�\����$FEAT_INDEX���~�� �搠ILECOM�P ;��)���"��SETUPo2 <��?�  N !��_AP2BCK �1=�  �)}6/E+%,/i/��W/�/~+/�/O/ �/s/�/?�/>?�/b? t??�?'?�?�?]?�? �?O(O�?LO�?pO�? }O�O5O�OYO�O _�O $_�OH_Z_�O~__�_ �_C_�_g_�_�_	o2o �_Vo�_zo�oo�o?o �o�ouo
�o.@�o d�o���M� q���<��`�r� ���%���̏[���� ���!�J�ُn����� ��3�ȟW������"� ��F�X��|����/� ��֯e������0��� T��x������=�ҿ �s�ϗ�,ϻ�9�b�t� P/ 2) *.VRiϳ�!�*���������Ɲ�PC�7�!�F'R6:"�c��χ��T��߽�Lը����x���*.F���>� �	N�,�k�x�ߏ��STM �⠸���Qа���!��iPendant? Panel���H��F���4������GIF�������pu����JPG&�P��<����	�PANEL1.D	T��������2�Y�G��
3w�����//�
4�a/��O///�/�
TP�EINS.XML�/���\�/�/�!�Custom T?oolbar?��PASSWOR�D/�FRS:�\R?? %Pa�ssword Config�?��? k?�?OH�6O�?ZOlO �?�OO�O�OUO�OyO _�O�OD_�Oh_�Oa_ �_-_�_Q_�_�_�_o �_@oRo�_voo�o)o ;o�o_o�o�o�o*�o N�or��7� �m��&���\� ����y���E�ڏi� �����4�ÏX�j��� �����A�S��w�� ���B�џf������� +���O��������� >�ͯ߯t����'��� ο]�򿁿�(Ϸ�L� ۿpς�Ϧ�5���Y� k� ߏ�$߳��Z��� ~�ߢߴ�C���g��� ��2���V����ߌ� ��?����u�
��� .�@���d������)� ��M���q�����< ��5r�%�� [�&�J� n��3�W� ��"/�F/X/�|/ /�/�/A/�/e/�/�/ �/0?�/T?�/M?�?? �?=?�?�?s?O�?,O >O�?bO�?�OO'O�O KO�OoO�O_�O:_�O ^_p_�O�_#_�_�_Y_��_}_o�_�_Ho)f��$FILE_DG�BCK 1=���5`��� ( �)
S�UMMARY.DyGRo�\MD:�o��o
`Diag� Summary��o�Z
CONSLOG�o�o�a
J�a�ConsoleO logK�[�`�MEMCHECK�@'�o�^qMe�mory Dat�a��W�)>�qHADOW����P��sShad�ow Chang�esS�-c-��)	FTP=��9�����w`qmmen�t TBD׏�W0�<�)ETHERNET̏�^�q��Z��aEther�net bpfiguration[���P��DCSVRF�ˏ��Ïܟ�q%��� verify� allߟ-c1P{Y���DIFFԟp��̟a��p%��diffc���q���1X�?�Q�� �����X��CH�GD��¯ԯi��px��� ���2`�G�Y��� ��� �GAD��ʿܿq��p���Ϥ�FY3h�O�aώ�� ��(�GAD������y��p�����0�UPDAT�ES.�Ц��[FORS:\�����a�Updates �List���kPS�RBWLD.CM�.��\��B��_pP�S_ROBOWEL���_����o��,o !�3���W���{�
�t� ��@���d�����/ ��Se����� N�r� =� a�r�&�J� ��/�9/K/�o/ ��/"/�/�/X/�/|/ �/#?�/G?�/k?}?? �?0?�?�?f?�?�?O �?OUO�?yOO�O�O >O�ObO�O	_�O-_�O Q_c_�O�__�_:_�_ �_p_o�_o;o�__o �_�o�o$o�oHo�o�o ~o�o7�o0m�o � ��V�z� !��E��i�{�
��� .�ÏR���������� .�S��w������<� џ`������+���O� ޟH������8���߯�n����$FIL�E_��PR����������� �MDONL�Y 1=4�� 
 ���w�į�� 诨�ѿ�������+� ��O�޿sυ�ϩ�8� ����n�ߒ�'߶�4� ]��ρ�ߥ߷�F��� j�����5���Y�k� �ߏ���B�����x� ���1�C���g���� ��,���P����������?��Lu�VI�SBCKR�<�a��*.VD|�4 OFR:\��4 �Vision VD file�  :LbpZ�# ��Y�}/$/� H/�l/�/�/1/�/ �/�/�/�/ ?�/1?V? �/z?	?�?�???�?c? �?�?�?.O�?ROdOO �OO�O;O�O�OqO_ �O*_<_�O`_�O�__�%_�_�MR_GR�P 1>4�L~�UC4  B�P�	 ]�ol`��*u����RHB ��2 ���� ��� ���He�Y�Q`ork bIh�oJd�o�Sc�o��oMS��O|�N$L���F�{5U�aT�˱�o��o^`��C%�љCre�*~��G86X=5���}?�]�A��\blq>����A�W�xq}E�?� F@ �r�d��a}J��NJk��H9�Hu���F!��IP��sX~�`�.9��<9�8�96C'6<�,6\b~AL�opB*�~Bo�$A�~/A�J4B2v ����A�_�B<�`�AF��<�׃����,.��PA�����|�ݏx����%���p�A6Β@U��{�v� a�������П����ߟ���<�'�hzBH�P �a`�Q�H��,�qK���ï�T
�6�PJ��PJ�`Ɂ��o�o)�B��P<5���@�33@����4�m�,�@UUU�U�~w�>u.�?!x�^��ֿ����3��=[z��=�̽=V6�<�=�=��=$q��~��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�O� Cϫo4z��P��P'�6��_V� m �o��To��xo�ߜo�� ����A�,�e�P�b� ������������ �=�(�a�L���p��� ������.�������* ��N9r]��� �����8# \nY�}���� ���/ԭ//A/� e/P/�/p/�/�/�/�/ �/?�/+??;?a?L? �?p?�?�?�?�?�?�? �?'OOKO6OoO�OH� �Ol��ߐߢ��O�� _ ��G_bOk_V_�_z_�_ �_�_�_�_o�_1oo Uo@oyodovo�o�o�o �o�o�oN u������ ���;�&�_�J��� n�������ݏȏ�� %�7�I�[�"/�描� ����ٟ�������3� �W�B�{�f������� կ�������A�,� e�P�b��������O�O �O��O�OL�_p� :_�����Ϧ������ ��'��7�]�H߁�l� �ߐ��ߴ�������#� �G�2�k�2��Vw� ����������1�� U�@�R���v������� ������-Q� u���r��6� �)M4q\ n������/ �#/I/4/m/X/�/|/ �/�/�/�/�/?ֿ� B?�f?0�BϜ?f��? ���/�?�?�?/OOSO >OwObO�O�O�O�O�O �O�O__=_(_a_L_ ^_�_�_�_���_��o �_o9o$o]oHo�olo �o�o�o�o�o�o�o# G2kV{�h �������C� .�g�y�`��������� �Џ���?�*�c� N���r��������̟ ��)��M�_�&?H? ���?���?�?�?��� �?@�I�4�m�X�j��� ��ǿ���ֿ���� E�0�i�Tύ�xϱϜ� ��������_,��_S� ��w�b߇߭ߘ��߼� ������=�(�:�s� ^��������� �'�9� �]�o���� ~������������� 5 YDV�z� �����1 U@yd��v�� ���/Я*/��
/� u/��/�/�/�/�/�/ �/??;?&?_?J?�? n?�?�?�?�?�?O�? %OOIO4O"�|OBO�O >O�O�O�O�O�O!__ E_0_i_T_�_x_�_�_ �_�_�_o�_/o��?o eowo�oP��oo�o�o �o�o+=$aL �p������ �'��K�6�o�Z�� ����ɏ��폴� � �D�/ /z�D/��h/ ş���ԟ���1�� U�@�R���v�����ӯ ������-��Q�<� u�`���`O�O�O��� ޿��;�&�_�J�o� �πϹϤ�������� %��"�[�F��Fo�� �����ߠo��d�!�� �W�>�{�b���� ����������A�,� >�w�b����������������=��$�FNO ����\��
F0l q  oFLAG>�(R�RM_CHKTY/P  ] ��d ��] ��OM�� _MIN� 	����� �  X�T SSB_CFG� ?\ �����OTP_DEF�_OW  	�|�,IRCOM� �>�$GENOV�RD_DO���<�lTHR� dz�dq_ENB]� qRAVC_?GRP 1@�I X(/ %/7/ /[/B//�/x/�/�/ �/�/�/?�/3??C? i?P?�?t?�?�?�?�? �?OOOAO(OeOLO�^O�OoROU�F\\� �,�|B,�8�?����O�O�O	__  D��UPE_�Hy_�\@@m_B�=�vR/��I\�O�SMT�G����
�oo+l��$HOSTC�19H�I� ��zM�SM�l[�bo�	127.�0�`1�o  e �o�o�o#z�oF�Xj|�l60s	a�nonymous�������-(ao�&�&��o� x��o������ҏ�3 ��,�>�a�O���� ������Ο�U%�7�I� �]����f�x����� ���ү����+�i� {�P�b�t�������� ����S�(�:�L� ^ϭ�oϔϦϸ���� ��=��$�6�H�Zߩ� ��Ϳs���������� � �2���V�h�z�� �߰���������
�� k�}ߏߡߣ���߬� ��������C�*< Nq�_����� �-�?�Q�c�eJ�� n������ �/"/E�X/j/|/ �/�/�%'/? [0?B?T?f?x?��? �?�?�?�??E/W/,O�>OPObO�KDaENT� 1I�K P!\�?�O  �P�O �O�O�O�O#_�OG_
_ S_._|_�_d_�_�_�_ �_o�_1o�_ogo*o �oNo�oro�o�o�o	 �o-�oQu8n �������� #��L�q�4���X��� |�ݏ���ď֏7����[���B�QUICC0��h�z�۟��A1ܟ��ʟ+���2,����{�!ROU�TER|�X�j�˯!?PCJOG̯���!192.168.0.10���}GNAME !��J!ROBOT��vNS_CFG �1H�I ��Auto-s�tarted�$FTP�/���/�? ޿#?��&�8�JϏ? nπϒϤ�ǿ��[���`���"�4�G�#��� ��������������� �����&�8�J�\�n� ������������� �/�/�/F���j��ߎ� ������������ 0S�T��x��� ��!�3��G,{� Pbt��C�� ��/�:/L/^/ p/�/���	/�/ =?$?6?H?Z?)/~? �?�?�?�/�?k?�?O  O2ODO�/�/�/�/�? �O�/�O�O�O
__�? @_R_d_v_�_�O-_�_ �_�_�_oUOgOyO�O �_ro�O�o�o�o�o�o �_&8Jmo�o �����o)o;o MoO!��oX�j�|��� ��oď֏����/����B�T�f�x���^�S�T_ERR J�;�����PDUSI�Z  ��^P�����>ٕWRD �?z���  �guest ���+�=�O�a�s�*��SCDMNGRPw 2Kz�Ð���۠\��K��� 	P01.�14 8�q  � y��B    ;�����{ �����������������������~ �ǟI�4�m�X��|��  i�  �  
����� ����+��������
����l�.x��
��"�l�ڲ۰s��d�������_G�ROU��L�� e��	��۠07K�QUPD  ����PČ�TYg������TTP_A�UTH 1M��� <!iPen'dan���<�_��!KAREL�:*�����KC�%�5�G��VISION SETZ���|��Ҽߪ��� ������
�W�.�@����d�v���CTRL� N�������
��FFF9E�3���FRS:DEFAULT��FANUC �Web Server�
������q�������������W�R_CONFIGw O�� ����IDL_CPU�_PC"��B���= �BH#MI�N.�BGNR_�IO��� ���% N�PT_SIM_D�Os}TPMO_DNTOLs �_PRTY�=!OLNK 1P���'9K]|o�MASTEr ������O_CFG���UO����C�YCLE���_?ASG 1Q���
 q2/D/V/h/ z/�/�/�/�/�/�/�/p
??y"NUM����Q�IPCH���£RTRY_�CN"�u���SC�RN������ ���R����?���$J23_D_SP_EN������0OBPROC��3��JOGV�1�S_�@��8��?�';ZO'??0CP�OSREO�KANJI_�Ϡu�A$#��3T ���E�O�ECL_LM B2e?��@EYLOGGI�N�������L�ANGUAGE Y_�=� }Q���LG�2U������ �x�����PZC � �'0������MC:\RSCH\00\˝�LN_DISP V�������T�OC�4Dz\=�#�Q�?PBOOK W+��o���o�o���Xi�o�o�o�o�o~}	x(y��	ne�i�ekEl�G_BUFF 1%X���}2�� ��Ӣ������ '�T�K�]��������� ��ɏۏ���#�P���ËqDCS Z>xm =���%|d�1h`���ʟܟ�g�I�O 1[+ �?'����'�7�I�[� o��������ǯٯ� ���!�3�G�W�i�{�@������ÿ׿�El /TM  ��d��#� 5�G�Y�k�}Ϗϡϳ� ����������1�C߀U�g�yߋߝ߈t�S�EV�0m�TYP�� ��$�}��ARS"�(_�s�2F�L 1\��0� ��������������5�TP<P���>DmNGNAM�4�U��f�UPS`GI�5�A�5s�_LO{AD@G %j{%@_MOV�u�����MAXUALRMB7�P8��y��D�3�0]&q��Ca]s�3�~�� 8@=@]^+ طv	��+V0+�P�A5dƋr���U ������E (iTy���� ���/ /A/,/Q/ w/b/�/~/�/�/�/�/ �/??)?O?:?s?V? �?�?�?�?�?�?�?O 'OOKO.OoOZOlO�O �O�O�O�O�O�O#__ G_2_D_}_`_�_�_�_ �_�_�_�_o
ooUo 8oyodo�o�o�o�o�o��o�o�o-��D_L?DXDISA^��� �MEMO_AP�X�E ?��
 �0y�����������ISCw 1_�� � O����W�i����� Ə�����}��ߏD� /�h�z�a�������� ������@���O� a�5������������ u��ׯ<�'�`�r�Y� �����y�޿�ۿ� ��8Ϲ�G�Y�-ϒ�}� �ϝ�����m�����4���X�j�#�_MST�R `��}�SC/D 1as}�R��� N��������8�#�5� n�Y��}������� �����4��X�C�|� g��������������� 	B-Rxc� ������ >)bM�q�� ���/�(//L/ 7/p/[/m/�/�/�/�/ �/�/?�/"?H?3?l?�W?�?{?�?�?�?n�MKCFG b����?��LTARMu_�2cRuB� �3WpTNBpM�ETPUOp�2�����NDSP_CMNTnE@F�E��' d���N�2A��O�D�EPOSCF��G�NPSTOL� 1e-�4@�<#�
;Q�1;UK_YW 7_Y_[_m_�_�_�_�_ �_�_o�_oQo3oEo��oio{o�o�a�ASI�NG_CHK  y�MAqODAQ2C�fO�7J�eDEV� 	Rz	MC}:'|HSIZEn@�����eTASK �%<z%$123456789 ���u�gTRIG 1]g�� l<u%����3���>svvY�Paq��kEM_I�NF 1h9G� `)AT&FV0E0(����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ ߏP��t�������]� ί�����(�۟� ^��#�5�����k�ܿ � ϻ�ů6��Z�A� ~ϐ�C���g�y����� ���2�i�C�h�ό� G߰��ߩ��ߙϫ�� ������d�v�)ߚ��� ��y��������<� N��r�%�7�I�[��� ���9�&��J�[�g��>ONIwTOR�@G ?;{�   	EX�EC1�3�2�3��4�5��p�7*�8�9�3�n� R�R�RR RR(R4R@�RLR2Y2e2�q2}2�2�2��2�2�2�3�Y3e3��aR_�GRP_SV 1�it��q(�a?��ڿ
�3�8���1��۵M�O~q_DCd~�1P�L_NAME �!<u� �!D�efault P�ersonali�ty (from� FD) �4RR�2k! 1j)TE�X)TH��!�AX d�?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�Ox2-?�O�O�O__@0_B_T_f_x_�b<�O �_�_�_�_�_�_o o�2oDoVoho&xRj" �1o�)&0\�b,� �9��b�a �@D�  �a?�ľc�a?�`�a�aA'�6�ew;�	�l�b	 ��xJp���`�`	p �<w �(p� �.r�� K�K ���K=*�J����J���JV�`�kq`q�P�x��|5p@j�@T;;f�r�f�q�a�crs�I�� چ�p���p�r� h}��3��´  Æ�>��ph�`z���꜖"�3Jm�q� H�N���ac���dw�� ~ �  P� �Q� �� |  �а�m�Əi}	'�� � �I�� �  ��ވ�:�È�È�=���(�ts�a	����I  �n @H�i~�ab�ӋB�b�w��urN0��  'Ж�q�p�@2��@���X�r�q5�C�pC0C�@ C���=�`
�A1q   @B�UV~X�
nwB0"h�A��p�ӊ�p�`���aDz���֏����Я	�pv�( �� -���I��-�=��A�a���e_q�`�p �?�ff ��m��>� ����Ƽ�uq1!ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`�5p<
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC��������#/*/c/N/�wi�����v/C�`� CHs/`
=$�p��<!�!��ܼ�'��3A�A�AR�1AO�^?�$��?��5p±�
=ç>�����3�W
=�#��]�;e�׬a@�����{�����<�>(��B�u���=B0�������	R��zH�F��G���G���H�U`E����C�+��}I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*O ONO9OrO]O�O�O�O �O�O�O�O_�O8_#_ \_G_�_�_}_�_�_�_ �_�_�_"oooXoCo |ogo�o�o�o�o�o�o �o	B-fQ� u������� ,��P�b�M���q��� ��Ώ���ݏ�(�� L�7�p�[������ʟ ���ٟ���6�!�Z��E�W���#1($1�ٙ9�K���ĥ%�����ƯS�3��8���S�4Mgqs��,�IB+8��J��a���{�d�d�����ȿ��쿔ڼ%P8�P�= :GϚ�S�6�h�z���R�Ϯ����������  %�� ��h� Vߌ�z߰�&�g�/9�$�������7�����A�S�e�w�   ������������̿2 F�$�&Gb��������!C���@���8������F� Dz�N�� F�P �D�������)#�B�'9K]o#?_���@@v
$�8�8��8�.
 v��� !3EWi{�����:� ���ۨ�1��$M�SKCFMAP � ���� ���(.�ONREL  ��!9��EXC/FENBE'
#7%�^!FNCe/W$JO�GOVLIME'dtO S"d�KEYE'u�%�RUN�,��%�SFSP�DTY0g&P%9#S�IGNE/W$T1M�OT�/T!�_C�E_GRP 1p��#\x��?p� �?�?�?�?�?O�? OBO�?fOO[O�OSO �O�O�O�O�O_,_�O P__I_�_=_�_�_�_ �_�_oo�_:o��TCOM_CFG 1q	-�vo�o��o
Va_ARC_�b"�p)UAP_�CPL�ot$NOCHECK ?	+ �x�% 7I[m���������!�.+N�O_WAIT_L� 7%S2NT^ar�	+�s�_ERR�_12s	)9��  ,ȍޏ��x����&��dT_MO��t>��, �k*oq��9�PARAM��u	+��a�ß'g�{�� =?�345?678901�� ,��K�]�9�i�����`��ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDS�P�c#6p(OFFSET_CART�oη�DISƿ��PE?N_FILE尨!��ai��`OPTIO�N_IO�/��PW�ORK ve7�s# ��Vż�8�  � �<�p�4�p�	 ���p��<�� �C�_DSBL  ���P#��ϸ�R�IENTTOD �?�C�� !=#���UT_SIM_ED$�"���V��?LCT w}���6��a[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ����s��ڐH(���H3k7HSM�5G�22G���Gp
͜�'fc�/-,ڐCR�	>�D!�M#{Z/���3�����4 y H "�c/u/�/0�B_����j�c��t�!�/ �/�"t32����/�6  ��P�%�Q%��%�|T���S62�q?'e	'� �� �2I� �  ��+==��ͳ?�;	�h�	�0�I  �n @�2�.��O�v;��ٟ?&gN �[OaA''�uD@!� Cb@C�@F#H!�/�Oz�O sb
�Ab@*�@�@��@�e0@Bb@QA�0Yv:G �13Uwz$o�V_�/z_e_�_�_	���( �� -�2�1�1ta�Ua�"c���:A����. ? �?�ff���[o"o�_U�`oX�0A�8���o�j>�1  	Po�V(���eF0�f��Y���L�?�嚫�xb0@<
6�b<߈;܍��<�ê<� <�&�,/a�A�;r�@Ov0P?f7ff?�0?&ip�T�@�.{r�J<?�`�u#	�Bdq t�Yc�a�Mw� Bo��7�"�[�F�� j�������ُ�� ��3����,���(��E�� E��3G+� F��a��ҟ �����,��P�;���B�pAZ�>��B ��6�<OίD���P�� t�=���a�s�����6j��h��7o��>��S��O����όFϑ�A�a�_��C�3Ϙ�/�%?��?�A��������#	Ę�a�P �N||CH����Ŀ������@I��_�'�3A��A�AR1AO��^?�$�?������±
=���>����3�?W
=�#� U���e���B��@���{����<������(�B�u���=B0������	�b��H�F�G����G��H�U�`E���C�+���I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻���������  �9�$�]�H�Z���~� ������������#5  YD}h��� ����
C. gR������ �	/�-//*/c/N/ �/r/�/�/�/�/�/? �/)??M?8?q?\?�? �?�?�?�?�?�?O�? 7O"O[OmOXO�O|O�O �O�O�O�O�O�O3_Q�(������b�y�gUU��W_<i_2�3�8��_�_2�4Mgs�_�_�R�IB+�_�_�a���{�miGo@5okoYo�o}l��P'r	P�nܡݯ�o=_�o0�_�[R?Q`�u���  �p���o��/��S� �z
uүܠ�������ڱ�����������  /�M�w�e�𛟉����l2 F;�$��Gb��t�a�a�`�p�S�C�y��@p�5�G�Y�۠F�� Dz�� F�P D��]����پ��ʯܯ�� ��~�?���@U@�?�K�K�꺡K���
  �|�������Ŀֿ� ����0�B�T�fϽ��V� ���{��1���$PARAM�_MENU ?�3�� � DEFP�ULSEr�	W�AITTMOUT���RCV�� �SHELL_W�RK.$CUR_oSTYL��	��OPT��PTB�4�.�C�R_DECSN���e��ߑ� ������������!�3�\�W�i�{���U�SE_PROG �%��%�����C�CR���e����_HOST !��#!��:���T�`��V��/�X����_�TIME��^�� � ��GDEBU�G\�˴�GINP?_FLMSK����qTfp����PGA e ����)CH��^��TYPE�����������  -?hcu� ������// @/;/M/_/�/�/�/�/ �/�/�/�/??%?7?�`?��WORD ?}	=	RSfu_	PNSU��2JOK�DRTE�y�]TRACEC�TL 1x3��� �`. �&�`�`�>�6D/T Qy3�%@�0�D � �c7�a:@V�@BR�2ODOVOhO�zO�O�O�H�C�H�O�O�H
�B *TTT�L^� RTTT��L�L� R!T� �U�E�_�_�_�_�_�_ o o2oDoVohozo�o �o�o�o�o�o�o
 .@Rdv��� ������*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�.Iv� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��j� ���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�o�o�o�o ��o0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ����������*��$PGTR�ACELEN  �)�  ���(��>�_U�P z���2m�u�Y�n�>�_CFG {m�SW�(�n����PКӂ�DEFSP/D |��'�P���>�IN��TR�L }��(�8�����PE_CON�FI��~m���mњ��ղ�L�ID����=�G�RP 1��W���)�A ����&ff(�A+33�D�� D]� ?CÀ A@1����(�d�Ԭ��0�0�?� 	 1��8�֚��� ´�����B�9����O��9�s�(�>�T?��
5�������� �=��=#�
 ����P;t_�������� G Dz (�
 H�X~i��� ���/�/D///�h/S/�/��
V7�.10beta1���  A��E�"ӻ�A �(�� ?!G��!>����"����!{���!BQ��!�A\� �!���!2p
����Ț/8?J?\?�n?};� ���/� �/�?}/�?�?OO:O %O7OpO[O�OO�O�O �O�O�O_�O6_!_Z_ E_~_i_�_�_�_�_�_ �_'o2o�_VoAoSo �owo�o�o�o�o�o�o .R=v1�/�#F@ �y�}� �{m��y=��1�'� O�a��?�?�?������ ߏʏ��'��K�6� H���l�����ɟ��� ؟�#��G�2�k�V� ��z��������o� �ίC�.�g�R�d��� �������п	���-� ?�*�cώ���Ϯ� �����B�;�f� x�������DϹ��߶� �������7�"�[�F� X��|��������� ��!�3��W�B�{�f� �������� ����� /S>wbt� �����= OzόϾψ����� �� /.�'/R�d�v� �߁/0�/�/�/�/�/ �/�/#??G?2?k?V? h?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O���O�O�O__ ?_*_c_N_�_r_�_�_ �_�_�_o�_)oTf x�to���/�o />/P/b/t/m o�|����� ��3��W�B�{�f� x�����Տ������ �A�S�>�w�b����O ��џ������+�� O�:�s�^�������ͯ ���ܯ�@oRodo�o `��o�o�o��ƿ�o� ��*<N�Y��}� hϡό��ϰ������� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�c�N�ﲟ��� l��������;�&� _�J���n��������� ��,�>�P�:L�� ���������� (�:�3��0iT� x�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?a?s?��?�?X?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O *\&_8_r����_�_��$PLI�D_KNOW_M�  ��� Q�TSV ���P��?o"o4o�OXo�CoUo�o R�SM_?GRP 1��Z'U0{`�@�`uf
�e�`
�5� �gpk 'Pe] o�������X���SMR�c��m1T�EyQ}? yR�� ��������폯���ӏ �G�!��-������� ����韫���ϟ�C� ��)������������寧���QST�a1W 1��)���P;0� A 4��E 2�D�V�h�������߿ ¿Կ���9��.�o� R�d�vψ��ϬϾ�����2�0� Q�	<3��3�/�A�S߂�4l�~ߐߢ��5 ���������6
��.�@��7Y�k�}���8��������M_AD  )���PARNUM  !�}o+��WSCHE� S�
��pf���S��UPDf��x��_CM�P_�`H�� �'��UER_CHK-���ZE*<�RSr��_�Q_MO�G���_�X�_R/ES_G��!��� D�>1bU� y�����/�	/����+/� k�H/g/l/��Ї/�/ �/�	��/�/�/�X� ?$?)?���D?c?h?�����?�?�?�V �1��U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_�INRr�J�b�Ud�2FMASS?O Z�SGMN>OqCMON�_QUEUE a��U�V P~P X�N$ UhN�FV�@�END�A��IEX1E�O�E��BE�@�O>�COPTIO�G���@PROGRAM7 %�J%�@�?����BTASK_I�G�6^OCFG ኤOz��_�PDATuA�c��[@Ц2=�DoVohozo�j2o �o�o�o�o�o)x;M jINFO[��m��D��� �����1�C�U� g�y���������ӏ����	�dwpt�l �)�QE DIT ��_i��^WERF�LX	C�RGADoJ �tZA���¿�?נʕFA��IOORITY�GW���MPDSPNQ�����U�GD��OTO�E@1�X� (/!AF:@E� c�~Ч!tcpn�>��!ud����!icm���?<��XY_�Q�X�=��Q)� *�1�5��P��]�@�L� ��p��������ʿ� �+�=�$�a�Hυϗ�=*��PORT)QH���P�E��_C?ARTREPPX�>�SKSTA�H�
�SSAV�@�tZ	�2500H86A3���_x�
�'��X�@�swPtS��x�ߧ���URGE�@�B��x	WF��DO�F"[W\��������WRUP_DEL�AY �X���RO_HOTqX	B%��c���R_NORM�ALq^R��v�SE�MI�����9�QS�KIP'��tUr�x 	7�1�1�� X�j�|�?�tU������ ��������$J \n4����� ���4FX |j������ �/0/B//R/x/f/�/�/�/tU�$RCgVTM$��D�� �DCR'������!?�0�Cw���C��>��+=_��:��+:��ss������(Z�:��o?�� <
6b�<߈;܍��>u.�?!<�&�?h?�?�? �@>��?O O2ODOVO hOzO�O�O�O�O�O�? �O�O__@_+_=_v_ Y_�_�_�?�_�_�_o o*o<oNo`oro�o�o �o�_�o�o�o�o�o 8J-n��_�� �����"�4�F� X�j�U������ď�� �ӏ���B�T�� x���������ҟ��� ��,�>�)�b�M��� ���������ïկ� Y�:�L�^�p������� ��ʿܿ� ����6� !�Z�E�~ϐ�{ϴϗ� ����-�� �2�D�V� h�zߌߞ߰������� ��
���.��R�=�v� ��k��������� �*�<�N�`�r����� �����������& J\?���� ����"4F�Xj|��!GN_�ATC 1�	;� AT&F�V0E0�A�TDP/6/9/�2/9�ATA��,AT%G1%B960��++5;��H�/,�!IO_TY�PE  �%�#�t�REFPOS�1 1�V+ x�u/�n�/j �/
=�/�/�/Q?<?u? ?�?4?�?X?�?�?�+/2 1�V+�/�?��?\O�?�O�?�!3 1�O*O<OvO�O�O|_�OS4 1��O��O�O_�_t_�_+_S5 1�B_T_f_�_�o	oBo�_S6 1��_�_�_5o�o�o�o>UoS7 1�lo~o��o�oH3l�oS8 1�%_����SMASKw 1�V/  
?��M��XNOS/�r�������!MOTE�  n��$��_CFG ����q���"PL_RANG������POWER ������SM�_DRYPRG �%o�%�P��T?ART ��^�UME_PRO-��?����$_EXEC_ENB  ���GSPD��Րݘ���TDB��
�R�M�
�MT_'�T�����OBOT�_NAME �o����OB_O�RD_NUM ?��b!H?863  �կ����PC_TIMEOUT��{ x�S232Ă�1�� L�TEACH PE�NDAN��w���-��Mai�ntenance Cons���s��"���KCL/!Cm��

���t�ҿ� No Us�e-��Ϝ�0�NPqO�򁋁���.�CH_L�������q	��s�MAVAIL������糅��SPACE�1 2��, �j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��ߤ� �ߚ� �2�D���h� ��|��`������ ���� �2�D��h� ��|���`���������y���2����0� B���f�����{���3); M_����� �/� /44F Xj|*/���/�/@�/?(??=?5Q/ c/u/�/�/G?�/�/�?�O�?$OEO,OZO6 n?�?�?�?�?dO�?�? _,_�OA_b_I_w_7�O�O�O�O�O�_�O _(oIoo^oofo�o8�_�_�_�_�_�o o6oEf){����G �o�� ���
M� ���*�<�N�`�r� ������w���o������d.��%�S� e�w�����������Ǐ َ���Θ8�+�=�k� }�������ůׯ͟�� ��%�'�X�K�]��� ������ӿ�����p�#�E�W� `� @�������x�����\�e������ �����R�d߂�8�j� �߾߈ߒߤ������ ����0�r���X�� ����������8�����
�ύ�_MO�DE  �{��S ��{|�2�0�A����3�	S�|)CWORK_{AD��*K�+/R  �{�`� ��� _INTVA�L���d���R_O�PTION� ���H VAT_G�RP 2��up(N�k|��_�� ���/0/B/��h� u/T� }/�/�/�/�/ �/�/?!?�/E?W?i? {?�?�?5?�?�?�?�? �?O/OAOOeOwO�O �O�O�OUO�O�O__ �O=_O_a_s_5_�_�_ �_�_�_�_�_o'o9o �_Iooo�o�oUo�o�o �o�o�o�o5GY k-���u�� ���1�C��g�y� ��M�����ӏ叧�	� �-�?�Q�c������� ��������ǟ��;�M�_����$SC?AN_TIM��_%�}�R �(�#((�<04_d d 	
!D�ʣ���u�/������U��25�����d�A�8�H�g��]	 ���������dd�x��  P����; ��  8� ҿx�!���D��$� M�_�qσϕϧϹ���������ƿv���F�X��/� ;G�ob��pm���t�_Di�Q̡  � l �|�̡ĥ������� !�3�E�W�i�{��� ������������/� A�S�e�]�Ӈ����� ��������); M_q����� ��r���j�T fx������ �//,/>/P/b/t/��/�/�/�/�/�%�/  0��6��!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O*�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo�O�OJ�o�o �o�o�o�o�o 2 DVhz��������
�7?   ;�>�P�b�t������� ��Ǐُ����!�3� E�W�i�{�������ß �ş3�ܟ�� &�8�J�\�n�������������ɯ�����,� �+�	�1234567�8�� 	� =5���f�x�������������
��.� @�R�d�vψϚ�៾� ��������*�<�N� `�r߄߳Ϩߺ����� ����&�8�J�\�n� �ߒ����������� �"�4�F�u�j�|��� ������������ 0_�Tfx��� ����I> Pbt����� ��!/(/:/L/^/ p/�/�/�/�/�/�/�2�/?�#/9?K?�]?�iCz  B}p˚   ��h�2��*�$SCR�_GRP 1�(��U8(�\x�d�@} � ��'�	 �3�1�2�4(1*�&��I3�F1OOXO}m��D�@�0ʛ�)���HUK�LM�-10iA 89�0?�90;��F;�M61C D�:�CTP��1
\&V�1 	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^�o OUO>oPo#G�/����o'o�o�o�o�oB��0�rtAA�0*  @�Bu&"Xw?��ju�bH0{�UzAF@ F�`�r��o���� �+��O�:�s��mBq�rr����������B� ͏b����7�"�[�F� X���|�����ٟğ�� �N���AO�0�B�CU�
L���E�jqBq>33���$G@�@pϯ7 B���G�I�
E�0EL_DEFAULT  �T���E���MIPOWERFL  
E*���7�WFDO� �*��1ERVENT? 1���`(��� L!DUM�_EIP��>��j�!AF_INEx�¿C�!FT�������!o:� ���a�!RP?C_MAINb�D�q�Pϭ�t�VIS}��Cɻ����!TP&��PU�ϫ�d��E��!
PMON_POROXYF߮�e4ߐ���_ߧ�f����!�RDM_SRV��߫�g��)�!R��Iﰴh�u�!
�v�M�ߨ�id���!RLSYNC���>�8���!R3OS��4��4��Y� (�}���J�\������� ������7��[" 4F�j|�����!�Eio�I�CE_KL ?%�� (%SVCPRG1n>����3��3���4�//�5./3/�6V/[/�7~/�/��D$�/�9�/�+�@� �/��#?��K?� �s?� /�?�H/�? �p/�?��/O��/ ;O��/cO�?�O� 9?�O�a?�O��?_ ��?+_��?S_�O {_�)O�_�QO�_� yO�_��Os��� �>o�o}1�o�o�o�o �o�o�o;M8 q\������ ���7�"�[�F�� j�������ُď��� !��E�0�W�{�f��� ��ß���ҟ��� A�,�e�P���t�����࿯�ί�y_DE�V ���MC:�@`.!�OUT��2�~�REC 1�`e��j� �� 	 �����˿���8ڿ��
 �`e�� �6�N�<�r�`ϖτ� ���Ϯ�������&�� J�8�n߀�bߤߒ��� ��������"��2�X� F�|�j�������� ������.�T�B�x� Z�l������������� ,P>`bt ������( L:\�d�� ��� /�$/6// Z/H/~/l/�/�/�/�/ .��/?�/2? ?V?D? f?�?n?�?�?�?�?�? 
O�?.O@O"OdORO�O vO�O�O�O�O�O�O_ _<_*_`_N_�_�_x_ �_�_�_�_�_oo8o o,ono\o�o�o�o�o �o�o�o�o "4 jX������ ����B�$�f�T� v������������؏ ��>�,�b�P�r����p�V 1�}� P8
�ܟ��B���TYPE\��HE�LL_CFG �.��͟  �	�����RSR ������ӯ������ �?�*�<�u�`�����ཿ������  �%�3�E�(�Q�\�ҰM�o¦p��d��2Ұd�]�K�:�HK 1�H� u������ �A�<�N�`߉߄ߖ� ������������&��8��=�OMM �H���9�FTOV�_EN�(�1�O�W_REG_UI���8�IMWAITr��a���OUT������TIM��;���VAL����_UNIT��K�1��MON_ALIA�S ?ew� ( he�#�������� ��Ҵ��);M�� q����d�� %�I[m �<������ !/3/E/W//{/�/�/ �/�/n/�/�/??/? �/S?e?w?�?�?F?�? �?�?�?�?O+O=OOO aOO�O�O�O�O�OxO �O__'_9_�O]_o_ �_�_>_�_�_�_�_�_ �_#o5oGoYokoo�o �o�o�o�o�o�o 1C�ogy��H ����	��-�?� Q�c�u� �������Ϗ Ꮜ���)�;��L� q�������R�˟ݟ� ����7�I�[�m�� *�����ǯٯ믖�� !�3�E��i�{����� ��\�տ�����ȿ A�S�e�wω�4ϭϿ� ���ώ����+�=�O� ��s߅ߗߩ߻�f��� ����'���K�]�o� ���>��������� �#�5�G�Y��}���������n��$SM�ON_DEFPR�O ������ �*SYSTEM*�  d=��RECALL ?}��� ( �}4c�opy frs:�orderfil�.dat vir�t:\tmpba�ck\=>ins�piron:12�732��s�� � }+.mdb:*.*CUZ��l�/x.:\��8R�o���0.a6H__�/ /�-?�b/t/�/ �/�F/�a/�/?? )�M�/p?�?�?� 8?J?��? OO%/7/ �/�/lO~O�O�/�/PO �/�O�O_!?3?�?W? h_z_�_�?�?B_�?�_ �_
oO/OAOSOdovo �oo�OHo�O�o�o +_�_O_�or�� �_:L_���'o 9o�o�on������o� �o[�����#5� Yj�|�����D�� �����1���U�f� x�������J�ӏ��� ���-���Q�b�t��� ����<�ϟa���� )�;�į߿pςϔϧ� ��˯]��� ��%��� ʿ[�l�~ߐߣ���F� ٿ�����!�3ϼ�W� h�z��ϱ�L����� ��
��/���S�d�v� �����>������� +�=�����r�� ��D��_�'� ����]�n����6�H����/#
x�yzrate 61 ���n/�/�/�%.'R4804� H/Z/�/�/?"3 .@�-a?s?�?�?* *�I?�$Y?�?�?O�!�$SNPX_�ASG 1�����9A�� P 0 '�%R[1]@1�.1O 	?�#% dO�OsO�O�O�O�O�O �O __D_'_9_z_]_ �_�_�_�_�_�_
o�_ o@o#odoGoYo�o}o �o�o�o�o�o�o* 4`C�gy�� �����	�J�-� T���c�������ڏ�� ���4��)�j�M� t�����ğ������ݟ �0��T�7�I���m� �������ǯٯ��� $�P�3�t�W�i����� ���ÿ����:�� D�p�Sϔ�wω��ϭ� �� ���$���Z�=� dߐ�sߴߗߩ����� �� ��D�'�9�z�]� ���������
��� �@�#�d�G�Y���}� ������������* 4`C�gy�� ����	J- T�c����� �/�4//)/j/M/ t/�/�/�/�/�/�/�/�?0?4,DPARAoM �9ECA_ �	��:P�4��0$HOFT_�KB_CFG  �p3?E�4PIN_�SIM  9K��6�?�?�?�0,@RV�QSTP_DSBº>�21On8J0SR� ��:� &� MULTIR�OBOTTASK�=Op3�6TOP�_ON_ERR � �F�8�APTN� �5�@�A�BRING_�PRM�O J0V�DT_GRP 1y�Y9�@  	�7 n8_(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 Dkhz���� ���
�1�.�@�R� d�v���������Џ�� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\������� ����ȯگ����"� I�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� tߛߘߪ߼������� ��(�:�a�^�p�� ���������� �'� $�6�H�Z�l�~��������������3VPRG_COUNT�6���A�5ENB��OM=�4J_U�PD 1��;8  
p2��� ��� )$6H ql~����� /�/ /I/D/V/h/ �/�/�/�/�/�/�/�/ !??.?@?i?d?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_�_�_Y?SDEBUG" � ��Pdk	�PSP_�PASS"B?~�[LOG ��+m�P�X�_�  �g�Q
M�C:\d�_b_M�PCm��o�o��Qa�o �vfSAV �m:dUb�U�\gSV�\TE�M_TIME 1]�� (�`��S���o	T1SV�GUNS} #'�k�spASK_OPTION" �g�ospBCCFGg ��| �f��v`����a&� �#�\�G���k����� ȏ������"��F� 1�j�U���y���ğ�� �ӟ���0��T�f��UR���S���ƯA� ����� ��D��nd� �t9�l���������ڿ ȿ�����"�X�F� |�jϠώ��ϲ����� ����B�0�f�T�v� xߊ��ߦؑ������ �(��L�:�\��p� ����������� � 6�$�F�H�Z���~��� ����������2  VDzh���� �����4Fd v������ //*/�N/</r/`/ �/�/�/�/�/�/�/? ?8?&?\?J?l?�?�? �?�?�?�?�?�?OO "OXOFO|O2�O�O�O �O�OfO_�O_B_0_ f_x_�_X_�_�_�_�_ �_�_oooPo>oto bo�o�o�o�o�o�o�o :(^Lnp �����O��$� 6�H��l�Z�|����� Ə؏ꏸ����2� � V�D�f�h�z�����ԟ ����
�,�R�@� v�d���������ίЯ ���<��T�f��� ����&�̿��ܿ�� &�8�J��n�\ϒπ� �Ϥ����������4� "�X�F�|�jߌ߲ߠ� ����������.�0� B�x�f��R������� �����,��<�b�P� ������x��������� &(:p^� ������  6$ZH~l�� ������/&/D/ V/h/��/z/�/�/�/��/�&0�$TBC�SG_GRP 2���%� � �1 
 ?�  /?A?+?e? O?�?s?�?�?�?�?�;�23�<d,� �$A?1	 H�C���6>���@E�5CL  B�p'2^OjH4J��B�\)LFY  A��jO�MB��?�IBl�O�O�@�JG_�@�  D	�15_ __$YC-P{_F_`_j\	��_�]@0�>�X�U o�_�_6oSoo0o~o�o�k�h�0	�V3.00'2	�m61c�c	*`�`�d2�o�e>�JC20(�a�i ,p�m�-  �0�����omvu1JCFG� ��% 1 �#0vz��rBrv�x����z � �%��I�4�m�X� ��|��������֏� ��3��W�B�g���x� ����՟������� �S�>�w�b�����'2 A ��ʯܯ������ E�0�i�T���x���ÿ տ翢����/��?� e�1�/���/�ϜϮ� �������,��P�>� `߆�tߪߘ��߼��� �����L�:�p�^� ������������  �6�H�>/`�r���� ������������  0Vhz8��� ���
.�R @vd����� ��//</*/L/r/ `/�/�/�/�/�/�/�/ �/?8?&?\?J?�?n? �?�?�?�?���?OO �?FO4OVOXOjO�O�O �O�O�O�O__�OB_ 0_f_T_v_�_�_�_z_ �_�_�_oo>o,obo Poroto�o�o�o�o�o �o(8^L� p������� $��H�6�l�~�(O�� ��f�d��؏���2�  �B�D�V�������n� ���ԟ
���.�@�R� d����v�������� Я���*��N�<�^� `�r�����̿���޿ ��$�J�8�n�\ϒ� �϶Ϥ�������ߊ� (�:�L���|�jߌ߲� �����������0�B� T��x�f������ �������,��P�>� t�b������������� ��:(JL^ ������ � 6$ZH~l� �^���dߚ // D/2/h/V/x/�/�/�/ �/�/�/�/?
?@?.? d?v?�?�?T?�?�?�? �?�?OO<O*O`ONO �OrO�O�O�O�O�O_ �O&__6_8_J_�_n_ �_�_�_�_�_�_�_"o oFo��po�o,oZo �o�o�o�o�o0 Tfx�H��� ����,�>��b� P���t���������Ώ ��(��L�:�p�^� ������ʟ���ܟ�  �"�$�6�l�Z���~� ����دꯔo��&� ЯV�D�z�h������� Կ¿��
��.��R��@�v�dϚτ�  ���� ��������$TBJOP_�GRP 2ǌ���  �?�������������x�JBЌ��9� �< �X�ƞ�� @���	� �C�� t�b�  C����>ǌ�͘Րդ�>���йѳ33=��CLj�fff?>��?�ffBG���Ќ�����t�ц�>;�(�\)�ߖ��E噙�;��h{CYj��  @h�~�B�  A�����f��C�  D�hъ�1��O��4�N����
:�/��Bl^��j�i��l�l����Aə�3A�"��D���Ǌ=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������<$�6�>B�\��T����Q�tsx�@g33@���C����y�1����>��Dh����������O<{�h�@i�  ��t��	� ��K&�j� n|���p�/��/:/k/�ԇ����!��	V3.0}0J�m61cIԃ*� IԿ��/�'� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�I�!CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;��;Q�UT,8�4` *���?�2���3\�X/�O��ESTPAR�S  ��	���H�R@ABLE 1%����0��
H�7Q 8��9
G
H
H�����
G	
H

H�
HYE��
H
H:
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_�^:BS _� �JGoYo ko}o�o�o�o�o�o�o �o1CUgy ����`#oRL�y�_ �_�_�_�O�O�O�O�O�X:B�rNUM  ����P���� V@P:B_CF�G ˭�Z�h�@���IMEBF_T�T%AU��2@�VE�RS�q��R {1���
 (�/����b� ����J� \���j�|���ǟ��ȟ ֟�����0�B�T�@��x�������2�_����@�
��MI_�CHAN�� � >��DBGLV����������ETHE�RAD ?��
O�������h������ROUT�!���!������SN�MASKD��U�255.���#������OOLOFS_�DI%@�u.�OR�QCTRL � ����}ϛ3rϧϹ��� ������%�7�I�[��:���h�z߯�APE?_DETAI"�G��PON_SVOF�F=���P_MON� �֍�2��S�TRTCHK ��^�����VTCOMPAT��O������FPROG �%^�%MULTIROBOTTݱx���9�PLAY&H���_INST_M�ް ������US8�q��LCK���QUICKME��=���SCREZ�}G�tps� @���u�z����_���@@n�.�SR_GR�P 1�^� �O����
��@+O=sa�� ��
m������ L/C1gU� y�����	/��-//Q/?/a/�/	1234567�0h�/�/@Xt�1����
 �}ipn�l/� gen.htm�? ?2?D?V?�`Panel� setupZ<}�P�?�?�?�?�?�? �??,O>OPObOtO �O�?�O!O�O�O�O_ _(_�O�O^_p_�_�_ �_�_/_]_S_ oo$o 6oHoZo�_~o�_�o�o �o�o�o�oso�o2D Vhz�1'� ��
��.��R�� v���������ЏG����UALRM��G ?9� �1�#� 5�f�Y���}������� џן���,��P���SEV  �����ECFG C��롽�A���   BȽ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �(� ��'�/SOFTPAR�T/GENLIN�K?curren�t=menupage,71,1��p��'�9� �3����edit�ҡ���0����D�� P���936��
��.�@� ��W�i�{��������� R�����/A�� ew����N� �+=O�s@�����C��f ��f//'/9/K/]/ `�/�/�/�/�/�/j/ �/?#?5?G?Y?�/�/ �?�?�?�?�?�?x?O O1OCOUOgO�?�O�O �O�O�O�OtO�O_-_ ?_Q_c_u__�_�_�_ �_�_�_��)o;oMo _oqo�o�_�o�o�o�o �o�o%7I[m � ����� ��3�E�W�i�{��� ���ÏՏ����� ��A�S�e�w�����*� ��џ�����oo O�a�s���������ͯ ߯���'���K�]� o���������F�ۿ� ���#�5�ĿY�k�}� �ϡϳ�B�������� �1�C���g�yߋߝ� ����P�����	��-� ?�*�<�u����� ��������)�;�M� ��������������� l�%7I[�� �����hz !3EWi�� �����v//�//A/S/e/P���$�UI_PANED�ATA 1������!  	�}w/�/�/0�/�/?? )?>? V�/i?{?�?�?�?�? *?�?�?OOOAO(O eOLO�O�O�O�O�O�Op�O�O_&Y� b�>RQ?V_h_z_�_�_ �__�_G?�_
oo.o @oRodo�_�ooo�o�o �o�o�o�o*<#�`G��}�-\ �v�#�_��!�3�E� W��{��_����ÏՏ ���`��/��S�:� w���p�����џ���� ��+��O�a��� ������ͯ߯�D�� ��9�K�]�o������� �ɿ���Կ�#�
� G�.�k�}�dϡψ��� �Ͼ���n���1�C�U� g�yߋ��ϯ���4��� ��	��-�?��c�J� ������������ ���;�M�4�q�X��� ��������% 7��[����� ��@��3 WiP�t��� ��/�//A/���� w/�/�/�/�/�/$/�/ h?+?=?O?a?s?�? �/�?�?�?�?�?O�? 'OOKO]ODO�OhO�O �O�O�ON/`/_#_5_ G_Y_k_�O�_�_?�_ �_�_�_oo�_Co*o goyo`o�o�o�o�o�o �o�o-Q8u�O�O}��������)�>��U-� j�|�������ď+�� Ϗ���B�)�f�M� �������������ݟ���XS�K�$UI�_PANELIN�K 1�U�  � � ��}1234?567890s��� ������ͯդ�Rq��� �!�3�E�W��{���@����ÿտm�m�&�4���Qo�  �0� B�T�f�x��v�&ϲ� ��������ߤ�0�B� T�f�xߊ�"ߘ����� �����߲�>�P�b� t���0�������� ����$�L�^�p��� ��,�>������� $�0,&�[�XI �m������ �>P3t�i ��Ϻ� -n�� '/9/K/]/o/�/t�/ �/�/�/�/�/?�/)? ;?M?_?q?�?�UQ �=�2"��?�?�?OO %O7O��OOaOsO�O�O �O�OJO�O�O__'_ 9_�O]_o_�_�_�_�_ F_�_�_�_o#o5oGo �_ko}o�o�o�o�oTo �o�o1C�og y�����B� 	��-��Q�c�F��� ��|�������֏� )��M���=�?��? /ȟڟ����"�? F�X�j�|�����/�į ֯�����0��?�? �?x���������ҿY ����,�>�P�b�� �ϘϪϼ�����o�� �(�:�L�^��ςߔ� �߸�������}��$� 6�H�Z�l��ߐ��� ������y�� �2�D� V�h�z����-����� ����
��.Rd G��}���� c���<��`r� �������// &/8/J/�n/�/�/�/ �/�/7�I�[�	�"?4? F?X?j?|?��?�?�? �?�?�?�?O0OBOTO fOxO�OO�O�O�O�O �O_�O,_>_P_b_t_ �__�_�_�_�_�_o o�_:oLo^opo�o�o #o�o�o�o�o �� 6H�l~a�� ������2�� V�h�K�������1 �U
��.�@�R�d� W/��������П��� ���*�<�N�`�r��/ �/?��̯ޯ��� &���J�\�n������� 3�ȿڿ����"ϱ� F�X�j�|ώϠϲ�A� ��������0߿�T� f�xߊߜ߮�=����� ����,�>���b�t� �����+��� ���:�L�/�p���e� ���������� ���6���ۏ��$�UI_QUICK�MEN  ����}��R�ESTORE 1�٩�  �
�8m3\n��� G����/�4/ F/X/j/|/'�/�/�/ /�/�/??0?�/T? f?x?�?�?�?Q?�?�? �?OO�/'O9OKO�? �O�O�O�O�OqO�O_ _(_:_�O^_p_�_�_ �_QO[_�_�_I_�_$o 6oHoZoloo�o�o�o �o�o{o�o 2D �_Qcu�o��� ����.�@�R�d� v��������Џ⏜oSCRE� ?�u1sc� Wu2�3�4�U5�6�7�8��USER�����T���ks'���4���5��6��7��8���� NDO_CFoG ڱ  � � � PDATE� h��N�one�SEUFRAME  �ϖ��RTOL_�ABRT����E�NB(��GRP �1��	�Cz  A�~�|�%|�������į֦��X�� UH�X�7�MSKG  K�S�7�N�%uT�%������VISCAND_wMAXI�I�3����FAIL_IM)GI�z �% #S����IMREGNUMrI�
���SIZI��� �ϔ,�O�NTMOU'�K��Ε�&����a���a��s��FR:\�� �� MC:\�(�\LOGh�B@Ԕ !{��Ϡ������z M�CV����UD1& �EX	�z ���PO64_�Q�n�n6��PO!�CLI�Oڞ�e�V��N�f@`�I�� �=	_�SZVmޘ;��`�WAImߠ�STAT �k�B% @��4�F�T�$#��x �2DWP  ��P G���=��͎�������_JMPERRw 1ޱ
  �p�2345678901���	�:�-� ?�]�c������������������$�MLO�W�ޘ�����_TI�/�˘'��MPH?ASE  k�ԓ�� ��SHIFT�%�1 Ǚ��< z��_��� �F/|Se� ������0// /?/x/O/a/�/�/�/��/�/����k�	�VSFT1[�	uV��M+3 �5��Ք p����A� W B8[0[0�Πpg3a1Y2�_3Y�7#ME��K�͗	6eѮ��&%��M��ഠb��	��$��T?DINEND3�4���4OH�+�G1�OSp2OIV I���]LRELEvI��4.��@��1_ACTIV�IT��B��A �`m��/_��BRDB���OZ�YBOX ��ǝf_[��b�2��TI190�.0.�P83p\��V254p^�Ԓ	 �S�_�[b���robo�t84q_   �p�9o[�pc�PZoMh�]Hm�_Jkx@1�o�ZABCd��k�,���P[�Xo} �o0);M�q ��������$>��aZ�b��_V