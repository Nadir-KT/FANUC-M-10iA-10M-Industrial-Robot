��   %��A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING���< �PLC�L* ��ST�A� mTRQ_M<��LINK"2&�SX<*Y<*Z/)I�I*IW*Ie$ �R�V* $� E�NBpV_DEBuU��!PNU;%�� UNEVEox�  �$�AS�S  �����!����� VIRTUAL�/�!'� 1 5_� ��� ��R?=?v?a?�?�? �?�?�?�?�:HE� M�!8O&O ���߿����]B�   ^��MO�O�? KL�O�O�O�O�O�OzK1_7R _]_o_Z_�_���d�_�_�_�_��=gL���_o?�o��@�3oXojo|o�o �o�o5�o�o�o�o #�$�R)SAw62k������ �#�5�G��"� M�s� ��������͏ߏ����'�9��#�$% �1521D}U%a{����_��}_ ԟ��������R� =�v�a�������ͯ�� ������<�'�`�K� ]���������޿ſϯ �ӿ8�Ͽ\�Gπ�k� �Ϗϡ���������"� 	��U��|�ߠߋ� �߯��������	�B� -�f�M�Wߙ�[���W� �������,��)�b� M���q����������� ��(L7p[ m�������� !�H�lW�{ �����/�2/ /#e/'/�/#/�/�/ �/�/�/�/�/.??R?x=?v?;g�$RV[��b�8k?�?c?  BFo;gx�?O(O�:OLO^OpO�O�O  �h 
�  :�  B`����������S�������������@$���\��[���C���@�@6r���C��O_ _,_>_P_b_t_�_�_ �_�_�_�?�_�_o(o OLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��o=o2��V�1o z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�C�`�G�Y���q� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|σ��χ��ϟ��� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t��� ������������(� :�L�^�p��������� ������ $6H Zl~����� ����2�Bh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? <?N?5?r?M�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ jQ