��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1��GPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|�(�ARG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� � $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WA��471�8GW+0�$�Y $DB� 6CkOMW!2MO� �H.	 \rVE�1$F�RA{�$O�UDcB]CT_MP1_FtE2}G�1_�3�B�2?GX�D�#
 d �$CARD_E�XIST4$FSSB_TYP~!AHKBD_SNB֒1AGN Gn �$SLOT_N�UM�APREV4DEBU� g1G �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��U0LETE_O�K�BUS�P_CR�A$;4AV� 0/LACIw1�Rp�@k �1$@MEN�@$D�V�Q`Pv�VA{QL� OU&R ,A�0�!z� B� LM_O�z
eR�"CAM_;�1 xr$�ATTR4�@� A�NNN@5IMG_�HEIGH�AXcWoIDTH4VT� ��UU0F_ASP�EC�A$M�0E�XP�.@AX�f��CF�D X '$GR� � S�!.@=B�PNFLI�`�d� UIRE 3T!GOITCH+C�`N� MS�d_LZ`AC�"��`EDp�dL� J�4S�0� <za�!p�;G0 � 
?$WARNM�0f�!�@� -s�pNST�� CORN�"a1F�LTR{uTRAT�� T}p  $ACCa1�p��|{��rORI�P�C�kR�T0_S~B\qHG�,I1 [ Th�`�"3I�pTYD(�@*2 3`#@� X�!�B*HDDcJ* TCd�2_�3_�4_�U5_�6_�7_�8_��94? �CO�$ <� �o�o�hK3 1�#`O_Mc@AC �t � E#6NGPvABA� �c1�@Q8��`,��@nr1�� d�P�0e�]p� cvnpUP&Pb2�6���p�"J�p_R�rPBC��J�rĘߜJV�@U� B��s}�g�1�"YtP_*0OF�S&R @� RO1_K8T��aIT�3T�ONOM_�0�1p�p3� >��D �� �Ќ@��hPV��mEX�p� �0g0ۤ�p�r�
$TF�2C$M�D3i�TO�3�0U�� F� ��H�w2tC1(�Ez�g0�#E{"F�"F�40C�P@�a2 �@$��PPU�3N1)ύRևAX�!D�U��AI�3BU�F�F=�@1 |Xpp���pPIT� +PP�M�M�y���F�SIMQS@I�"ܢVAڤT�&=�Nw T�`(zM�x�P�B�qFACTb�@EW�P1�B�Tv?�MC� �$*1JB`p�*1�DEC��F���S.yS��� �H0�CHNS_EMP�1�$G��8��@_�4�3�p|@P��3�TCc�(r/�0-sx���ܐ� MBi��!����J�R� i�SEGFRR��Iv �aR�Tp�N�C��PVF4|?�bx &� �f{uJc!�Ja��� !2�8�ץ�AJ���SIZ�3S�c�B�TM���g�|��JaRSINFȑ b���q�۽�н�����L�3�B���CRC�e�3CCp��� �c��mcҞb�1J�c�P��.����D$ICb�Cq�5r�ե��@v�'����EV���zF��_J��F,pN��ܫ��?�4�0A�! � r���h�Ϩ��p�2@�͕a�� �د\q}R�Dx Ϗ ��o"27�!ARV�O`�C�$LG�pV�B@�1�P��@�t�aA�0�'�|�+0Ro�� M�Ep`"1 CRA 3 AZV�g6p��O �FCCb�`�`F��`K������ADI ��a�A�bA'�.p ��p�`�c�`S4PƑL�a�AMP��-`Y�3�P�M�]pUR��QU�A1  $@TITO1/S@S�!����"0�DBPXWO��zB0!5�$SK��L�2�DBq�!"�"v�PR�� 
� 8=����!# @q1�$2�$z�O�L�)$�/���� )%�/�$C�!&?�$gENE�q.'*?�PA
�!RE�p2(�H ��O�07#$L|3$$�#�B�[�;���FO_D��ROSr�#�������3RIGGE�R�6PApS����E�TURN�2�cMR-_8�TUw��0�EWM��M�GN�P���BLAH�<E��y�P��&$P�" �'P@�Q3�CkD{��DQ���4�11��FGO_AWAY�B�MO�ѱQ#!��DCS_�)  �PIS� I gb @{s�C��A��[ �B�$�S��AbP�@�EW�-�TNTVճ�BV �Q[C�(c`�UWr�P��J��P�$0��SAF�E���V_SV�bEOXCLU��n'ONL2��SY�*a�&�OT�a'�HI_�V�4��B���_ #*P0� 9�_z��po "�TSG�� +nrr�@6Acc *b��G�#@E�V.iHb>?fANNUN$0.$�fdID�U�2�S C@�`�i�a��j�f�"��pOGI$2,O�c$FibW$}�OT9@��1 $DUM�MYk��da��dn��� � �E- ` ͑HE4(sg�*b�S|AB��SUFFIW�[�@CA=�c�5�g6�a�"MSW��E. 8Q�KEYI5���TM�10s�qA�vIN��#�b��/ D��HOST_P!�rk��ta�`�tn��tsp�pEMӰ�V��� SBLc U}LI�0  8	�=ȳ#��!Tk0�!1� � $S��ESAMPL��j�۰f爒�f���I�0��[ $SUB�k�#0�Cp��T�r#a�SAVʅ ��c���C��P�f�P$n0E�w YN�_B#2 0Q�D�I{dlpO(��9#�$�R_I�� �ENC2_S� 3  5�C߰�f�- �SpU����!!4�"g�޲�1T���5X�j`ȷg��0��0K�4�AaŔAV�ER�qĕ9g�DSP�v��PC��r"�(���ƓVALU�ߗHE�ԕM+�I�Pճ��OPP ���TH��֤��P�SH� �۰F��df��J� ��q�C1+6� H�bLL_DU s�~a3@{��3:����OTX"���s�ʡR_NOAUT5O�!7�p$)�$�*��c4�(�Cy��8�C, �"ɢ'�L��� 8H *8�LH <6����c"� �`, `Ĭ�kª�q��@q��sq��~q��7���8��9��0����1���1̺1ٺ1�1��1 �1�1�2R(�2����2̺2ٺU2�2�2 �2�U2�3(�3��3���̺3ٺ3�3�3* �3�3�4(�a8��?��!9 <�9�&�z��I��1���M���QFE@'@� : y,6��Q? �@FP?9��5�9�E�@A��A� ;�p$TP�$�VARI:�Z���U�P2�P< ���TDe���K`Q����"���BAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�HH  ��P�ȢF@|`�!>t ;E�4�sC�ST�D� D���c�<� 	 C��{��_���l����R  ���FORC�EUP?b��FLUS�`H�N>�F ��^�RD_CM�@E������� ��@vMP��REMr F�Q��1��P���7Q
K4	NJ��5EFFۓ:�@I�N2Q��OVO�O{VA�	TROV���DTՀ�DTMX� ��@�
ے_P`H"p��CL��A_TpE�@�pK	_(�FY_T��v(��@%A;QD� �����`�!0tܑ0RQ��"�_�a����M�7�sCL�dρRIV'��{��EARۑIOFHPC�@����B�Bƅ�CM9@���R ��GCLF�e!DaYk(M�ap#5Tu�DG��� �%aFsSSD �s? P�a(�!�1���P_�!�(J�!1��E�3�!3�+=5�&�GRA��7��@��;�PW��OyNn��EBUG_S�D2H�P{�_E �A �p�Q _�TERM`5Bi5�K@�ORI#e0C�i5���SM_h�P��e0D�9TA�9�E�9UP\�F�3 -�A{�AdPw3>S@B$SEG�:� �EL{UUSE�@NFIJ�B$�;1�<�4�4C$UFlP=��$,�|QR@���_G90Tk�D�~SN;ST�PAT�����APTHJ3Q�E �p%B`�'EC����AR$P�I�aSH�FTy�A�A�H_SGHORР꣦6 �0�$�7PE��E�OV�R=��aPI�@�Uz�b �QAYLOW���IE"�r�A��?���ERV��XQ�Y ��mG>@�BN��U����R2!P.uASY1MH�.uAWJ0G�т�Eq�A�Y�R�U�d>@��EC���EP�;�uP;�6WOR>@Mv`�0SMT6��G3�GR��13�aP�AL@���`�q�uH ׸ ���TO�CA�`P	P�`$OP����p�ѡ�`e0O��RE�`�R4C�AO�p낎Be�`R�Eu�h�A���e$PWR�IM�u�RR_�c C�K�b=B I&2H|���p_ADDR��?H_LENG�B�q��q�q$�R��S�J6ڢSS��SKN��u`���u̳�uٳSE�~A�(�HS��[MN�!K���0��b����OLX���p����`ACRO 3pJ�@��X�+��Q���6�OUP3�b_"�IX��a�a1��}� ������(��H��D���ٰ��氋�IO
2S�D������`<�7�L $l��`�Y!_OFFr�P�RM_��ɡHT�TP_+�H:�M (|pOBJ]"�p��[$��LE~Cd�>��N � ��֑�AB_�TqᶔSؙ`H�LVh�KR�"uHITCOU���BG�LO�q ���h�����`��`sSS� ���HW��#A:�Oڠ<`IN�CPU2VISIOW�͑��n��to��t�o�ٲ�IOLN.��P 8��R��p�$SLob P7UT_n�$p���P& ¢ ��Y F_�AS�"Q��$L ������Q  U�0	P�q��^���ZPHY���-��y��UOI �#R `�K���@�$�u�"pP�pk���$�����Y�UeJ5�S-���NE6W�JOGKG̲DISĖ���Kp���#T �(�uAVF�+`�CTyR�C
�FLAG2v��LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w� m� _�{0a�^��cg���4� ����Ǝ���{0��� �SCH_���a�SLN�d�VW���AE�"����4��UM��Aљ`LJ�@�DAUf�EAU�p��d|�r��GH�bY���BOO>��WL ?�6 �IT��y0�REC��SCR ܓ��D
�\���MARG m�!��զ ��d%�����S����W���U�� �JGM[�MNC�HJ���FNKEY�\�K��PRG��UqF��7P��FWD��HL��STP��V`��=@��А�RS��HO`����C9T��b ��7�[�UL���6� (RD� ����Gt��@CPO��������MD��FOCU��RGE]X��TUI��I��4�@�L��� ��P����`��P��9NE��CANA��B�j�VAILI�CL� !�UDCS_HII4��s�O�(!�S���S��D�^��BUFF�!X�5?PTH$m����v`�ěԃ�AtrY��?P��j�3��`O+S1Z2Z3Z�|�� Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�C���K�&&8���![ LQ��+00� 	P���`#qdt
�U�dt�9��_ \ ��`4Г�\��Ѩ#\0C�4�] ��CLD�PL��UTRQLI��dڰ�)�$FLG &�� 1�#�D���'�B�LD�%�$�%ORGڰ5�2�PVŇVY8��s�T�r�$}d^ ����$6��$�%S�`T�� �B0�4�6RCLMC�4]?o?�9�渰MI�p}d_ d�=њRQ��DgSTB�p� ;Fl�HHAX�R JH>dLEXCESr��RBM!p�a`� /B��TE��`a�p=F_A7Ji��KbOtH:� K�db \Q��n�v$MBC�LI|�~)SREQUIR�R��a.\o�AXDEBUTZ�ALt M��c�b��{P����2ANDRѧ`�`d;�2��f�SDC��N�INl� K�x`��X� N&��atZ���UPST�w ezrLOC��RIrp�EX<fA�p�9AAODAQn��f XY�OND�rMF,Łf�s"���}%�e/� ��AFX�3@IGG�� g ��t"��ܓs#N�s$R�a%��iL���hL�v�@�DAT	A#?pE�%�tR���Y�Nh t W$MD`qI}�)nv� ytq�ytHP`�Pxux��(�zsANSW)�Pyt@��yuD+�)\b����0o�i �@C�Uw�V�p 0XeRR2��j Du�{Q��~7Bd$CALIA@���G��2��RI�N��"�<E�NTE��Ck�r^�آXb]���_N�qlk���9��D���Bm��DIVFFDH�@���qnI�$V,��S�$��$Z�X�o��*����oH ?�$BELT�u!_ACCEL�.�~�=�IRC�� ����D�T�8�$PS�@�"L  Šp��#�^�S�Eы T�PAT!H3���I���3x�p�A_W��ڐ���2n�C��4�_MG��$DD��T���$FW�Rp9��I�4���DE7�PPAB�N��ROTSPE!E�[g�� J��[��C@4�x�$US�E_+�VPi��S�YY���1 qYNr!@A�ǦOFF�qnǡMOU��NG����OL����INC �tMa6��HB��0HBENCS+�8q9Bp�X4�FDm�IN�Ix�0]��B��VE��#�>y�23_UP񕋳/LOWL���p� B���Du�9B#P`��x ���BCv�r�MO3SI��BMOU��@��7PERCH  ȳOV��â
ǝ� ���D�ScF�@MP����� Vݡ�@y�j��LUk��Gj�p�UPp=ó���ĶTRK�>�AYLOA�Qe� �A��x�����N`�F��RTI�A$��MO UІ�HB�BS0�p7D5����ë�Z�DU�M2ԓS_BCKLSH_Cx�k�� ��ϣ���=���ޡ< �	ACLAL"q�p�1м@��CHK� :�S�RTY���^�%E1Qq_�޴_�UM�@�C#��S�CL0�r�LMT_OJ1_L��9@H��qU�EO�p�b�_�e�k�e�SPC��u�L��N�PC�N�Hz �\P��C�0~"XT\��CN_:�N9�L�I�SF!�?�V����U�/���x�T���CB!�SH�:��E� E1T�T����y���T�f�PA ��_P��_� =������!����J6 L�@���OG�G�TORQU��ONֹ��E�R0��H�E�g_W2��ā_郅���I*�I�I��Ff`xaJ�1�~1�VC3�0BD:B�1�@SBJRKF9~�0DBL_SM�:�2M�P_DL2GRV�����fH_��d���CcOS���LNH ��������!*,�aZ���fcMY�_(�TH���)THET0��N�K23���"��C-B�&CB�CAA�B��"��!��!�&SB8� 2�%GTS�Ar�CIMa�����,4#<97#$DU���H�\1� �:Bk62�:AQ�(rSf$NE�D�`I ��B+5��$̀�!�A�%�5�7���LCPH�E�2���2S C%C%�2-&FC0JM&̀V�8V�8߀LUVJV!KV/KV=KUVKKVYKVgIH�8@FRM��#X!KH/KUH=KHKKHYKHgI�O�<O�8O�YNO�JO!KO/KO=KO*KKOYKOM&F�2�!�+i%0d�7SPBA?LANCE_o![c�LE0H_�%SP�c� &�b&�b&PFULC�h�b�g�b%�p�1k%�UTO_<��T1T2�i/�2N��"�{�t#�Ѡ�`�0�*�.�T��O�À<�v INSEG"�ͱREV4vͰl�gDIF�ŕ�1lzw6��1m�0OBpq�ь�?�MI{���nL�CHWARY�_�A�B��!�$MEC�H�!o ��q�AX���P����7Ђ�`n� 
�d(�U�RO�B��CRx�H���(�MSK_f`��p P �`_���R/�k�z�����1 S�~�|�z�{���z��q�INUq�MTC�OM_C� �q � ���pO�$ONOREn����p�Ђr 8p GRle�uSD�0AB��$XYZ_DAx�1a���DEBUUqX������s z`$��wCOD�� L����p�$BU�FINDX|� � <�MORm�t $فUA��֐�Р�\�<��rG��u� � $SIMUL  S�*�Y�̑a��OBJE�`̖AD�JUS�ݐAY_	IS�D�3���_FI�=��T u 7�~�6�'��p} =��C�}p�@b�D��FRiIr��T��RO@ �\�E}��y�OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1�0e��M��ED}�*�p ��N�PMֲ�����x�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B��2�G�B�_�M��y�q�E� x �Hw��p��ATUS
W���C�0o�s��çBTM�ǌ�I��k�4��x�԰q�y �Dw�E&���@E��r��7��жЗ�EXE��ἱ�����f �q�z @w���UP�'��$�pQ�XN����������� ��PG΅{ h �$SUB����0_����!�MPWAI2v�P7ã�LOR����F\p˕$RCV?FAIL_C����BWD΁�v�DE�FSP!p | Lw���Я�\���UNI+�����H�RX�+�}_L\pP��x�t���p�}H�> *�j�(�s`~�N�`KSETB�%�J�PE �Ѓ~��J0SIZAE\���X�'���S��OR��FORMA�T�`��c ��WrEeM�t��%�UX���G��PLI��p��  $ˀP_�SWI�pq�J_P�L��AL_ ������A��B��� C���D�$E���.�C_�U�� ?� � ����*�J3K0����TI�A4��5��6��MOM��������ˀB��AD������l����PU� NR������u��m��� A$PI�6 q��	�����K4��)6�U��w`��S/PEEDgPG�� ������Ի�4T��� � @��SA�Mr`��\�]��MOV_�_$�npt5�H�5���1���2��@������'�S�Hp�IN�'�@�+�����4($4+T+G�AMMWf�1'�$GGET`�p���Da�z��

pLIBR>ѺII2�$HI=�_�g�t��2�&E;��(A�.� �&LW�-6<��)56�&]��v�p��V���$PDCK���q��_?�����q�&���7��4����9+� �$_IM_SR�pD�s0�rF��r�rLE���!Om0H]��0����ܬpq��PJqUR_SCRN�FA����S_SAVE_DX��dE@�NOa�CA A�b�d@�$q�Z�Iǡ s	�I� �J�K� ��� �H�L��>�"hq� �����ɢ�� @bW^US�A�,M4���a��)q`��3�W@W�I@v�_�q���MUA�o�� � $P9Y+�$W�P�vNG�{��P:��RA�0�RH��RO�PL������q� ��s'�X;�O�I�&�Zxe ���m��# p��ˀ�3s�O@�O�O�O�O�aa�_т� |��q�d@��.v ��.v��d@��[wFv��9E���% 
��rJ;B�w�|�tP���PMA�QUa ���Q8��1�Q�TH�HOLW�Q7HYS��ES��q�UE�pZB��Oτ�  ـPܐ(�A��(��v�!�t�O`�q���u�"���FA��IR#OG�����Q2����o�"��p��INF�Oҁ�׃V����R�vH�OI��� (�0SLEQ������BY�����Á��P�0Ow0���!E�0NU��AUT<�A�COPY�=�(/�'��@Mg�N��=��}1������ ��RG4��Á���X_�P�C$;ख�`��W���P��@�������E�XT_CYC b�HᝡRpÁ�r��_NAe!А����ROv`	�� �s ���POR_�1�E2�SRV �)l_�I�DI��T_� k�}�'���dЇ�����U5��6��7��8i��H�SdB���2�$R��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,�0FL`�o@SYN��K�M��Ck��PWR+�9ᘐ���DELA}�dY֟pAD�a�qQSwKIP4� �A�Z$�OB`NT����P_$�M�ƷF@\b Ipݷ�ݷ�ݷd�� ��빸��Š�Ҡ��ߠ�9��J2R�� ��� 4V�EX� TQQ����TQ������� ��`�#�RD�C�V� �`��X)�R�p�����r��~m$RGEAR_� sIOBT�2FLG��LfipER�DTC����Ԍ���2TH2N<S}� 1���uG T\0 ����u�M\Ѫ`I�d	ּ�EF�1Á� yl�h��ENAB��cTPE�04�]�� ��Y�]��ъQn#��*���"���ҏP��2�Қ �߼�����������3�қ'�9�K�]�o����4�Ҝ����������� I��5�ҝ!�3�E�W�i�{�
��6�Ҟ��������(������7�ҟ-�?Qcu��8�Ҡ��������SWMSKÁ�l��a��EkA�rREMO[TE6�����@0�݂TQ�IO}5�QISTP�QR�W@��� �pJ�����p����E�"$DSB_SIGN�1�UQ�x�C\��S2�32���R�iDE?VICEUS�XR>SRPARIT��4!_OPBIT�QI�OWCONTR+��TQ��?SRCU� M~pSUXTASK�3�N�p�0p$TATU��P �H �0������p_XPC)�$�FREEFROMqS	pna�GET�0.��UPD�A�21��RSP� :���� !$USA�N�na&����ERI��0�RpRYq5*"_�j@�Pm1�!�6WR	K9KD���6��Q?FRIEND�Q�R�UFg�҃�0TOO�L�6MY�t$L�ENGTH_VT\�FIR�pC�@ˀyE> +IUFIN-R:M��RGI�1ÐOAITI�$GXñl3IvFG2v7G1�0��p3�B�GPR�p�1�F�O_n 0��!R�E��p�53҅U�TCp��3A�A�F�G(��":���e1n!���J�8�%���%]� ��%�� 74�X �O0�L��T�3H@&��8���%b453GE�IW�0�WsR�TD�� ��T��M����Q�T]�{$V 2���H�1�а91�8�02�;2k3�;3�:ifa �9-i�aQ��NS��ZRS$V��2BVwEV��2A Q�B;���� �&�S�`��F�"�k�@��2a�PS�E ��$r1C��_$Aܠ6wPR��7vMU�cqS�t '�|(�529�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx_�����BSOC����N��DUMMY�14�p@SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW_C��U��S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}����_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�S�A�pC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EG� �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G + AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC  o�ER|f�5� � $�@�_ A��!�PO���à�0#�
�_M�RAt�� d r� T��ٔERR��L��;TY&���I��qV�0�cz�TOQ�d�PL[ �d�"�� ?�|w�! � pp`qT)0���_V1VrP�aӔ����2ٛ2薈E����@�H�E����$W�����V!��$�P��o�cI���aΣ	 HELL�_CFG!�� 5��B_BAS�q�SR3��� Ea#Sb���1�U%��2��3��4��U5��6��7��8����RO����I0�0NL�\CAB+�����ACK4�����,�\@p2@�&�?�_PUﳳCO. U�OUG�P�~ ����m�������T=Pհ_KAR�l�&_�RE*��P���|�QUE���uP�����CSTOPI_AL7�l�k0��h��]�l0SEM�4�(��M4�6�TYN�SO���DIZ�~�A������m_TM�MA'NRQ��k0E�����$KEYSWI�TCH�ӵ�m���H=E��BEAT��|�E- LE~�����U±�F!Ĳ���B�O_�HOM=OGREFUPPR&��y!� �[�C��O��-EC�OC��Ԯ0_IOC1MWD
�a�	�m��� � Dh1���	UX���M�βgPgC�FORC��� ���OM.  �� @�5(�U�#P�, 1��, 3��4�5	�NPX_A�St�� 0��AD�D���$SIZ>��$VAR����TIP/�.��A�ҹM�ǐ��/�1�+ �U"S�U!Cz���F'RIF��J�S���5Ԓ�NF�� �� �� xp`SI��TqE�C���CSGL��	TQ2�@&����� ���STMT��,�P� �&BWuP��SHsOW4���SV��$�� �Q�A00�@Ma}���� ������&���5��6���7��8��9��A ��O ���Ѕ�Ӂ���0��F��� G��0G ���0G���@G��PTG��1	1	1	U1+	18	1E	2��U2��2��2��2��U2��2��2��2��U2��2	2	2	U2+	28	2E	3��U3��3��3��3��U3��3��3��3��U3��3	3	3	U3+	38	3E	4�U4��4��4��4��U4��4��4��4��U4��4	4	4	U4+	48	4E	5�U5��5��5��5��U5��5��5��5��U5��5	5	5	U5+	58	5E	6�U6��6��6��6��U6��6��6��6��U6��6	6	6	U6+	68	6E	7�U7��7��7��7��U7��7��7��7��U7��7	7	7	�7+	78	7E��V�P��UPDs� � �`NЦ�5�Y�SLOt�� � �L��d���A�aT�A�0d��|�ALU�:ed�~�CUѰjgF�!aID_L�ÑeH�I�jI��$FILcE_���d��$2��SeSA>�� h�O��`E_BLCK���b$��hD_CPUyM�yA��c�o�dxb����R �Đg
PW��!� oqLA��S=�ts�q~tRUN�qst�q~t����qst�q~t ��T��ACCs���X -$�qLE�N;��tH��ph�_�I���ǀLOW_AXMI�F1�q�d2*�AMZ���ă��W�Im�8ւ�aR�TOR��p�g�D�Y���LAC�Ek�ւ�pV�ւ~�_�MA2�v�������T#CV��؁��T��ي �����t�V����V�IJj�R�MA���J���m�u�b����q2�j�#�U�{�t�K�JK���VK;���H���3f��J0����JJ��;JJ��AAL��ڐ(��ڐԖ4Օ5����N1���ʋƀW�LrP�_(�g�k(�q�r�� `�`GR�OUw`��B��N�FLIC��f�RE�QUIRE3�EB�U��qB���w�2�����p���q5�p��{ \��APPR��iC}�Y�
ްEN٨�CLO7��S_M���H���u�
�qu�7� ���MC������9�_MG��C�C�o��`M�в�N�BRKL�NOL|�N�[�R��_LINђ�|�=�J����Pܔ������������������6ɵ�̲8k�+��q���� ��
��q�)��7�PATH 3�L�B�L��H�wࡠm�J�CN�CA��ؒ�ڢB�IN�rUChV�4a��C!�UM��!Y,���aE�p�����ʴ���PAYL�OA��J2L`R'_AN�q�Lpp����$�M�R_F2�LSHR��N�LO�ԡ�Rׯ�`ׯ�ACRL_G�ŒЛ� �r�Hj`߂$HM�^��FLEXܣ�q}J�u� :� ������������1�F1�V�j�@�@R�d�v�������E�� ��ȏڏ����"�4� q���6�M���~��U��g�y�ယT��o�X ��H������藕?� ����ǟِݕ�ԕ�����%�7��JJ�� � V�h�z����`AT�採@�EL��� S��J|��v��JEy�CTR���~�TN��FQ��H�AND_VB-����v`�� $��Fa2M����ebSW?���'��� $$	MF�:�Rg�(x�,4�%��0&A�`�=���aM)F�AW�Z`i�A�w�A��X X�'pi�D*w�D��Pf�G�p�)CSTk��!x��!N��DY�pנM�9$`%� ��H��H�c�׎���0� ��Pѵڵ������������� ���1��R�6��QOASYMvř����v��J���cі�_SH>��ǺĤ�ED����������J�İ%�p�C�IDِ�_VI��!X�2PV_UN!IX�FThP�J��_R �5_Rc�cTz�pT�V�݀@���İ�߷��U $�������Hqpˢ3��aEN�3�SDI����O4d��`J�� x g"IJAAȱz�aabp�coc��`a�pdq�a� �^�OMME��� h�b�RqAT(`PT�@ � S��a7�;�Ƞ�@ȷh�a�iT�@<� �$DUMMY9�Q�$PS_��R�FC�  S�v ��p���Pa� XXƠ���STE����SBRY�M21_�VF�8$SV_E�RF�O��LsdsCLRJtA��Odb`�O�p � D ?$GLOBj�_LO���u�q�cAp�rܛ@aSYS�qADqR``�`TCH  � ,��ɩb�oW_NA����7��SR���l ���
*?�& Q�0"?�;'?�I)?�Y) ��X���h���x����� �)��Ռ�Ӷ�;��Í�v�?��O�O�O�D�XOSCRE栘p�����ST��s}�y`���p�/_:HA�q� TơgpTYP�b���G�aG���Od0I�S_䓀d�p�UEMd� ����ppyS�qaRSM_�q�*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCO�U��S�Ԕ 1�!�UE&��Ubwr���PROGM�FL�@$CUgpPO��Q���UI_�`H>� � 8�� �_HE�PS�#��`?RY ?�qp�b���dp�OUS>�� � @6p�v�$BUTTp�R|pR�COLUMq�<e��SERV5��PANEH�q� w� �@GEU��Fy��)$HE�LPõ)BETERv�)ෆ���A  � ��0��0��0�ҰIN簪c�@N(��IH�1��_�o ֪�LN�r'� �qpձ_ò=��$H��TEX8l����FLA@��/RELV��D`���������M��?,@�ű�m����"�USRVIEW�q�� <6p�`U�`��NFI@;�FOsCU��;�PRI@�m�`�QY�TRI}P�qm�UN<`�Md� #@p�*eW�ARN)e�SRT+OL%��g��ᴰ�ONCORN��RA�U����T���w�V�IN�Le� =$גPATH9�ג�CACH��LOG�!�LIMKR���x�v���HOST��!�b�R��OgBOT�d�IM>�	 �� ���Zq��Zq;�VCPU_�AVAIL�!�EX	�!AN���q�`�1r��1r��1��\��p�  #`C�����@$TOOLz�$��_JMP�� ���e$S�S����VSHI9F��Nc�P�`ג��E�ȐR����OS�UR��Wk`RADILѮ��_�a��:�`9a��`a�r��LULQ�$OUTPUTg_BM����IM��AB �@�rTILNSCO��C7� ������&�� 3��A���q���4m�I�2G�W(��prLe�}��yDJU��~N�WAIT֖��}��{�%! NE޿u�YBO�� ?�� $`�tv�SB@TPE��NECp�J^FY�.nB_T��R�І �a$�[YĭcB��dM�,�F� �p�$�pb�OP?�MAS��_DO�!QT�pD��ˑ#%��p!"DELAY�:`7"JOY�@(�nCE$���3@ �xm��d�pY_[�!"�`�"��[����P? S� Z�ABC%��  �$�"R��
E`��$$CLAS������!pn�� � VIRT]��/ 0gABS����1 5�� < `D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX8i}0-�AXL�p���"�63  �{tIqN��qztPRE�����v�p�uLAR�MRECOV �9�rwtNG�� �.;	 =#��
�.�0PPLIMC��?5�p��Handl�ingTool �o� 
V7.5�0P/23 �!��PB��
��_�SWt� UP�!� x�F0��t����An�v� 8[64�� �it��y� N2 �7DA5�� �j� QBy@��o�Noneis�ͅ˰ ��T��]�!LAA[xyrP_l�V�utT��s9�UTO�"�Њt�y��HGAPCON
0g�1��Uh�oD 1581����̟ޟry����/Q 1���p �,�蘦���;�@���q_��"�" g�c�.�H����D�HTTHKYX��"�-�?�Q��� ɯۯ5����#�A�G� Y�k�}�������ſ׿ 1�����=�C�U�g� yϋϝϯ�����-��� 	��9�?�Q�c�u߇� �߽߫���)����� 5�;�M�_�q���� ����%�����1�7� I�[�m���������� !����-3EW i{����� �)/ASew ����/��/ %/+/=/O/a/s/�/�/ �/�/?�/�/?!?'? 9?K?]?o?�?�?�?�? O�?�?�?O#O]����TO�E�W�DO_CLEAN��7��C�NM  � �__/_A_S_�DSPDRYR�O&��HIc��M@�O�_ �_�_�_oo+o=oOo aoso�o�o���pB��v# �u���aX�t�������9�PLUGGp���G��U�PRCvPB�@��_�or�Or_7�SEGF}�K[mwxq�O�O������?rqLAP�_�~q�[�m���� ����Ǐُ����!�|3�x�TOTAL�f| yx�USENU�p��� �H���B��R�G_STRING� 1u�
�kMn�S5�
ȑ�_ITEM1Җ  n5�� ��$�6� H�Z�l�~�������Ư�د���� �2�D��I/O SIG�NAL̕Tr�yout Mod�eӕInp��S�imulated�בOut���OVERR�P =� 100֒In� cycl��ב�Prog Abo�r��ב��Sta�tusՓ	Hea�rtbeatїMH Faul��Aler'�W�E� W�i�{ύϟϱ������� �CΛ�A�� ��8�J�\�n߀ߒߤ� �����������"�4��F�X�j�|���WOR {pΛ��(ߎ����� � �$�6�H�Z�l�~��� ������������ 2PƠ�X �� A{������ �/ASew������SDEV[�o�#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g?>y?PALTݠ1 ��z?�?�?�?�?O"O 4OFOXOjO|O�O�O�O��O�O�O�O_�?GRI�`ΛDQ�?_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|� ���������0�B�T��oPREG �>�� f���Ə؏� ��� �2�D�V�h�z� ������ԟ���Z���$ARG_��D ?	���;���  �	$Z�	[�O�]O��Z�p�.�S�BN_CONFIOG ;��������CII_SA_VE  Z������.�TCELLSETUP ;��%HOME_I�OZ�Z�%MOVq_��
�REP�l�U�(�UTOBAC�Kܠ���FRA:\z� �\�z�Ǡ'`�pz���ǡi�INI�0�z���n�MESSAG���ǡC�>��ODE_D����ą�%�O�4�n�PA�USX!�;� ((O>��Ϟˈ� �Ϭ���������� *�`�N߄�rߨ߶�g�~l TSK  w�x��_�q�UPDT+���d!�A�WSM�_CF��;����'�-�GRP 2�:�?� N�BŰA|��%�XSCRD1�;1
7� �ĥĢ����������*� ������r��������� ��7���[�&8J�\n��*�t�GR�OUN�UϩUP�_NA�:�	�t��_ED�1�7�
 �%-B?CKEDT-�2��'K�`���-(t�z�q�q�z���2t1�����q�k�(/��ED3/��/�.pa/�/;/M/ED4�/ t/)?�/.?p?�/�/ED5`??�?<?.p�?O�?�?ED6O �?qO�?.MO�O'O9OED7�O`O_�O.p�O\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o��_	-9o�oo%oCR_ 9]�oF�o�k� � NO_D�EL��GE_U�NUSE��LA�L_OUT �����WD_AB�ORﰨ~��pIT_R_RTN��|ONONSk����˥CAM_PAR�AM 1;�!�
� 8
SONY� XC-56 2�34567890� ਡ@����?��( С�\�
���{����^�HR5q�̹��ŏ�R57ڏ�Af�f��KOWA �SC310M
��x�̆�d @ <�
���e�^��П \����*�<��`��r�g�CE_RIA�_I�!�=�Ff��}�z� ���_LIU�]������<��FB�GP� 1��Ǯ��M�_�q�0�C* Y ����C1��9���@��G���CR�CU]��d��l��s��QR�����[Դm���v���������W C����(���숁=�HE�`ONF�Iǰ�B�G_PR/I 1�{V�� �ߖϨϺ�����������CHKPAUS��� 1K� , !uD�V�@�z�dߞ߈� ���߾������.��R�<�b���O���������_MOR��� ���B�Z?����� 	 �����*��N�`��������?��q?$;�;����K��9��P���çaÃ-:���	�

 ��M���pU�ð��<���,~��DB����튒)
mc:c?pmidbg�f~�:�  ���¥�p�/�O  �U�U�	s�� )� �s>_�  .�/UX�?��p#�pE$Ug�/���p�Uf�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����o=L���*MC��1����?43���1��t�īCz�  BHH�CPU�eB��CF��;.<C����C5rY
K�D��nyDQ��D���>��D�;D���=�F��>F�$�G}RB�7Gz�0��Y	��Y!�&w�1����s�������b���BDw�M@x8�ʊ1Ҩ����g@D��p@�0EYK�EX��EQ�EJ�P F�E�F�� G��>^�F E�� FB�� H,- Ge���H3Y��:��  >�33 s���~  n8�~@��5Y�E>�ðyA��Y<#�
"Q� ���+_�'RS/MOFS�p�.8���)T1��DE ���F 
Q��;�(P  B_<_���R����	op6C4RP�Y
s@ ]AQ��2s@C�0B3�MaCR{@@*cw��UT�p�FPROG %�z�o�oigI�q���v���ldKEY_TB�L  �&S�#� ��	
�� �!"#$%&'(�)*+,-./0�1i�:;<=>?�@ABC� GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�������������������s���p`LCK�lx4�p`�`STAT ���S_AUTO_D�O���5�IND�T_ENB!���R��Q?�1�T2}�^�S�TOPb���TRL^r`LETE��Ċ�_SCREEN ��Zkcs�c��U��MMEN�U 1 �Y  <�l�oR�Y1� [���v�m���̟���� �ٟ�8��!�G��� W�i��������ïկ ��4���j�A�S��� w�����迿�ѿ��� �T�+�=�cϜ�sυ� �ϩϻ�������P� '�9߆�]�o߼ߓߥ� �������:��#�p� G�Y��������� ��$����3�l�C�U� ��y����������� ���	VY)�_MA�NUAL��t�DB;CO[�RIGڇ
��DBNUM� ���B1 e
�PXWO_RK 1!�[�_�U/4FX�_�AWAY�i�G�CP  b=�Pj_CAL� #�j�Y���܅ `�_�  1">�[ , 
�m�g�&/~&lMZ�I�dPx@P@#ONT�IMه� d��`&�
�e�MOT�NEND�o�RECORD 1(�[qg2�/{�O��! �/ky"?4?F?X?�( `?�?�/�??�?�?�? �?�?)O�?MO�?qO�O �O�OBO�O:O�O^O_ %_7_I_�Om_�O�_ _ �_�_�_�_Z_o~_3o �_Woio{o�o�_�o o �oDo�o/�oS �oL�o����@ ���+�yV,�c� u��������Ϗ>�P� ����;�&���q��� 򏧟��P�ȟ�^�� ����I�[����� � ��$�6�������j�TOLERENC�wB���L���� CS_CFG �)�/'dM�C:\U�L%04�d.CSV�� cl��/#A ��CH��z� //.ɿ��(�S�RC_OUT �*��1/V�S�GN +��"���#�17-FE�B-20 18:�57027-JA}Np�21:48+ P;�����/.��f�pa��m��PJP�����VERSIO�N Y�V�2.0.�ƲEF�LOGIC 1,^� 	:ޠ�=�ޠL��PROG�_ENB��"p�U�LSk' ����_?WRSTJNK ���"fEMO_OPT_SL ?	��#
 	R575/#=�����0��B����TO  ��ݵϗ��V_F E�X�d�%��PA�TH AY�A�\�����5+ICTZ�Fu-�j�>#egS�,��STBF_TTS��(�	d���l#!w��� MAU��z�^"MKSWX�.�<�4,#�Y�/�
!J� 6%ZI~m��$�SBL_FAUL�(�0�9'TDIAb[�1<�<� ����123456�7890
��P ��HZl~��� ����/ /2/D/�V/h/�� P� ѩ�yƽ/��6�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�?��,/�UMP���� �ATR���1O�C@PMEl�OOY_�TEMP?�È��3F���G�|DUNI���.�YN_BRK� 2_�/�EMG?DI_STA��]���ENC2_SCR 3�K7(_:_ L_^_l&_�_�_�_�_)��C�A14_�/o@o/oAoԢ�B�T5�K�ϋo~ol�{_ �o�o�o'9K ]o������ ���#�5��/V�h� z��л`~�����ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T���x��� ������ү����� ,�>�P�b�t������� ��ο����(�f� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��:� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ���������* <N`r���� ���&8J \n�������� ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? ��?�?�?�?�?OO ,O>OPObOtO�O�O�O��O�O�O�O__NoE�TMODE 16v�5�Q �d��X
X_j_|Q�PR�ROR_PROG7 %GZ%�@��_�  �UTABLE  G[�?oo�)oRjRRSEV_?NUM  �`WP��QQY`�Q_�AUTO_ENB�  �eOS�T_N�Ona 7G[�Q�Xb  *��`�J�`��`��`d`+�`p�o�o�o�dHISUc��QOP�k_ALM �18G[ �A��l�P+�ok}������o_Nb�`  G[�a�R
�:P�TCP_VER �!GZ!�_�$E�XTLOG_RE�Qv�i\�SI�Ze�W�TOL  ��QDzr�=�#דQXT_BW�D�p��xf́t�_D�I�� 9�5��d�T�QsRֆSTE�P��:P�OP_�DOv�f�PFA�CTORY_TU�NwdM�EATU�RE :�5̀�rQHand�lingTool� �� \sfm�English� Diction�ary��rodu�AA Vis��� Master�����
EN̐n�alog I/O�����g.fd̐u�to Softw�are Upda�te  F OR��matic B�ackup��H5�96,�gro�und Edit�ޒ  1 H5Camera�F��OPLGX�e�ll𜩐II) nX�ommՐshw�n��com��co����\tp���pa�ne��  opl���tyle se�lect��al �C��nJ�Ցoniwtor��RDE���tr��Reli�ab𠧒6U�Diagnos(�푥��5528�u��h�eck Safe�ty UIF��E�nhanced �Rob Serv>%�q ) "S�r�User Fr[������a��xt. oDIO �fiG�s sŢ��endx��Err�LF� p$Ȑĳr됮� �����  !��FCTN_ Menu`�v-��ݡ���TP In�ېfac�  E�R JGC�p�בk Exct�gޠ�H558��ig�h-Spex�Sk�i1�  2
P���?���mmunic'�ons��&�l��ur�ې��ST xǠ��conn���2��TXPL��n{cr�stru�����"FATK�AREL Cmd�. LE�uaG�5�45\��Run-�Ti��Env��dG
!���ؠ++��s)�S/W��[��License�Z��� 4T�0�ogBook(Syڐ�m)��H54O�M�ACROs,\�/�Offse��Lo�a�MH������r�, k�MechS�top Prot����� lic/�M=iвShif����ɒMixx��)����xSPS�Mode Switch��7 R5W�Mo�:�=.�� 74 ����g��K�2h�ul�ti-T=�M���L�N (Pos�Regiڑ�������d�ݐt Fun��ǩ�.�����Nu�m~����� lne���ᝰ Adju�p�����  - =W��tatuw᧒}T�RDMz��ot��scove
 U�9���3����uest 49�2�*�o�����62~;�SNPX b Ҟ��8 J7`���Lgibr��J�48��D�ӗ� �Ԅ�
�6O��� Parts in VCCMt�32���	�{Ѥ�J�990��/I� �2 P��TMILKIB��H���P��AccD�L�
T�E$TX�ۨ�ap�1S�Te����pkCey��wգ�d���Unexce{ptx�motnZ�0�������є��� O���� 90�J�єSP CSX�C<�f��Ҟ� P�y�We}���PRI��>vr�t�me�n�� ��iP�ɰa�����vGr{id�play�İv��0�)�H1�M�-10iA(B2�01 �2\� 0�\k/�Ascii��l�Т�ɐ/�Coyl��ԑGuar�� 
�� /P-�ޠ"�K��st{Patt ��!S�Cyc�҂�orie��I�F8�ata- qu�Ґ�� ƶ��mH5�74��RL��am����Pb�HMI �De3�(b����P�CϺ�Passw�o+!��"PE? S1p$�[���tp��� �ven��Tw�N�p��YELLOW sBOE	k$Arc��'vis��3*�n0�WeldW�cia�l�7�V#t�Opd����1y� 2F�=a�portN�(�p�T1�T� �� f��xy]�&TX��tw�igj�1� b�� ct\�JPN� ARCPSU cPR��oݲOL� wSup�2fil� p&PAɰאcro�� "PM(����O$�SS� eвtexF�� r���=�t�OssagT��P���P@�Ȱ�锱�r�tW��H'>r�dp9n��n1
t�!� z ��ascbin4psyn���+Aj�M HEL��NCL VIS� PKGS PL;OA`�MB �,��4VW�RIPE� GET_VAR� FIE 3\t���FL[�OOL:� ADD R72�9.FD \j8�'�CsQ�QE��DV�vQ�sQNO WT�WTE��}PD  �^��biRFOR ��ECTn�`���ALSE ALA�fPCPMO-130  M" #h��D: HANG �FROMmP�AQf�r��R709 D�RAM AVAILCHECKSO!���sQVPCS S�U�@LIMCHK� Q +P~dFF P�OS��F�Q R5�938-12� CHARY�0�P?ROGRA W��SAVEN`AME.�P.SV��7��$�En*��p?FU�{�T�RC|� SHAD�V0UPDAT K�CJўRSTATI��`�P MUCH �y�1��IMQ MOTN-003���}�ROBOGUI�DE DAUGHp�a���*�tou�����I� Šhd�AT�H�PepMOVET��ǔVMXPAC�K MAY AS�SERT�D��YC�LfqTA�rBE ?COR vr*Q3r�AN�pRC OP�TIONSJ1vr�̐PSH-171ZZ@x�tcǠSU1��1Hp^9R!�Q�`_TP�P��'�j�d{t�by app w�a 5I�~d�PHI����p�aTEL�MXSPD TB5b�Lu 1��UB6@�qEmNJ`CE2�61���p��s	�may 1n�0� R6{�R�} �Rtraff)��� 40*�p��f�r��sysvar scr J7��cj`DJU��bH� V��Q/�PSET� ERR`J` 6�8��PNDANT� SCREEN UNREA��'�J`MD�pPA���pR`�IO 1���PFI��pB�pGROUN�PD��G��R�P�QnRSVIP !p�a�P�DIGIT VE�RS�r}BLo�UE�Wϕ P06  �!��MAGp�ab�ZV�DI�`� S�SUE�ܰ�EP�LAN JOT` 'DEL�pݡ#Z�@=D͐CALLOb�Q� ph��R�QIP�ND��IMG�R�719��MNT/��PES �pVL�c��Hol�0Cq���t�PG:�`C�M�c�anΠ��pg.v~�S: 3D mK�view d�` L�p��ea7У�b� �of �Py���AN�NOT ACCE�SS M��Ɓ*�tn4s a��lok�^�Flex/:�Rmw!mo?�PA?��-�����`n�pa �SNBPJ AUTO-�06f����T|B��PIABLE1q� 636��PLN�: RG$�pl;pNnWFMDB�VI��>�tWIT 9x�0@o��Qui#0�ҺP�N RRS?pUS�B�� t & r/emov�@ )�_�v�&AxEPFT_=�� 7<`�pP:�O�S-144 ��h� s�g��@OST�� � CRASH� DU 9��k$P�pW� .$��_LOGIN��8&��J��6b046 i�ssue 6 J�g��: Slow� �st��c (�Hos`�c���`I�L`IMPRWtSPOT:Wh:0�T��STYW ./�VM�GR�h�T0CAT.��hos��E�q�T�� �O�S:+p�RTU' k�-S� ,����E:��pv@�2��� t\hߐ��m� ��all��0� 9 $�H� WA͐���3 CNT0 T��� WroU�al�arm���0s�d �� �0SE1���r R{�OMEBp���K�7 55��REàSE�st��g   �  �KANJI��no���INISITALIZ-p��dn1weρ<��d�r�� lx`�SC�II L�fai/ls w�� ��`�YSTEa���o��PNv� IIH���1W��Gro>Pm ol\wpSh@�P��Ϡ?n cflxL@А�WRI �OF Lhq��p?�F�up��de-rela�_d "APo SY��ch�Abetwe>:0IND t0$FgbDO���r� `��GigE�#op�erabilf  �PAbHi�H`��c�l�ead�\etfp�Ps�r�OS 0�30�&: fig��GLA )P ��i��}7Np tpswx�-B��If�g�������5aE�a EX�CE#dU�_�tPCL{OS��"rob�+NTdpFaU�c�!����PNIO V750�Q1��QaN��DB ��P M��+P�QED�DET���-� \rk��O�NLINEhSBU�GIQ ߔĠi`Z�I�B�S apABC? JARKYFq�9 ���0MIL�`� �R�pNД �p0G+AR��D*pR��PN�"! jK�0cT�P�Hl#n�a�ZE }V�� TASK�$VP2(�4`
�!�$��P�`WIBPK0�5�!FȐB/��B�USY RUNN��� "�򁐈��R�-p�LO�N�DI�VY�CUL��f3sfoaBW�p����30	V��ˠIyT`�a505.�@{OF�UNEX�P�1b�af�@�E��S�VEMG� NML�q� D0pCC_SGAFEX 0c�08"q]D �PET�`N@N�#J87����RsP��A'�M�K�`K��H GUNCH�G۔MECH�pM�c� T�  y, �g@�$ ORY L�EAKA�;�ޢS�PEm�Ja��V�tG�RIܱ�@�CTLN�TRk�FpepnR�j50�EN-`#IN�����p �`�Ǒk!��T3/dqo��STO�0A�#�L��p �0�@�Q�АY0�&�;pb1TO8pP�s���FB�@Yp`�`DU��aO�supk��t4 � P�F� Bn�f�Q�PSVGN-q1��V�SRSR)J�UP�a2�Q�#D��q l O��QBRKCTR5Ұ�|"�-�r�<pc�j!IN=VP�D ZO� ���T`h#�Q�cHset�,|D��"DUAL�� w�2*BRVO1/17 A]�TNѫt8�+bTa2473��q.?��sAUz�i�B��complete���604.� �-�`hanc�U�� F��e8�� 	 ��npJtPd!q��`���� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP���R(}\xPe� aʰI���E��1��p�� j  �� xSP�'^P �A�AxP�q\ 5 sig��a��"AC;a��
�b�CexPb_p��.p�c]l<bHbcb_c�irc~h<n�`tl 1�~`xP`o�dxP�b]o2�� �cb�c�ixP>�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`>�cptlibxzxP�lcr�xrxP\�b�lsazEdxP_fm �}gcxP�x���o|sp��o�mc(��ob_jDzop�u6�wf���t��wms�1q��s1ld�)��jmc�o\��n��nuhЕ��|st�e��>�pl�qp�iwcck���uvf0uxߒ��lvisn��CgaculwQ
E� F  ! Fc.sfd�Qv�� qw����Data Ac_quisi��nF�<|1�RR631`��T}R�QDMCM ��2�P75H�1�P5k83xP1��71��k59`�5�P57<P xP�Q����(���Q̖�o pxP!da�q\�oA��@��y ge/�etdms�?"DMER"؟,�GpgdD���.�m��8�-��qaq.<᡾FxPmo��h���f{��u�`13��MACR�Os, Sksaf�f�@z����03�SR��Q(��Q6��1�Q9�ӡ�R�ZSh��PxPJW643�@7ؠ6�P,�@�PRS�@���e x�Q�UС PIK�Q52 PTLC�W���xP3 (��p/O��!�Pn �xP�5��03\sfm�nmc "MNM�Cq�<��Q��\$AcX�FM���ci,Ҥ��X����cdpq+�
�s�k�SK�xP�SH560,P��,�y��refp "RE�Fp�d�A�jxP	�o�f�OFc�<gy�to�TO_����ٺ���+je�u��caxis2�xPE��\�e�q"ISDT�c��]�prax ���MN��u�b�isde܃h�\�w�xP�! isbasi5c��B� P]��QoAxes�R6��8����.�(Ba�Q�ess��xP����2�D�@�z�atis ���(�{�����~��m��FMc�u�{�<
ѩ�MNIS��ݝ ����x����ٺ���x� j75��De�vic�� Interfac�RȔQJ754��� xP�Ne`��xP�ϐ`2�б����dn� �"DNE���
t�pdnui5UI��ݝ	bd�bP>�q_rsofOb~
dv_aro��u�����stchkc��z	 �(�}onl��G!ffL+H�J(��"l"�/�n�b��z�h�amp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!�2��xpc_2pcc{hm��CHMP_�|8бpevws��2�쳌pcsF��#C� SenxPacrao�U·�-�R6�P�d�xPk�����p��g8T�L��1d M�2`���8�1c4ԡ�3 qem��GEM,\i(�>�Dgesnd�5��`�H{�}Ha�@sy����c�Isu�xD��Fmd��I��7�4���u����AccuCal �P�4� ��ɢ7ޠBU0��6+6f�6��C99\aFF q�S(�U��2�
X�p�!Bdf��cb_�SaUL��  �� ?�ܖt�o��otplus\tsrnغ�qb��Wp��t���1��T�ool (N. �A.)�[K�7�Z�(P�m����bfc�ls� k94�"Kp4p��qtpap�� "PS9H�stpswo��p�L7��t\�q����D�yt 5�4�q��w�q��� ��M�uk��rkey�����s��}t�sfoeatu6�EA��� cf)t\Xq�����̜d�h5���LR0C0�md�!�587���aR�(����2V���8c?u3l\�pa�3}H�&r-�Xu���t,�� �q "�q�Ot� �~,���{�/��1c�}����y�p�r��5� ��S�XAg�-�y���W�j874�- i�RVis���Queu�� Ƒ�-�6H�1���(����u����tӑ����
�tp�vtsn "VTCSN�3C�+�� v\p�RDV����*�pr�dq\�Q�&�vs�tk=P������n�m&_�դ�clrq8ν���get�TX��Bd���aoQϿ�0qstr�D[� ��at�p'Z����npv��@�enlIP0��`D!x�'�|���sc ����tvo/��2�q���vb����q ���!���h]��(�� Control^�PRAX�P5��g556�A@59�P[56.@56@5A��J69$@982� J552 IDVR7�hqA���16��H���La�� ���Xe�frlpa�rm.f�FRL��am��C9�@(F�����w6{���A<��QJ643�� �50�0LSE
�_pVAR $SG�SYSC��RS_?UNITS �P�2��4tA�TX.$V�NUM_OLD �5�1�xP{�50�+�"�` Funct���5tA� }��`#@��`3�a0�cڂ��9���@H5נ� �P���(�A����۶�}����ֻ}��bP�Rb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`��2�1���96����@�%C�� Aف��J�bIncr�	����\����1o5qni4�MNINp	xP�`���!��Hour�  � �2�21 ��AAVM���0y ��TUP ��J545 ���6162�V�CAM  (��CLIO ���R6�N2�MS�C "P ��STYL�C�2�8~ 13\�NRE "FHRM �SCH^�DC�SU%ORSR �{b�04 �oEIOC�1 j o542 � os| ~� egist������7�1��MASK�93�4"7 ��OCO) ��"3�8��12���� 0 HB���� 4�"39N� �Re�� �LCH=K
%OPLG%��3"%MHCR.%M�C  ; 4? ��6 6dPI�54�s� �DSW%MD� pQ�K!637�0�0p"��1�Р"4 �6~<27 CTN K V� 5 ���"7���<25�%/�T�%FRDM� �Sg!���930 FB( NB�A�P� ( HLB o Men�SM$@<jB( PVC ��s20v��2HTC�~CTMIL��~\@PAC 16U��hAJ`SAI \@EL�N��<29s�U�ECK �b�@FR3M �b�OR����IPL��Rk0CS�XC ���VVF�naTg@HTTP ��!26 ��G��@obIGUI�"%IPGS�r� H863 qb�!�07rΈ!34 �r�84 \so`! Qx`CC�3 Fb�21�!9s6 rb!51 ����!53R% 1!s(3!��~�.p"9js �VATFUJ775�"��pLR6^RP�W;SMjUCTO�@xT158 F!80���1�XY ta3!770� ��885�UO	L  GTSo
�{` �LCM �r| TS�S�EfP6 W�\@C�PE `��0VR�� l�QNL"��@001 imrb�c3 =�b�0���0�`�6 w�b-P- Ru-�b8n@5EW�b9 �Ґa� ���b�`�ׁ�b2 2000$��`3��`4*5�`A5!�c�#$�`7.%~�`8 h605? ;U0�@B6E"aRpm7� !Pr8 t��a@�tr2 iB�/�1vp3�vp5 �Ȃtr9Σ�a4@-�p�r3 F��r5`&�re`u��r7 ��r8�U�p9 \h�738�a�R2DK7"�1f��2&�y7� �3 7iCЊ�4>w5Ip�Or6�0 C�L�1bEN�4 I�pyL�uP��@LN�-PJ8�N�8Ne�N�9 H�r`�E"�b7]�|���8�В����9 2��a`0�qЂ5�%U097 0��@1�0����1 (�q�3 5R���0���mpU��0�0�7*�H@x(q�\P"RB6�q124�b;��@���f@06� x�3 p�B/x�u ��x�6 /H606�a1� ����7 6 ���<p�b155 ����}7jUU162 ��3 g��4*�6?5 2e "_��PF�4U1`���B1��z�`0'�174 �q���P�E186 R� ��P�7 ��P�8�&�3 (�90 B/�s191����@�202��6 30���A�RU2� d���2 b2h`��4Ģ᪂2�4���19�v Q�2��u2d�TRpt2� ��H�a2hPd�$�5���!U2�pD�p
�2�p��@5�0H-@��8 @�9��TX@�� �e5�`rb26Af�2^R�a�2 Kp��1y�b5Hp�`

�5�0@�gqGA��F�a52ѐ�Ḳ6�K60ہ5� ׁ2��i8�E��9�EU5@�ٰ\�q5hQ`S�2
ޖ5�p\w�۲�pJh �-P��5�p1\t�ZH�4��PCH�7j��phiw�@��P�x�~�559 ldu�  P�D���Q�@�������� �`.��P>��8��581�"�q58�!AM۲T�A iC�a589��@�x�����5 �a��12@׀0.�1���,�2��8��,�!P\h8��Lp� ��,�7��6�08�40\��ANRS 0C}A��p��{��ran��FRA ��Д�е���A% ���ѹ�Ҍ�����( ����Ќ���З��� ������ь����$�!G��1��ը���������� xS�`q�  �����`�64��M��iC/50T-H������*��)p46��� C���N����m75s�֐� Sp��b4�6��v����ГM-71?�7�З�����42������C��-��а�70�r�E��/h����O$���rD���c7c7C@�q��Ѕ���L���/��2\imm7c7�g������`���(��e����� "�������a r�L�c�T,�Ѿ�"��,�� ��x�Ex�m77t����k���a5�����)�iC��-HS-� B
_�@>���+�Т�7U��]���Mh7�s�7������-9~?�/260L_� �����Q������4��]�9pA/@���q�S�х鼔��h621��c��92������.�)92c0�g$�@ �����)$��5$����pylH"O"
�21p���t?�350� ���p��$�
��� �350!���0���9�U/0\m9��M9A3��4%� s��3M$��X%yu���"him98 J3����� i d�"m4~�103p�� ����h794̂�&R���H�0����\���g� 5AU��՜��0���*2@��00��#06�`�АՃ�է!07{r ��������kЙ @����EP�#�� ����?��#!�;&�07\;!�B1P��߀A��/ЁCBׂ2��!�:/��?�ҽCD2C5L����0�"l�2BL
#��B��\20�2_�r�re ���X��1��N����A$@��z��`C�p0U��`��04��DyA�\�`fQ����sU���\�5  ���� p�^P��<$85���+�P=�ab1l��1LT��lA8�!uDnE\(�20T��J�1 e�bH85���b����5[�16Bs��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3� � ��b�s��-`�_�Wa8�_����6I	$2�X5�1�U85��R�p6S����/�/+q��!�q��`�6o��58m[o)�m6sW��Q��?��set06�p ��3%H�5��10�p$����g/�JrH~��  ��A�856����F�� ���p/2��h�܅�✐)�5��̑v0��(��m6��Y�!H�ѝ̑m�6�Ҝ���a6�DM����-S�+��H2������ ��� �r̑��✐0��l���p1���Fx���2�\t6h T6H����Ҝ�'V l���ᜐ�V7ᜐP/����;3A7��@p~S��������4�`@圐�V���!3��2�PM[��%ܖO�7chn��vel5�p���Vq���_arp#���̑�.���2l_�hemq$�.�'�6415���5���?�� ��F�����5g�L�ј[���1��𙋹y1����M7NU�@�М��eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h����� �u���㜐��`ZS�!ܑ4���M-����S�$̑�ք �� �0��<�����07shJ�H�v�À�sF ��S*󜐳���̑�� �vl�3�A�T�#��`QȚ�Te��q�pr��,��T@75j�5�dd� ̑1�(UL�&�(�,����0�\�?���̑�a��? xSP���a��e�w�2��(�	�2�C��A/���\�+px�����21 (ܱ�CL S����B�̺��7F���?�<�lơ1L����c� ��b�u9�0����e/q���O���9�K��r9 (��,�Rs�ז�x5�G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O����1!41w���2<T@� _std��G��y� �ң�H� jdgm����w0\� �1 L���	�P�~�W*�b��t 5������%3�,���E{�������L��5\L��3�L�|#~���~!���4�#��O����h�L6A������2璥���44������[6\j4s��·���#��ol�E"w�8Pk�����?0 xj�H1�1Rr�>��6]�2a�2Aw�P ��2��|41�8��ˡ���{� �%�A<���  +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R� �ˑb�W���Fs��� �)�ѐ�!���a�1��ڛ�5��16�16�C��C����0\imBQ��d����b���\B5�-���DiL ���O�_�<ѠPEtL�E�RH�ZǠPgω�am1l��u���̑��b�<����<�$�T �̑�F����Ȋ�D�pb��X"��hr��pw� ���^P���9�0\� j971\kckrcfJ��F�s�����c��e "CTME�r��������a�`main.p[��g�`run}�_vc�#0�w�1O�ܕ_u����bctm�e��Ӧ�`ܑ�j7�35�- KAREL Use {�	U���J��1��
�p� Ȗ�9�B@���L�9��7j[�a�tk208 "KP��Kя��\��9���a��̹����cKRiC�a�o ��kc�q J�&s�����Grſ� fsD��:y��s�ˑ1X3\j|хrdtB�,� ��`.v�q�� ��sǑIf�Wfj52��TKQuto S�et��J� H5nK536(�932�Z��91�58(�9�BA�1(�74O,A$�?(TCP Ak��В/�)Y� �\t�pqtool.v��v���! co�nre;a#�Control Re��ble��CNRE (�T�<�4�2���D�)����S�552��q(g�� (򭂯4X�cO�ux�\sfuts�UTS`�i�栜����t�棂��? 68�T�!�SA OO+D6���������,!��6c+� ig.t�t6i��I0�TW8 ���la��vo58�o�bFå򬡯i�Xh��!Xk�0Y!�8\m6e�!6EC���v��6���������<16�A���A�6s����U�g�TX|ώ���r1�qR��˔Z4�T�����,#�eZp)g����<O NO0���uJ��tCR;�x�F�a� xSP�f���prdsuchk �1��2&&?���	t��*D%$�r(��@���娟:r��'�s�q8O��<scrc�C�<\At�trldJ"�o�\�V����Pa�ylo�nfir1m�l�!�87��7� �A�3ad�! ��?ވI�?plQ��3���3"�q��x p�l�`���d7��l�calC�uDu���;���mov�����i'nitX�:s8O�p�a�r4 ��r67A4�|�e GenerGatiڲ���7g2�q$��g R� (#Sh��c ,|�bE��$Ԓ\�:�"��4��4�4�. sg��5�F$d6�"e;Qp "SH�AP�TQ ngcr pGC�a(�&"<� ��"GDA¶��r6�"aW�/�$�dataX:s�"t�pad��[q�%tput;a__O7;a�o8(�1�yl+s�r�?�:H�#�?�5x�?�:c O��:y O�:�IO�s`O%g�qǒ�?�@08\��"o�j92;!�P�pl.Colli=s�QSkip#��@ 5��@J��D��@\ވP�C@X�7��7��|s2��ptclsF�LS�DU�k?�\_ ets�`�< \�Q��@���`dc�KqQ�FC;��J,�n��` (��4eN����T�{��� 'j(�c�����/IӸaxȁ��̠H������зa�e\mc�clmt "CL�M�/��� mate�\��lmpALM0�?>p7qmc?����2vm�q��%�3s���_sv90�_x_m#su�2L^v_� K�o�{in�8(3r<�c_logr�N�rtrcW� �v_3�~yc��d��<�te��derv$cCe� Fiρ�R��Q�?�l�enter߄|��d(Sd��1�TX�+�fK�r�a99sQ9x+�5�r\tq\�� "FNDR����STDn$�LANG�Pgui��D⠓�S����Ơ�sp�!ğ֙uf �ҝ�s����$�����e+�=����������ࠓ���w�H�r\f�n_�ϣ��$`x�tc�pma��- TC�P�����R638� R�Ҡ��38
��M7p,���Ӡ�$Ӏ��8p0Р�VS,�>�tk��99�a��B3�� �PզԠ��D�2�����UI��t���hqB���8��������p���rqe�ȿ��exe@ 4φ�B���e38�ԡG��rmpWXφ�var@�φ�3N������vx�!ҡ��q��RBT $cO�PTN ask �E0��1�R MA�S0�H593/�9�6 H50�i�48
0�5�H0��m�Q�QK��7�0�g�Pl��h0ԧ�2�ORD�P��@"��t\mas��0�a��"�ԧ�����k�գR�����¹`m��b��7�.f���u�d��r��splayD�E���1>w�UPDT Ub���887 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q `�䗣�#��К�`2�� vlv��Ù�`$�>�b���! S���Easy/К�U�til��룙�51G1 J�����R7 Θ�Nor֠��inGc),<6Q�� �`�c��"4�[���98Q6FVRx So����q�nd6����P�� 4�a\ (��
  ����D���d��K�bdZ����men7���- Me`tyFњ�Fb¨0�TUa�57	7?i3R��\��5�u?��!� n����f������l\mh�Ц�űE|Ghmn�	��<\HO���e�1�� l!D��y��Ù�\|�p����B���Ћmh�@��:.aG! ���/�t�55�6�!X�l�.us��Y/k)�ensubL���eK�h�� �B\1;5�g?y?�?�?D��?*r�m�p�?Ktbox  O2K|?�G��C?A%�ds���?1ӛ#�  �TR��/��P�4B�`��U�P�V�P"�Q�P0@�U�PO��P�"�T3�U@�P�f�Pk"�2}�4�T@�P�f�P2�"�Q5�S��Q���R?Ă�Q3t.��P׀al��P+O�P517��IN�0a��Q(}g��PESTf3ua�PB�l��ig�h�6�aq��P? � xS��`�  n�0mbum�pP�Q969g�6!9�Qq��P0�baAp|�@Q� BOX��,>vche�s�>v�etu㒣=wffse�3���]�;u0`aW��:zol�sm�<ub�a-��]D�K�ibQ�c����Q<twaǂ� tp�Q҄Tar�or Recov�b�O�P�642 ����a�q��a⁠Q3Erǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>�pjot��PXc���C�1�adb -�ail��nag���b�QR629�a�Q��b��P  �
�  �P��$$C�L[q ���t������$�PS_DIGIT�.��"�!� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv��������*璬1:PRODUCT�Q0\PGSTK�bqV,n�99��\���$FE�AT_INDEX���~��� 搠ILECO_MP ;��)���"��SETU�P2 <�~��  N !��_AP2BCK� 1=�  #�)}6/E+%,/i/��W/�/~+/�/ O/�/s/�/?�/>?�/ b?t??�?'?�?�?]? �?�?O(O�?LO�?pO �?}O�O5O�OYO�O _ �O$_�OH_Z_�O~__ �_�_C_�_g_�_�_	o 2o�_Vo�_zo�oo�o ?o�o�ouo
�o.@ �od�o���M �q���<��`� r����%���̏[��� ����!�J�ُn��� ����3�ȟW������ "���F�X��|���� /���֯e������0� ��T��x������=� ҿ�s�ϗ�,ϻ�9��b�� P/ 2>) *.VRiϳ�!�*�������ߌ��PC�7�!�OFR6:"�c������T��߽�Lը���ܮx���*.F��>� �	N�,�k���ߏ��STM @�����Qа���!��iPendant Panel���H��F���4�������GIF��������u����JPG &P��<�����	PANEL1.DT��������2�Y�G��
3w�� ���//�
4�a/��O///�/�
T�PEINS.XM)L�/���\�/�/��!Custom Toolbar?��PASSWO�RD/�FRS�:\R?? %P�assword ?Config�?� �?k?�?OH�6O�?ZO lO�?�OO�O�OUO�O yO_�O�OD_�Oh_�O a_�_-_�_Q_�_�_�_ o�_@oRo�_voo�o )o;o�o_o�o�o�o* �oN�or��7 ��m��&��� \�����y���E�ڏ i������4�ÏX�j� �������A�S��w� ����B�џf����� ��+���O������� ��>�ͯ߯t����'� ��ο]�򿁿�(Ϸ� L�ۿpς�Ϧ�5��� Y�k� ߏ�$߳��Z� ��~�ߢߴ�C���g� ����2���V����� ����?����u�
� ��.�@���d������ )���M���q����� <��5r�%� �[�&�J �n��3�W ���"/�F/X/� |//�/�/A/�/e/�/ �/�/0?�/T?�/M?�? ?�?=?�?�?s?O�? ,O>O�?bO�?�OO'O �OKO�OoO�O_�O:_ �O^_p_�O�_#_�_�_ Y_�_}_o�_�_Ho)f��$FILE_D�GBCK 1=���5`��� ( �)
�SUMMARY.�DGRo�\MD:�o�o
`Dia�g Summar�y�o�Z
CONSLOG�o�o�a
J��aConsol�e logK�[��`MEMCHEC�K@'�o�^qM�emory Da�ta��W�)}�qHADOW���P��sSha�dow Chan�gesS�-c-�?�)	FTP=���9����w`qmme?nt TBD׏�W�0<�)ETHERNET̏�^�q��Z��aEthe�rnet bpfi�guration�[��P��DCSVR�Fˏ��Ïܟ�q%��� verif�y allߟ-c1�PY���DIFF�ԟ��̟a��p%��diffc���q¡�1X�?�Q�� �����X��CHGD��¯ԯi��p!x��� ���2`�G�Y�� ��� ��GD��ʿܿq��p8���Ϥ�FY3h�O�a��� ��(σGD������y��p��ϡ�0�UPDA�TES.�Ц��[�FRS:\������aUpdates� List���kP�SRBWLD.C	M.��\��B��_p�PS_ROBOWEL���_����o�� ,o!�3���W���{�
� t���@���d����� /��Se���� �N�r� = �a�r�&�J ���/�9/K/� o/��/"/�/�/X/�/ |/�/#?�/G?�/k?}? ?�?0?�?�?f?�?�? O�?OUO�?yOO�O �O>O�ObO�O	_�O-_ �OQ_c_�O�__�_:_ �_�_p_o�_o;o�_ _o�_�o�o$o�oHo�o �o~o�o7�o0m �o� ��V�z �!��E��i�{�
� ��.�ÏR�������� ��.�S��w������ <�џ`������+��� O�ޟH������8����߯n����$FI�LE_��PR����������� �MDON�LY 1=4�� 
 ���w�į ��诨�ѿ������� +Ϻ�O�޿sυ�ϩ� 8�����n�ߒ�'߶� 4�]��ρ�ߥ߷�F� ��j�����5���Y� k��ߏ���B����� x����1�C���g��� ����,���P����������?��Lu�VISBCKR�<�a�*.VD|�4 �FR:\���4 Vision� VD file � :LbpZ� #��Y�}/$/ �H/�l/�/�/1/ �/�/�/�/�/ ?�/1? V?�/z?	?�?�???�? c?�?�?�?.O�?ROdO O�OO�O;O�O�OqO _�O*_<_�O`_�O�_�_%_�_�MR_G�RP 1>4��L�UC4  B��P	 ]�ol`��*u����RHB ��2� ��� ��� ���He�Y�Q`o rkbIh�oJd�o�Sc��o�oL,�M�V`KGXF��5U�aS����o�o E=�aEP��E!��-���9?6�">_Z`}@�6�A�j0lq?_��A�e�xq�0~�� F@ �r�d�a}J��N�Jk�H9��Hu��F!��/IP�s}?�`��.9�<9���896C'�6<,6\b ~+A�,�e�P���t�A�PA�����|�ݏ x���%��I�4�F� �j�����ǟ���֟���!��E�`r�UBH�P �~��������W
6�PJ��PQ��˯�o�o�B��P5���@�3�3@���4�m�T�U�UU��U�~w�>u?.�?!x�^���ֿ���3��=[�z�=�̽=�V6<�=�=��=$q��~���@8�i7G���8�D�8?@9!�7ϥ��@Ϣ���cD�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p������������� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__/  D�UPE_�Hly_�\@@m_B�=��vR/��I�O�SMT*�G���
�o�o+l�$HOST�C�1H�I� Ĺ�zMSM��l[bo�	1�27.0�`1�o  e�o�o�o #z�oFXj|�l6�0s	anonymous�����F�%ao�&�&��o�x��o������ ҏ�3��,�>�a� O����������Ο�U %�7�I��]����f� x��������ү��� �+�i�{�P�b�t��� ���������S� (�:�L�^ϭ�oϔϦ� �������=��$�6� H�Zߩ���Ϳs����� ������ �2���V� h�z��߰������� ��
��k�}ߏߡߣ� ���߬���������C� *<Nq�_�� ����-�?�Q�c� eJ��n���� ���/"/E� X/j/|/�/�/� %'/?[0?B?T?f? x?��?�?�?�?�?? E/W/,O>OPObO�KDa�ENT 1I�K� P!�?�O  �P�O�O�O�O�O#_ �OG_
_S_._|_�_d_ �_�_�_�_o�_1o�_ ogo*o�oNo�oro�o �o�o	�o-�oQ u8n����� ���#��L�q�4� ��X���|�ݏ���ď�֏7���[���B�?QUICC0��h�z�۟��1ܟ��ʟ+��2,���{�!?ROUTER|�X��j�˯!PCJO�G̯��!19�2.168.0.�10��}GNAME� !�J!RO�BOT�vNS_C�FG 1H�I ��Aut�o-starte�d�$FTP�/ ���/�?޿#?��&� 8�JϏ?nπϒϤ�ǿ ��[������"�4�G�#������������ �����������&�8� J�\�n������� ������/�/�/F��� j��ߎ����������� ��0S�T��x �����!�3�� G,{�Pbt�� C����/� :/L/^/p/�/��� 	/�/=?$?6?H? Z?)/~?�?�?�?�/�? k?�?O O2ODO�/�/ �/�/�?�O�/�O�O�O 
__�?@_R_d_v_�_ �O-_�_�_�_�_oUO gOyO�O�_ro�O�o�o �o�o�o�_&8 Jmo�o����� o)o;oMoO!��oX� j�|�����oď֏� ���/���B�T�f�x����^�ST_ERR� J;�����PDUSIZ  ���^P����>ٕW�RD ?z����  guest���+�=�O��a�s�*�SCDMN�GRP 2Kz�;Ð��۠�\��K�� 	P01.14 8�q�   y���B    �;����{ ����������������������~ �ǟI��4�m�X�|�� � i  � � 
���� �����+��������
���l�.Vx����"�l�ڲ۰s�d��������_GROU��L.�� ��	��۠�07K�QUPD � ���PČ�T�Yg�����TT�P_AUTH 1�M�� <!i?Pendan����<�_�!KAREL:*����݇KC%�5�G���VISION SCETZ���|��� �ߪ���������
�W�.�@��d�v���C?TRL N��������
�FF�F9E3���F�RS:DEFAU�LT�FAN�UC Web S_erver�
�� ����q��������������WR_CON�FIG O�� ����IDL_�CPU_PC"���B��= �BH�#MIN.�BGNR_IO��� ����% NPT_SI�M_DOs}T�PMODNTOL�s �_PRTY��=!OLNK 1P���'�9K]o�MAS�TEr �����O_gCFG��UO��|��CYCLE����_ASG 19Q���
 q2/ D/V/h/z/�/�/�/�/��/�/�/
??y"N�UM���Q�I�PCH��£RTRY_CN"�u���SCRN������� ���R���?��$J2�3_DSP_EN������0OBP�ROC�3��JO�GV�1S_�@��8�?�';ZO'?}?0CPOSREO~�KANJI_� Ϡu�A#��3T ����E�O�ECL_L�M B2e?�@EYLO�GGIN��������LANGUA�GE _�=�� }Q��LG�2U������ �x������PC � �'0������MC�:\RSCH\0�0\˝LN_DISP V��������TOC�4D�z\=#�Q�?PB?OOK W+��`o���o�o���Xi��o�o�o�o�o~}	x(y��	ne�i��ekElG_BUF/F 1X���}2����Ӣ��� ���'�T�K�]��� ��������ɏۏ����#�P��ËqDCS� Zxm =���%|d1h`���ʟܟ|�g�IO 1[+G �?'����'� 7�I�[�o�������� ǯٯ����!�3�G� W�i�{�������ÿ׿z�El TM  ��d��#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝߜ�t�SEV�0m.�TYP�� �0�$�}�ARS"�(_|�s�2FL 1\��0���������0�����5�TP<P����DmNGNA�M�4�U�f�UPSF`GI�5�A�5s��_LOAD@G �%j%@_M�OV�u����MAXUALRMB7�P8 ��y���3�0]&q
��Ca]s�3�~��� 8@=@^+ �Z�v	��V0+�P1�A5d�r���U����� �E(iTy� ������/ / A/,/Q/w/b/�/~/�/ �/�/�/�/??)?O? :?s?V?�?�?�?�?�? �?�?O'OOKO.OoO ZOlO�O�O�O�O�O�O �O#__G_2_D_}_`_ �_�_�_�_�_�_�_o 
ooUo8oyodo�o�o �o�o�o�o�o�o-���D_LDXDIS�A^�� �MEMO�_APX�E ?��
 �0y� ���������ISC 1_�� �O����W�i� ����Ə�����}� �ߏD�/�h�z�a��� ����������� @���O�a�5������� �����u��ׯ<�'� `�r�Y������y�޿ �ۿ���8Ϲ�G�Y� -ϒ�}϶ϝ�����mπ����4��X�j�#�_MSTR `��~}�SCD 1as}�R���N�������� 8�#�5�n�Y��}�� �����������4�� X�C�|�g��������� ������	B-R xc������ �>)bM� q�����/� (//L/7/p/[/m/�/ �/�/�/�/�/?�/"? H?3?l?W?�?{?�?�?��?n�MKCFG �b���?��LT�ARM_�2cRu;B �3Wp|TNBpMETPUOp��2����NDS?P_CMNTnE@8F�E�� d���N��2A�O�D�EPO�SCF�G�NPS�TOL 1e-�4=@�<#�
;Q�1 ;UK_YW7_Y_[_m_�_ �_�_�_�_�_o�_o Qo3oEo�oio{o�o�a��ASING_CH�K  �MAqODAQ2CfO�7J�e�DEV 	Rz	�MC:'|HSI�ZEn@����eTA�SK %<z%$�12345678�9 ��u�gTRI�G 1g�� l<u%���3����>svvYPaq��kE�M_INF 1h�9G `�)AT&FV0�E0(���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ���ڄH�� ����G�ֈAO�w� 2�������џ ���� ����͏ߏP��t��� ����]�ί����� (�۟�^��#�5��� ��k�ܿ� ϻ�ů6� �Z�A�~ϐ�C���g� y��������2�i�C� h�ό�G߰��ߩ��� �ϫ��������d�v� )ߚ��߾�y����� ���<�N��r�%�7� I�[������9�& ��J[�g��>�ONITOR�@G� ?;{   	?EXEC1�3�U2�3�4�5�T�p�7�8�9�3�n�R�R�R RRR(R@4R@RLR2YU2e2q2}2�U2�2�2�2�U2�3Y3e3���aR_GRP_SOV 1it��q(�5�
��5��m۵MO~q_DC�d~�1PL_NAM�E !<u� ��!Defaul�t Person�ality (f�rom FD) ��4RR2k! 1j�)TEX)TH��!�AX d�?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO�O�O�Ox2-?�O�O �O__0_B_T_f_x_�b<�O�_�_�_�_�_ �_o o2oDoVoho&x�Rj" 1o�)&0=\�b, �9��b��a @D�  &�a?��c�a?�`�a�aA'�6�ew�;�	l�b	 ��xJ�p��`�`	p �< �(p�� �.r� K��K ��K=*��J���J���JV��kq`q�P��x�|� @j��@T;f�r�f��q�acrs�I5�� ��p���p�r��ph}�3��´7  ��>��p�h�`z��Ꝝ�"�Jm�q� H�N��ac��$�dw���  �  �P� Q� �� |  а�m�Əi}	'� � ��I� �  �����:�È~�È=���(��#�a	���I  ?�n @H�i~�ab�Ӌ�b�$w���"N0��  '�Ж�q�p@2��@Ǔ���r�q5�C��pC0C�@ C�����`
��A1]w@B�V~JX�
nwB0h�A���p�ӊ�p@����aDz���֏���Я	��pv�( �� -��I��-��=��A�a�we_q��`�p �?�ff� ��m��� ����Ƽ�!@ݿ:�>1�  P�apv(�`ţ� �=�qs�t��?���`x�`�� <
6b<�߈;܍�<��ê<� <�#&P�ό�AO��c�1��ƍ�?fff?�O�?&��qt@�.��J<?�`��wi4����dly�e ߾g;ߪ�t��p�[� ��߸ߣ����� ��0��6�wh�F0%� r�!��߷�1ى���~�E�� E�O�?G+� F�!��� /���?�e�P���t���lyBL�cB��Enw 4�������+��R�� s����������h�Ô�>��I�mXj���A�y�we�C�������A�#/*/c/N/wi������v/C�`� C!Hs/`
=$�p�<!�!���ܼ�'�3A��A�AR1AO��^?�$�?����±
=���>����3�?W
=�#�]�;�e��?������{����<����>(�B�u���=B0������	R���zH�F�G����G��H�U�`E���C�+���}I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0w/O*OONO9OrO ]O�O�O�O�O�O�O�O _�O8_#_\_G_�_�_ }_�_�_�_�_�_�_"o ooXoCo|ogo�o�o �o�o�o�o�o	B -fQ�u��� ����,��P�b� M���q�����Ώ��� ݏ�(��L�7�p�[� �����ʟ���ٟ� ��6�!�Z�E�W���#1�( ��9�K��y�ĥ �����<Ư!3�8���!4Mgs��,��IB+8�J��a���{�d�d���@��ȿ���ڼ%P8�	P�=:GϚ�S�06�h�z���R�Ϯ�`���������  %�� ��h�Vߌ�z߰� &�g�/9�$�������7����A�S�e�w�  ��������������2 F;�$�&Gb����a�����!C����@���8�����F�� DzN�� F�P D�������)#B�'9K�]o#?���@U@v
4$8�8���8�.
  v���!3E Wi{����:� ��ۨ�1���$MSKCF�MAP  ��?� ����(.�ONREL7  �!9���EXCFENB�E'
#7%^!FNC�e/W$JOGOVLKIME'dO S"d�WKEYE'�%�WRUN�,�%�SFSPDTY0xg&P%9#SIGNE/>W$T1MOT�/T!��_CE_GRoP 1p��#\x��?p��?�?�? �?�?O�?OBO�?fO O[O�OSO�O�O�O�O �O_,_�OP__I_�_ =_�_�_�_�_�_oo��_:o�TCOM_CFG 1q	-��vo�o�o
Va_/ARC_b"�p)UAP_CPL�o�t$NOCHECK� ?	+  �x�%7I[m ���������!�.+NO_WA�IT_L 7%S2NMT^ar	+�s�o_ERR_12s	)9�� ,ȍޏ���x���&��dT_�MO��t��, �S�*oq�9�PAR�AM��u	+���a�ß'g{�� =�?�345678901��,��K�]� 9�i�������ɯۯ��&g�����C��c�UM_RSPAC�E/�|����$ODRDSP�c#6p(�OFFSET_C�ART�o��DIS�ƿ��PEN_FI�LE尨!�ai��`O�PTION_IO��/��PWORK kve7s# �� V�ؤ��p�4�p��	 ���p��<����RG_DSBL'  ��P#������RIENTTO�D ?�C�� !=�#��UT_SIM_D$�"����V��LCT w�}�h�iĜa[�1�_P�EXE�j�RAT�vШ&p%� ��2^3j�)TEX)TH�>)�X d3��� ����%�7�I�[�m� ������������ �!�3�E���2��u� ��������������c�<d�ASew ���������Ǎ�^0OUa0o(��(����}u2, ����O H @D�  &[?�aG?��c�c�D][�Z�;��	ls���xJ���������<; ��� ��2��H(��H3k7�HSM5G�22�G���Gp
͜�'f�/-,2�KCR�>�D!�M#�{Z/��3�����4y H "�c/�u/�/0B_�����jc��t�!�/ �/�"t3�2����/6  U��P%�Q%��%��|T��S62�q?'e	�'� � �2�I� �  {��+==��ͳ?��;	�h	�0�I  �n @�2 �.��Ov;��ٟ?&&gN [OaA''�uDt@!� Cb@C�@F#�H!�/�O�O sb
S�Ab@�@�@���@�e`0Bb@QA8�0Yv: �13Uwz$oV_�/z_e_�_��_	��( �� -�2�1�1ta�Ua�c���:A-����.  �?�fAf���[o"o�_Uʈ`oXÜQ8���o�j>N�1  Po�V(�� �eF0�f�Y���L�/?����xb�P�<
6b<߈�;܍�<�ê�<� <�&�,/aA�;r�@Ov�0P?fff?�0?y&ip�T@�.{r�J<?�`�u #	�Bdqt�Yc�a �Mw�Bo��7�"� [�F��j�������ُ ����3�����,���(�E�� E���3G+� F� �a��ҟ�����,���P�;���B�pA Z�>��B��6�<OίD� ��P��t�=���a�s�x����6j�h��7o��>�S��O�`����Fϑ�A�a�_��C3Ϙ�/�%?��?���������
#	Ę��P �N||#CH���Ŀ����ރ�@I�_�'��3A�A�AR�1AO�^?�$��?��� �±�
=ç>�����3�W
=�#�� U��e���B���@��{�����<���(��B�u��=�B0�������	�b�H�F��G���G���H�U`E����C�+��I#��I��HD��F��E���RC�j=[�
�I��@H��!H�( E<YD0߻���� ����� �9�$�]�H� Z���~����������� ��#5 YD}h ������� 
C.gR��� ����	/�-// */c/N/�/r/�/�/�/ �/�/?�/)??M?8? q?\?�?�?�?�?�?�? �?O�?7O"O[OmOXO �O|O�O�O�O�O�O�O��O3_Q(�������b��gUU���W_i_2�3�8���_�_2�4Mgs8�_�_�RIB+�_�_��a���{� miGo5okoYo�o}lJ��P'rP�nܡݯ��o=_�o�_�[R?Q�u���  �p���o�� /��S��z
uүܠ�������ڱ������p�����  /��M�w�e��������l2� F�$��Gb	��t��a�`�p�S�C�y�@p�5�G�Y�~۠F� Dz���� F�P DC��]����پ���ʯܯ� ��~�?̯��@@�?�RK�K���K���
 �|������� Ŀֿ�����0�B�pT�fϽ�V� ���{���1��$PA�RAM_MENU� ?3���  DEFPULSEr��	WAITTM�OUT��RCV��� SHEL�L_WRK.$CUR_STYL��;	�OPT�ߧPTB4�.�C�R?_DECSN���e ��ߑߣ��������� ��!�3�\�W�i�{�����USE_PR_OG %��%��\���CCR���e�����_HOST !��!��:���AT�`�V��/�X�|����_TIME���^��  ��GD�EBUG\�˴�G�INP_FLMS�K����Tfp����P+GA  ����)�CH����TYPE
�������� ��� -?h cu������ �//@/;/M/_/�/ �/�/�/�/�/�/�/?�?%?7?`?��WOR�D ?	=	�RSfu	PNS2UԜ2JOK�DR�TEy�]TRA�CECTL 1xv3��� �`_l m&�`�`|�>�6DT Qy3��%@�0D � o `2@U,6D-6D.6D/6De06D16A�c2@ �`8BV�8BR�8BM 8BPJ�8BF�8B6D6DU	6D
6D6D6D6D6D6D^�8BU6D6D6D6DQ6D�8B6D6D~P8B6DV�8Bj�8B6D6DҀ8B�8B!6D"6D#6D�8BU%6D&6D'6D(6D)6D*6D5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐن.A �v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ��r����� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����������� �*��$P�GTRACELE�N  )�  ���(���>�_UP z����m�u�Y��n�>�_CFG �{m�W�(��n���PКӂ�DEFSPD |����aP��>�IN~��TRL }���(�8����PE__CONFI��~m՟�mњ�\�ղ�LID�����=�GRP 1���W��)�A ����&ff(�A�+33D�� D�]� CÀ A)@1��Ѭ(�d�Ԭ����0�0�� 	 �1�ح֚��� �������B�9�����O�9�s�(�>�?T?�
5��������� =��=#�
����P ;t_�����<��  Dz (�
H�X~i ������/��/D///h/S/�/���
V7.10be�ta1��  �A�E�"ӻ�A (�� ?!G���!>���"�܇��!���!BQ��!A\� �!��T�!2p����Ț/ 8?J?\?n?};� ����/��/�?}/�?�? OO:O%O7OpO[O�O O�O�O�O�O�O_�O 6_!_Z_E_~_i_�_�_ �_�_�_�_'o2o�_ VoAoSo�owo�o�o�o �o�o�o.R=�v1�/�#F@  �y�}��{m��y=� �1�'�O�a��?�?�? ������ߏʏ��'� �K�6�H���l����� ɟ���؟�#��G� 2�k�V���z������� �o��ίC�.�g� R�d����������п 	���-�?�*�cώ� ��Ϯ������ B�;�f�x�������D� ���߶��������7� "�[�F�X��|��� ��������!�3��W� B�{�f��������� � ����/S>w bt������ =OzόϾψ ����ϼ� /.�'/ R�d�v߈߁/0�/�/ �/�/�/�/�/#??G? 2?k?V?h?�?�?�?�? �?�?O�?1OCO.OgO RO�OvO�O�O���O�O �O__?_*_c_N_�_ r_�_�_�_�_�_o�_ )oTfx�to�� �/�o/>/P/ b/t/mo�|�� �����3��W� B�{�f�x�����Տ�� �����A�S�>�w� b����O��џ����� �+��O�:�s�^��� ����ͯ���ܯ�@o Rodo�o`��o�o�o�� ƿ�o���*<N� Y��}�hϡό��ϰ� �������
�C�.�g� Rߋ�v߈��߬����� 	���-��Q�c�N�� �����l������� �;�&�_�J���n��� ��������,�>�P� :L��������� ���(�:�3��0 iT�x���� �/�///S/>/w/ b/�/�/�/�/�/�/�/ ??=?(?a?s?��? �?X?�?�?�?�?O'O OKO6OoOZO�O~O�O �O�O�O*\&_8_�r���_�_��$�PLID_KNO�W_M  ��� Q�TSoV ���P��?o"o 4o�OXoCoUo�o R��SM_GRP 1���Z'0{`�@R�`uf�e�`
�5 � �gpk' Pe]o�����������SMR��c��mT�EyQ}? yR����������� ����ӏ�G�!��-� ����������韫��� ϟ�C���)������������寧���QS�T�a1 1���)���P0� A 4��E2�D�V�h��� ����߿¿Կ���9� �.�o�R�d�vψ���P�Ͼ����2�0�N Q�<3��3�/�A�S��4l�~ߐ����5���������A6
��.�@��7Y�k�}���8���������MAD  �)��PAR�NUM  !��}o+��SCHE� �S�
��f���S��UPDf�x��_CMP_�`H�� ��'�UER_wCHK-���ZE*<RSr��_�QG_MOG���_�~X�_RES_G��!���D�>1 bU�y������/�	/��� �+/�k�H/g/l/� �Ї/�/�/�	��/�/ �/�X�?$?)?��� D?c?h?����?�?�?�V 1��U�ax�@c]�@t@(�@c\�@�@D�@c[�*@��T?HR_INRr�J���b�Ud2FMASS6?O ZSGMN>OqC�MON_QUEUE ��U�V P~P� X�N$ UhN8�FV�@END�A���IEXE�O�E��B�E�@�O�COPTI�O�G��@PROG�RAM %�J%��@�?���BTAS�K_IG�6^OCFG ��Oz��_�P�DATA�c��[@Ц2=�DoVoho zo�j2o�o�o�o�o�o�);M jIN+FO[��m��D �������� 1�C�U�g�y����������ӏ���	�dwpt��l )�QE DI�T ��_i��^W�ERFLX	C�RGADJ �tZA�����?נʕFA~��IORITY�G�W���MPDSP(NQ����U�GD��oOTOE@1�X� (!AF:@�E� c�Ч!t�cpn���!u�d����!icm����?<�XY_�Q�X���Q)� a*�1�5��P�� ]�@�L���p������� �ʿ��+�=�$�a��Hυϗ�*��POR�T)QH��P�E���_CARTRE�PPX��SKSTyA�H�
SSAV�@��tZ	2500H863���_x�
Ԫ'��X�@�s�wPtS�ߕߧ���UR�GE�@B��x	WFF��DO�F"[W\��������WRUP_�DELAY �|X���R_HOTqX�	B%�c���R_NORMALq^R��v�SEMI�����9�QSKIP'��vtUr�x 	7� 1�1��X�j�|�?�tU �������������� $J\n4�� ������4 FX|j��� ����/0/B//�R/x/f/�/�/�/tU�?$RCVTM$��D��� DCR'����Ў!C`N��C�d�C��o�?��>��L�<|�{:��g��&��/����%�t����|��}'�:�o?��� <
6b<�߈;܍�>u�.�?!<�&�?h?�?�?�@>� �?O O2ODOVOhOzO �O�O�O�O�O�?�O�O __@_+_=_v_Y_�_ �_�?�_�_�_oo*o <oNo`oro�o�o�o�_ �o�o�o�o�o8J -n��_���� ���"�4�F�X�j� U������ď���ӏ ���B�T��x��� ������ҟ����� ,�>�)�b�M������� �����ïկ�Y�:� L�^�p���������ʿ ܿ� ����6�!�Z� E�~ϐ�{ϴϗ����� -�� �2�D�V�h�z� �ߞ߰���������
� ��.��R�=�v��k� ����������*� <�N�`�r��������� ��������&J \?������ ��"4FXj�|��!GN_AT�C 1�	; �AT&FV0�E0�ATD�P/6/9/2/�9�ATA��,AT%G1�%B960�W+++�,�H/�,�!IO_TYPOE  �%�#t��REFPOS1� 1�V+ x	�u/�n�/j�/ 
=�/�/�/Q?<?u??��?4?�?X?�?�?�+2 1�V+�/�?�?�\O�?�O�?�!3 1�O*O<OvO�O�O_>�OS4 1��O�O��O_�_t_�_+_S5 1�B_T_f_�_o�	oBo�_S6 1� �_�_�_5o�o�o�oUoS7 1�lo~o�o��oH3l�oS8 1�%_����SMASK ;1�V/  
?�M�N�XNOS/�r�������!MOTE � n��$��_CFG� ����q���"P?L_RANG������POWER 壧���SM_�DRYPRG �%o�%�P��TA�RT ��^�U?ME_PRO-�?�����$_EXEC_?ENB  ���GSPD��Րݘ���TDB��
�RM\�
�MT_'�T�����OBOT_NAME o�����OB_OR�D_NUM ?��b!H863  �կ����PC_T�IMEOUT�� �x�S232Ă1��� LT�EACH PEN�DAN��w���-��Main�tenance �Cons���s�"����KCL/C�m��

���t�ҿ �No Use�-��Ϝ�0�NPO��򁋁���.�CH_L���̫��q	��s�MA�VAIL�����������SPACE1w 2��, j�@߂�D��s�߂� ��{S�8�?� k�v�k�Z߬��ߤ��� �� �2�D���hߊ� |��`������� ��� �2�D��h�� |���`���������y�
��2����0�B� ��f�����{���3);M _������/� /44FX j|*/���/�/�/ ?(??=?5Q/c/ u/�/�/G?�/�/�?O@�?$OEO,OZO6n? �?�?�?�?dO�?�?_�,_�OA_b_I_w_7 �O�O�O�O�O�_�O_ (oIoo^oofo�o8�_�_�_�_�_�oo 6oEf){����G �o�� ���
M�  ���*�<�N�`�r��� ����w���o�収���d.��%�S�e� w�����������Ǐَ ���Θ8�+�=�k�}� ������ůׯ͟��� �%�'�X�K�]����� ����ӿ�������#�E�W� `� @�������x�����\�e�������� ���R�d߂�8�j߬� �߈ߒߤ�������� ��0�r���X���� ��������8�����
�ύ�_MOD�E  �{��S ���{|�2�0� ����3�	S|�)CWORK_A�D��=9(+R  �{�`� ��� _INTVAL����d���R_OPoTION� ���H VAT_GR�P 2��u�p(N� k|��_��� ��/0/B/��h�u/ T� }/�/�/�/�/�/ �/?!?�/E?W?i?{? �?�?5?�?�?�?�?�? O/OAOOeOwO�O�O �O�OUO�O�O__�O =_O_a_s_5_�_�_�_ �_�_�_�_o'o9o�_ Iooo�o�oUo�o�o�o �o�o�o5GYk -���u��� ��1�C��g�y��� M�����ӏ叧�	�� -�?�Q�c��������� ������ǟ�;��M�_����$SCAN_TIM��_%�}�R �(ӿ#((�<04�d d 
!D�ʣ��u�a/�����U�E�25�����dA�D8�H�g��]	����������dd�x� � P���� ��  8� ҿ�<!���D��$�M� _�qσϕϧϹ���������ƿv���F�X��/� ;��ob��pm��t�_DiQ|̡  � l� |�̡ĥ�������!� 3�E�W�i�{���� ����������/�A� S�e�]�Ӈ������� ������);M _q������ �r���j�Tf x������� //,/>/P/b/t/�/��/�/�/�/�%�/  0��6��!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O*�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo�O�OJ�o�o�o �o�o�o�o 2D Vhz�����`��
�7?  ;� >�P�b�t��������� Ǐُ����!�3�E��W�i�{�������ß �ş3�ܟ��&� 8�J�\�n�������������ɯ�����,� �+�	�12345678^�� 	� =5���f�x�������������
��.�@� R�d�vψϚ�៾��� ������*�<�N�`� r߄߳Ϩߺ������� ��&�8�J�\�n�� ������������� "�4�F�u�j�|����� ����������0 _�Tfx���� ���I>P bt������ �!/(/:/L/^/p/��/�/�/�/�/�/� 2�/?�#/9?K?]?��iCz  Bp�˚   ��h2���*�$SCR_�GRP 1�(��U8(�\x�d�@ >� �'��	  �3�1�2�4(1*�&�I�3�F1OOXO}m��D�@�0ʛ)����HUK�LM-�10iA 890�?�90;��F;�M61C D�:�CP�*�1
\&V�1	��6F��CW�9)A7Y	�(R�_�_�_�_�_�\���0i^�oO UO>oPo#G�/���o�'o�o�o�o�oB�B0�rtAA�0*  @�Bu&Xw?��ju�bH0{Uz�AF@ F�` �r��o����� +��O�:�s��mBqrr`����������B�͏ b����7�"�[�F�X� ��|�����ٟğ���N����AO�0�B�CU
�L���E�jqBq>HE����$G@�@pϯ B���G�I
E��0EL_DEFA�ULT  �T�_�E���MIPOWERFL  
E*��7�oWFDO� *���1ERVENT �1���`(��� L!DUM_�EIP��>��j!AF_INE�<¿C�!FT�������!o:� ���a�!RPC�_MAINb�DȺ8Pϭ�t�VIS}�C�y�����!TP���PU�ϫ�d��E�!�
PMON_PR'OXYF߮�e4ߑ���_ߧ�f����!RDM_SRV��r��g��)�!R�dIﰴh�u�!
v��M�ߨ�id���!?RLSYNC��>��8���!ROS��4��4��Y�(� }���J�\��������� ����7��["4 F�j|�����!�Eio�ICE_KL ?%�� (%SVCPRG1n>���3D��3���4/D/�5./3/�6V/[/�7~/�/��D�/�9�/�+�@��/ ��#?��K?�� s?� /�?�H/�?� p/�?��/O��/;O ��/cO�?�O�9? �O�a?�O��?_� �?+_��?S_�O{_ �)O�_�QO�_�yO �_��Os���� >o�o}1�o�o�o�o�o �o�o;M8q \������� ��7�"�[�F��j� ������ُď���!� �E�0�W�{�f����� ß���ҟ���A� ,�e�P���t���������ί�y_DEV� ��M{C:�@`!�OUT��2��?REC 1�`e��j� �� 	 �����˿���ڿ��
 �`e��� 6�N�<�r�`ϖτϦ� �Ϯ�������&��J� 8�n߀�bߤߒ��߶� ������"��2�X�F� |�j���������� ����.�T�B�x�Z� l������������� ,P>`bt� �����( L:\�d��� �� /�$/6//Z/ H/~/l/�/�/�/�/.� �/?�/2? ?V?D?f? �?n?�?�?�?�?�?
O �?.O@O"OdORO�OvO �O�O�O�O�O�O__ <_*_`_N_�_�_x_�_ �_�_�_�_oo8oo ,ono\o�o�o�o�o�o �o�o�o "4j X������� ���B�$�f�T�v� �����������؏� �>�,�b�P�r���p�oV 1�}� P
��l!����� ����TYPE�\��HELL_C�FG �.���� ��r�����RSR������ӯ�� �����?�*�<�u� `�����������ο�  �%@�3�E��Q�\�Ӑ1M�o�p��d���2Ӑd]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&��1�OW_REG�_UI���IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he�#�� ��������Ӕ��) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������o���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( ��}/xcopy �fr:\*.* �virt:\tm�pback7=>�inspiron:12732 Ypbt�� }0.a6HZ_���
xyzrate 61 ����n���.M4804 HZ���/�3/s:or�derfil.dat<�a/s/�/�/z� */mdb:9@�Y/�/�/?�	.. A��/n?�?�?�- �G?�^?�?OO&/ 8/�/�/mOO�O�/�/ �/ZO�O�O_"?4?�? X?i_{_�_�?�?C_�? �_�_oO0OBOTOeo wo�o�O�OIo�O�o�o ,_�_P_as� ��_;�_`��� (���o������M
28�Y����� !o3o�o��a�s����� �oE���Y�����! 3F�ݟn������ 6�H�ŀ^����&� 8���ܟm�������� ȟZ�����"�4�ǯ X�i�{ύϠ���C�֯ ������0�����e�`w߉ߜ����06� X������ �2Թ������n���߷2076G�Y������!� 3�����a�s������� E���Y�����!�3� F�����n����6 H��^�&�8� ����m������� Z��/"4�X i/{/�/��C/��/ �/?0BTe?w? �?��I?��?�?O�O�$SNPX_�ASG 1�����9A�� P 0 '�%R[1]@1�.1O 9?�$3% dO�OsO�O�O�O�O�O �O __D_'_9_z_]_ �_�_�_�_�_�_
o�_ o@o#odoGoYo�o}o �o�o�o�o�o�o* 4`C�gy�� �����	�J�-� T���c�������ڏ�� ���4��)�j�M� t�����ğ������ݟ �0��T�7�I���m� �������ǯٯ��� $�P�3�t�W�i����� ���ÿ����:�� D�p�Sϔ�wω��ϭ� �� ���$���Z�=� dߐ�sߴߗߩ����� �� ��D�'�9�z�]� ���������
��� �@�#�d�G�Y���}� ������������* 4`C�gy�� ����	J- T�c����� �/�4//)/j/M/ t/�/�/�/�/�/�/�/�?0?4,DPARAoM �9ECA_ �	��:P�4��0$HOFT_�KB_CFG  �q3?E�4PIN_�SIM  9K��6�?�?�?�0,@RV�QSTP_DSBº>�21On8J0SR� ��;� & �MULTIROBOTTASK=O�q3�6TOP_�ON_ERR  ��F�8�APTN ��5�@�A�BRING_P�RM�O J0VD�T_GRP 1�<Y9�@  	�7n8 _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D khz����� ��
�1�.�@�R�d� v���������Џ��� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\��������� ��ȯگ����"�I� F�X�j�|�������Ŀ ֿ����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�a�^�p��� ��������� �'�$� 6�H�Z�l�~���������������3VPRG�_COUNT�6q��A�5ENB�O�M=�4J_UP�D 1��;8  
q2���� �� )$6Hq l~�����/ �/ /I/D/V/h/�/ �/�/�/�/�/�/�/!? ?.?@?i?d?v?�?�? �?�?�?�?�?OOAO <ONO`O�O�O�O�O�O �O�O�O__&_8_a_�\_n_�_�_�_YS�DEBUG" � ��Pdk	�PSP_PwASS"B?�[�LOG ���m�P�X�_ � �g�Q
MC�:\d�_b_MPACm��o�o�Qa��o �vfSAV ��m:dUb�U�\gSV�\TEM�_TIME 1��� (�`�Q�a��2o	T1SVGU�NS} #'k��spASK_OPT�ION" �go�spBCCFG ��| �b�{�}`����a&�� #�\�G���k�����ȏ ������"��F�1� j�U���y���ğ��� ӟ���0��T�f��UR���S���ƯA��� ��� ��D��nd��t 9�l���������ڿȿ �����"�X�F�|� jϠώ��ϲ������� ��B�0�f�T�v�x� ���ߦؑ������� (��L�:�\��p�� ���������� �6� $�F�H�Z���~����� ��������2 V Dzh����� ����4Fdv ������/ /*/�N/</r/`/�/ �/�/�/�/�/�/?? 8?&?\?J?l?�?�?�? �?�?�?�?�?OO"O XOFO|O2�O�O�O�O �OfO_�O_B_0_f_ x_�_X_�_�_�_�_�_ �_oooPo>otobo �o�o�o�o�o�o�o :(^Lnp� ����O��$�6� H��l�Z�|�����Ə ؏ꏸ����2� �V� D�f�h�z�����ԟ ����
�,�R�@�v� d���������ίЯ� ��<��T�f����� ��&�̿��ܿ��&� 8�J��n�\ϒπ϶� �����������4�"� X�F�|�jߌ߲ߠ��� ��������.�0�B� x�f��R��������� ���,��<�b�P��� ����x��������� &(:p^�� ����� 6 $ZH~l��� �����/&/D/V/ h/��/z/�/�/�/�/��&0�$TBCS�G_GRP 2���%� � �1 
 ?�  /?A?+?e?O? �?s?�?�?�?�?�;2�3�<d, ��$A?1	 HC{���6>��@E~�5CL  B�'2�^OjH4J��B�\)LFY  A��jO�MB��?�IBl��O�O�@�JG_�@�  D	�15_ __�$YC-P{_F_`_j\��_�]@0�>�X�Uo �_�_6oSoo0o~o�o��k�h�0	V�3.00'2	mw61c�c	*�`0�d2�o�e>�JC0(�a�i ,p�m-w  �0����o�mvu1JCFG [��% 1 #0Vvz��rBrv�x����z�  �%��I�4�m�X��� |��������֏��� 3��W�B�g���x��� ��՟�������� S�>�w�b�����'2A  ��ʯܯ������E� 0�i�T���x���ÿտ 翢����/��?�e� 1�/���/�ϜϮ��� �����,��P�>�`� ��tߪߘ��߼����� ���L�:�p�^�� ����������� � 6�H�>/`�r������ ���������� 0 Vhz8���� ��
.�R@ vd������ �//</*/L/r/`/ �/�/�/�/�/�/�/�/ ?8?&?\?J?�?n?�? �?�?�?���?OO�? FO4OVOXOjO�O�O�O �O�O�O__�OB_0_ f_T_v_�_�_�_z_�_ �_�_oo>o,oboPo roto�o�o�o�o�o �o(8^L�p �������$� �H�6�l�~�(O���� f�d��؏���2� � B�D�V�������n��� �ԟ
���.�@�R�d� ���v��������Я ���*��N�<�^�`� r�����̿���޿� �$�J�8�n�\ϒπ� �Ϥ�������ߊ�(� :�L���|�jߌ߲ߠ� ���������0�B�T� �x�f�������� �����,��P�>�t� b��������������� :(JL^� ����� � 6$ZH~l�� ^���dߚ //D/ 2/h/V/x/�/�/�/�/ �/�/�/?
?@?.?d? v?�?�?T?�?�?�?�? �?OO<O*O`ONO�O rO�O�O�O�O�O_�O &__6_8_J_�_n_�_ �_�_�_�_�_�_"oo Fo��po�o,oZo�o �o�o�o�o0T fx�H���� ���,�>��b�P� ��t���������Ώ� �(��L�:�p�^��� ����ʟ���ܟ� � "�$�6�l�Z���~��� ��دꯔo��&�Я V�D�z�h�������Կ ¿��
��.��R�@�pv�dϚτ�  ����� ��������$TBJOP_G�RP 2ǌ���  ?i������������x�JBЌ��9� �_< �X����� @���	 ߐC�� t�b � C����>�c�͘Րդ�>̚���ѳ33=�{CLj�fff?��?�ffBG��ь������t�ц�>�(�\)�ߖ�E�����;��hC=Yj��  @h��?B�  A�����f��C�  Dphъ�1��O�4��N����
:���Bl^��j�i�l��l����Aə�A��"��D��֊�=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������$�6�>B�\��T����Q�tsx�@333@���C���y��1����>��D�h����������<'{�h�@i�  ��t��	�� �K&�j�n |���p�/�P/:/k/�ԇ���!���	V3.00�J�m61cI��*� IԿ��/�' �Eo�E���E��E��F��F!��F8��FT��Fqe\F�N�aF���F�^�lF���F�:�
F�)F���3G�G���G��G,I��!CH`�C��dTDU�?D���D��DE(�!/E\�E���E�h�E��ME��sF�`F+'\FD���F`=F}�'�F��F��[
F���F���M;��;Q�*T,8�4` *�ϴ?
�2���3\�X/O���ESTPARS�  ��	���HR�@ABLE 1ʒ���0��
H�7 (8��9
G
H
H��T��
G	
H

H
HTYE��
H
H
H�6FRDIAO��XOjO|O�O�O�ETO "_4[>_P_b_t_�^:B	S _� �JGoYoko }o�o�o�o�o�o�o�o 1CUgy� ���`#oRL�y�_�_ �_�_�O�O�O�O�OX�:B�rNUM  V���P���� V@P:B_CFGG ˭�Z�h�@���IMEBF_TT�%AU��2@�VER�S�q��R 1=���
 (�/��	��b� ����J�\� ��j�|���ǟ��ȟ֟ �����0�B�T��� x�������2�_����@�
��MI_CWHAN�� � ���DBGLV����������ETHER_AD ?��O�������h�����oROUT�!���!������SNM�ASKD��U�255.���#������OOLOFS_D�I%@�u.�ORQCTRL ��� ��}ϛ3rϧϹ����� ����%�7�I�[�:����h�z߯�APE_�DETAI"�G�P�ON_SVOFF�=���P_MON ��֍�2��ST�RTCHK ��^�����VTCOMPAT��O������FPROG %�^�%MULTI?ROBOTTݱ��<��9�PLAY&H��_INST_Mްe ������US��q��LCK���Q?UICKME�=�ރ�SCREZ�>G�tps� �� �u�z����_��@@�n�.�SR_GRP� 1�^� �O����
��+ O=sa�쀚 �
m������L/ C1gU�y �����	/�-/�/Q/?/a/�/	1?234567�0�/��/@Xt�1���
� �}ipnl�/� gen.htm�? ?2?D?V?`�Panel _setupZ<}P���?�?�?�?�?�?  �??,O>OPObOtO�O �?�O!O�O�O�O__ (_�O�O^_p_�_�_�_ �_/_]_S_ oo$o6o HoZo�_~o�_�o�o�o �o�o�oso�o2DV hz�1'�� �
��.��R��v����������ЏG���U�ALRM��G ?9� �1�#�5� f�Y���}�������џ�ן���,��P��S�EV  �����ECFG ���롽�A�� �  BȽ�
  Q���^����	��-� ?�Q�c�u������������� ������I��?���(% D�6� �$�]�Hρ�l� �ϐ��ϴ�������#�0�G���� �߿�U�I_Y�HIST� 1��  �(�� ��3/�SOFTPART�/GENLINK�?current�=editpage,��,1���!�3��� ����mwenu��962�߀�����K�]�o�36u�
��.�@���W� i�{���������R��� ��/A��ew ����N�� +=O�s��������f��f //'/9/K/]/`�/ �/�/�/�/�/j/�/? #?5?G?Y?�/�/�?�? �?�?�?�?x?OO1O COUOgO�?�O�O�O�O �O�OtO�O_-_?_Q_ c_u__�_�_�_�_�_ �_��)o;oMo_oqo �o�_�o�o�o�o�o �o%7I[m�  ������� 3�E�W�i�{������ ÏՏ�������A� S�e�w�����*���џ �����ooO�a� s���������ͯ߯� ��'���K�]�o��� ������F�ۿ���� #�5�ĿY�k�}Ϗϡ� ��B���������1� C���g�yߋߝ߯��� P�����	��-�?�*� <�u��������� ����)�;�M����� ������������l� %7I[��� ����hz! 3EWi���� ���v////A/�S/e/P���$UI�_PANEDAT�A 1������!  	�}w/�/�/�/�/?? )?>?��/ i?{?�?�?�?�?*?�? �?OOOAO(OeOLO �O�O�O�O�O�O�O�O\_&Y� b�>R Q?V_h_z_�_�_�__ �_G?�_
oo.o@oRo do�_�ooo�o�o�o�o �o�o*<#`G ��}�-\�v�# �_��!�3�E�W�� {��_����ÏՏ��� `��/��S�:�w��� p�����џ������ +��O�a������� ��ͯ߯�D����9� K�]�o��������ɿ ���Կ�#�
�G�.� k�}�dϡψ����Ͼ� ��n���1�C�U�g�y� ���ϯ���4�����	� �-�?��c�J��� ������������� ;�M�4�q�X����� ������%7�� [������� @��3Wi P�t����� /�//A/����w/�/ �/�/�/�/$/�/h? +?=?O?a?s?�?�/�? �?�?�?�?O�?'OO KO]ODO�OhO�O�O�O �ON/`/_#_5_G_Y_ k_�O�_�_?�_�_�_ �_oo�_Co*ogoyo `o�o�o�o�o�o�o�o -Q8u�O�O}��������)�>��U-�j�|� ������ď+��Ϗ� ��B�)�f�M����� ���������ݟ�&��S�K�$UI_P�ANELINK �1�U � �  ���}1234567890s������� ��ͯդ�Rq����!� 3�E�W��{�������ÿտm�m�&����Qo�  �0�B�T� f�x��v�&ϲ����� ����ߤ�0�B�T�f� xߊ�"ߘ��������� �߲�>�P�b�t�� ��0���������� ��$�L�^�p�����,� >������� $�0,&�[gI�m ������� >P3t�i�� Ϻ� -n��'/9/ K/]/o/�/t�/�/�/ �/�/�/?�/)?;?M? _?q?�?�UQ�=�2 "��?�?�?OO%O7O ��OOaOsO�O�O�O�O JO�O�O__'_9_�O ]_o_�_�_�_�_F_�_ �_�_o#o5oGo�_ko }o�o�o�o�oTo�o�o 1C�ogy� ����B�	�� -��Q�c�F�����|� ������֏�)�� M���=�?��?/ȟ ڟ����"�?F�X� j�|�����/�į֯� ����0��?�?�?x� ��������ҿY��� �,�>�P�b��Ϙ� �ϼ�����o���(� :�L�^��ςߔߦ߸� ������}��$�6�H� Z�l��ߐ������� ��y�� �2�D�V�h� z����-��������� 
��.RdG� �}����c� ��<��`r��� �����//&/8/ J/�n/�/�/�/�/�/ 7�I�[�	�"?4?F?X? j?|?��?�?�?�?�? �?�?O0OBOTOfOxO �OO�O�O�O�O�O_ �O,_>_P_b_t_�__ �_�_�_�_�_oo�_ :oLo^opo�o�o#o�o �o�o�o ��6H �l~a���� ����2��V�h� K�������1�U 
��.�@�R�d�W/�� ������П������ *�<�N�`�r��/�/? ��̯ޯ���&��� J�\�n�������3�ȿ ڿ����"ϱ�F�X� j�|ώϠϲ�A����� ����0߿�T�f�x� �ߜ߮�=�������� �,�>���b�t��� ���+������ :�L�/�p���e����� ������ ��6��🯡�ۏ��$UI�_QUICKME�N  ����}��RESTORE 1٩��  ��
�8m 3\n���G� ���/�4/F/X/ j/|/'�/�/�//�/ �/??0?�/T?f?x? �?�?�?Q?�?�?�?O O�/'O9OKO�?�O�O �O�O�OqO�O__(_ :_�O^_p_�_�_�_QO [_�_�_I_�_$o6oHo Zoloo�o�o�o�o�o {o�o 2D�_Q cu�o����� ��.�@�R�d�v���������Џ⏜SC�RE� ?��u1sc� uU2�3�4�5��6�7�8��UGSER����T����ks'���4��5*��6��7��8��� �NDO_CFG �ڱ  �  �� PDATE �h��Non�e�SEUFRA_ME  ϖ���RTOL_AB�RT����ENB�(��GRP 1���	�Cz  A�~�|�%|��������į֦��X�� U�H�X�7�MSK  �K�S�7�N�%�uT�%�����VI�SCAND_MA�XI�I�3���FAIL_IMGI��z �% #S���IM�REGNUMI�
����SIZI�� ��ϔ,�ONT�MOU'�K�Ε��&����a���a��s�F�R:\�� � �MC:\(�\wLOGh�B@Ԕ !{��Ϡ������z MCV�����UD1 �E�X	�z ��PO�64_�Q���n6��PO!�LI��Oڞ�e�V�N��f@`�I�� =	�_�SZVmޘ���`�WAImߠ�ST�AT �k�% @��4�F�T�$#�x� �2DWP  ���P G��=���͎���_�JMPERR 1�ޱ
  �p23�45678901 ���	�:�-�?�]� c���������������x��$�MLOW��8������_TI/�˘�'��MPHASOE  k�ԓ� ���SHIFT%�15 Ǚ��<z� �_����F /|Se��� ����0///?/ x/O/a/�/�/�/�/�/�����k�	VSwFT1\�	V���M+3 �5�Ք �p����A�  BU8[0[0�Πpg3�a1Y2�_3Y�7ME���K�͗	6e���&+%��M���b���	��$��TDI�NEND3�4��4O H�+�G1�OS2OI�V I���]LRELEvI��4.�@��1?_ACTIV�IT�<�B��A �m��/_��BRDBГOZ�YBOX �ǝ�f_\��b�2�T�I190.0m.�P83p\�V�254p^�Ԓ	� �S�_�[b��robot84�q_   px�9o\�pc�P ZoMh�]Hm�_Jk@1�o^�ZABCd��k�,���P\�Xo}�o0 );M�q�� ������>��a	Z�b��_V