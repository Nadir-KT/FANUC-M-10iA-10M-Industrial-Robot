��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ����ALRM_�RECOV1   $ALMO�ENB��]ON�i�APCOUPwLED1 $[�PP_PROCE�S0  �1�(|URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y12 � u3�|4|GRG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WAx�471�:OFF_ �N�3DELHLO�Gn25Aa2?i1@N?�� -M��H W+0�$Y �$DB� 6COMW!2MO� 21\D�.	 \rVE��1$F��A{�$O��D�B�CTM�P1_F�E2�G1�_�3�B�2�"XD��#
 d $�CARD_EXI�ST4$FSS�B_TYPuAH�KBD_S�B�1A�GN Gn $�SLOT_NUM�JQPREV,DB�U� g1G ;1_ED�IT1 � *1G=� S�0�%$EP�$�OP�AEToE_OKRUS�oP_CRQ$;4x�V� 0LACIw�1�RAPk �1x@M}E@$D�V��Q�Pv�A{oQLv� OUzR ,mAЧ0�!� B� LM�_O�^eR�"CAsM_;1 xr~$ATTR4�NP� ANN�@5I�MG_HEIGH|Q�cWIDTH4�VT� �UU0F_�ASPECQ$�M�0EXP��@A�X�f�CFT ?X $GR� � �S�!�@B@NFL�I�`t� UIREx 3dTuGITCHCj�`N� S�d_L�`2�C�"�`EDlpE
� J�4S�0� �zsa�!ip;G0 �� 
$WARNM��0f�!,P� �s�pN{ST� CORN�"�a1FLTR�uTRkAT� T�p H0ACCa1���{��ORI
`"S={R�T0_S�B�qHG�,I1 [ Thp�"3I9�TY�D(,P*2 �`w@� X�!R*HD�cJ* TC��2��3��4��U5��6��7��8���94�qO�$ <� $6xK3 1w`�O_M�@�C t� � E#6NGP�ABA� �c��ZQ ���`���@nr���� ��P�0����x�p�PzPb26��4��"J�_R��B�C�J��3�JV P��tBS��}Aw��"v�tP_*0OFSzRw @� RO_K8̨��aIT�3��NO�M_�0�1ĥ38���T �� $�d��AxP��K}EX��� �0g0I01��p�
�$TFa��C$MDM3��TO�3�0U� ^�� �Hw2J�C1|�EΡg0wE�{vF�vF�40CPhp@�a2 
P$A`�PU�3N)#�dR*�AX�!sDEwTAI�3BUFV8��p@1 |�p۶��pPIdT� PP�[�MZ�Mg�Ͱj�F>[�SIMQSI�"0��A.���� ��lw' Tp|zM��P��B�FACTrbHPEW7�P1Ӡ��vv��MCd� ��$*1JB�p<�*1D#ECHښ�H���b�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF4��� &k�Bv�u�cu��a E�� !2��+�MQ��EчSIZ�3����T��P�����aRSINF�����kq��������LX������F�CRCMu�3CC lpG��p���O}���b��1�������2�V�D
xIC��C���r����0P��{� EV �zUF_��F�pNB
0�?������A�! �r�Rx���� V�lp�2��aR�t�,��g�RTx �#�5�5"2��uARt���`CX�$LG�p��B�1 `s�P�t�a!A�0{�У+0R���tME�`!BupCr3RA 3tAZ�л4�pc�OT�FC�b�`��`FNp���1��ADI+�a%��b��{��p$�pSp�c�`S0�P��a,QMP6�`IY�3��M'�pU���aU  $m@TITO1�S�S�!���$�"0�DBPXW�O��!��$S�K��2�P� �"��"@�PR8� 
p� ���# m@6q1$��$��+ЅL9$?(�V�%�@?R4C&_?R4E3NE��'~?(��� RE�pY2(H� �OS��#$L�3$$3R��;43�MVOk_D@!V�ROScrr�w�S���~CRIGGER2F�PA�S��7�ETUsRN0B�cMR_���TUː[��0EW5M%���GN>`��FRLA���Eݡ�P��&$P�t�'��@4a��C�DϣV�D�XQ��4�1��MVGO�_AWAYRMO�#�aw!�DC{S_)  `IS#� �� �s3S�AQ汯 4Rx�ZS W�AQ�p�@1UW��cT'NTV)�5RV
a�@��|c�éWƃ��JBx��x0��SAFEۥ��V_SV�bEXC�LUU�;��ON�L��cYg�~az�OyT�a{�HI_V? ���R, M�_ *Ȥ0� ��_z�2� �p�QSGO  +�rƐm@�A�c~b����w@��V�i�b�fA�NNUNx0�$�dI%DY�UABc�@Sp �i�a+ �j�f�!�p�OGIx2,��$1F�b�$ѐOT�@A� $DUMMAY��Ft��Ft±� |6U- ` !�HE�|s��~bc�B�@ SUFFI���4PCA�Gs5�Cw6CrZ� MSW�U. 8!�KEYI��5�TM�1�s�qoA�vINޱE��!, �/ D��HOST�P!4���<���`<�°<��p<�EM'����Z�� SBL� U}L��0  �	8����DT�0?1 � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0�QS�����#��SAV �����c�S< 9�`��fP$�0E!� YwN_B�#2 0�`DI�d�pO|�m��#�$F�R_IC�� �ENC2_Sd3  ��< 3�9���� cgp����B4�"��2�A��ޖ5���`ǻ��@Q@K&D-!�a�A�VER�q����D3SP
���PC_�q���"�|�ܣ�VALMU3�HE�(�M�sIP)���OPPm �TH�*���S" T�/�Fb�;�d����d D����1�6 H(rLL_DUǀ�a�@��k���֠OT�"U�/���@@NOAUT5O70�$}�x�~�@s��|�C� ���C� 2iaz�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|�pw�����9 <���z�ΓKI����H猡�BaFEq@{@:� ,��&a? �P_P?��>�����E�@��	r�RP��z;fp$TP�?$VARI����n,�UP2Q`< W�߃TD��g���`��p����ia��BAC�"G= T2����$)�,p+r³�p IFI�� �p�� q M�P"$��Fl@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� FW�@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(��a�#5T�DG���� �%��FSS� )�?C P(q1�1�`Q_1"811�EC�13D;5D6�GR)A���@�����P�W�ON2EBUG�S�2�C`gϐ_E A ���?�WA�TERM�5B�5���ORI�w�0C�5X��SM�_-`���0D�52��TA�9EIU}P��F� -Q�ϒA�P�3�@B$gSEGGJ� EL�UwUSEPNFI��pBx��1@��4>DC�$UF�P��$���Q�@C���G�0qT�����SNSTj��PATۡg��APTHJq�A�E*�Z%qB�\`F�{E��F�q�pARxxPY�aSHFT͢�qA�AX_SHOR($�>��6 @$GqP9E���OVR���aRZPI@P@$U?r *a�AYLO���j�I��"��Aؠ��ؠERV��Qi�[Y)��G�@@R��i�e��i�R�!=P�uASYM���uFqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P��֊WOR�@M���k0SMT��G��G1R��3�aPA�@���p5�'�H � :j�A�TOCjA7pyP]Pp$OPd�O��C�%�p�O,!��RE.pR�C�A�O�?��Be5pR��EruIx'QG�e$P�WR) IMdu�RR�_$s �05��B �Iz2H8�=�_A�DDRH�H_LE�NG�B�q�q:�x�Rj��So�J.�SS��SK������ ���-�SE*����HS�N�MN1K	�`j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ����Q8� ��OUPW3�bE_>�I��!q�a1�� ������|���������-���:���iIOX2S=�D�e��<]���L $��p��!_OFF[r_�P�RM_��aT�TP_�H��M (�pOBJ�"�pG�[$H�LE�C��>ٰN � 9�*��AB_�T��
�S��`�S��LV��KR�W"duHITCOU�?BGi�LO�q ����d� Fpk�GpsSS� ���HWh��wA��O.��`IN�CPUX2VISIO��!��¢.�á<��á-� �IOLN.)�P 87�R'�[p�$SL�bd P7UT_��$dp��Pz �� F_AuS2Q/�$LD���D�aQT U�0]P�Aa������PHYG�d��Z�Ͱ5�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp����x��ٶ%�UJ���S����NE�WJsOG�G �DIS��b&�KĠ��3T |���AV��`_�CTR<!S^�FLAGf2&�;LG�dU �n�:���3LG_SIZ���ň��=���FD��I����Z �ǳ� �0�Ʋ�@s��-ֈ�-ր=�-���-��0-�ISGCH_��Dq��N?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHrܵ�I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn瘱I�BU�FF1XY��PT�$�� �v��f�QL6q1YY��Pp �����pOS1�%2�3���_�0Z �  ��aiE��*��IDX�dP��RhrO�+��A&S�T��R��Yz�<! _Y$EK&CK+����Z&m&KF�1[ L��o�0��]PL� 6pwq�t^����t�7�?_ \ �`�Р瀰�7��#�0C��]{ ��CLDP��>;eTRQLI�jd8.�094FLGz�0�r1R3�DM�R7��LqDR5<4R5ORG.� ��e2(`���V�8.��T8<�4�d^ �q�<4(��-4R5S�`T00m���0DFRCLM�C!D�?�?3I@��M9IC��d_ d����RQm�q�DSTB	�  �Fg�H�AX;b �H�LE�XCESZr�rBMup�a`Z��B;d��rB`��`a��F_�A�J��$[�O�H0K��db \��ӂS�$�MB��LIБ}SREQUIR�R>q�\<Á�XDEBU��oAL� MP�c�ba��Ph؃ӂ!BoAND�ф�`�`d�҆�c�cDC1��IN�����`@�(h?Nz�@q��o�w �SPST8�w e�rLOC��RI�p�EX�fA��p��AoAODAQnP�f X��ON��[rMF�����f)�"�I��%�e��T��FX�@IGG� g �q��"E�0��#���$R�a%;#7y���Gx��VvCPi�DAT	Aw�pE:�y��RF����NVh t W$MD�qIё)�v+�tń�tH�`�P�ux�|��sANSW}�P�t�?�uD�)�b��	@Ði �@C�U��V�T0�eRR2�j Dɐ�Qނ~�Bd$CALI�@�F�G�s�2�RI�N��v�<��NTE���kE���,��b����_Nl��ڂ���kDׄRm�DIVFiFDH�@ـn��$V��'c!$��$Z������~�[��oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS�@#2L  �Ė83ಀ����� ��PAT!H��������3̒Vp�A_�Q�.�4�B��Cᐈ�_MGh��$DDQ���G�$FWh��p��m������b�DE��PPAB�NԗROTSPE!ED����00J�Я�8��@��̐$US�E_��P��s�S�Y��c�A kqYNru@Ag��OFF�qn�MOUN�NGg��K�OL�H�INC *��a��q��Bj�L@�BENCS��q�BđX���D��IN#"I̒0��4�\BݠVEO�w�>Ͳ23_UPE�߳/LOWL���00����D���BwP���� �1RCʀƶMO3SIV�JRMO���@�GPERCH  �OV��^��i� <!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸUPp������TRKr�>"AYLOA'a��  Q-�̒<�1Ӣ`0 ���RTI$Qx�0 MO ���МB R�0J��D���s�H����b�DU�M2(�S_BCKLSH_C̒��>� =�q�#�U��ԑ���2�<t�]ACLALvŲp�1n�P�CHK00:'%SD�RTY4�k���y�1�q_6#2�_�UM$Pj�Cw�_�S�CL��ƠLMT_OJ1_LO��@���q��E�����๕�幘SPC��7���L���PCo���H� ȰPU�m�C/@�"XT\_�c�CN_��N��Le���SFu���V��&#����9�̒��=�C�u�SH6#��c��� �1�Ѩ�o�0�͑
��f_�PAt�h�_Ps�W�_10��4�R�01D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�sR0Hљ��_W��-ԁ_=��C��I��I*�I�II�F�`�aJLA.�1[�VC��0�D�BO1U�@i�B\JRKU��~	@DBL_SMd�:BM%`_DLC�BGRV��C��I���H_� �*CcOS+\�(LN� 7+X>$C�9)I�9)u*c,)�Z2 HƺcMY@!�( "TH&-��)THET0�N�K23I��"=�A C-B6CB=�C�A�B�(261C�616SB8C�T25GTS QơC��aS$" �4c#<�7r#$DUD�EX��1s�t��B�6���AQ�|r�f$NE�DpI B U�\B5��$!��!�A�%E(G%(!LCPH$U�2׵�2SX pCc%pCr%�2�&�C�J�&!�VAHV6H3�YLUVhJVuKV�KV�KUV�KV�KV�IHAH@ZF`RXM��wXuKH�KUH�KH�KH�KH�I�O2LOAHO�YWNO�hJOuKO�KO�KO*�KO�KO�&F�2#1�ic%�d4GSPBA?LANCE_�!�c�LEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%�Ċ1ky�UTO_<?�jT1T2Cy��2N&�v�ϰctw�gѠp�0Ӓ~���T��O����� INSEGv�!�REV�v!���gDIF��1l�w6�1m
�OB�q
����MIϰ1��L�CHWAR����A�B&u�$MEC�H,1� :�@�U�AX�:�P��Y�G$�8pn� 
Z��|���RO�BR�CR̒��N��'�MSK_�`�f�p P Np_���R����΄ݡ�1 ��ҰТ΀ϳ��΀"��IN�q�MTC�OM_C@j�q � L��p��$ONORE³5����$�r 8� GRl�E�SD�0ABF��$XYZ_DAx5A���DEBU�qXI��Q�s �`$�wCOD�� ���k�F�f�$BU�FINDXР � ��MOR��t $-�U��)��rРB��Ӱ��Gؒu� � $SIMULT ��~�� ����OBJE�` �AD�JUS>�1�AY_	Ik��D_����C��_FIF�=�T � ��Ұ��{��p� ��З��p�@��D�FRiI��ӥT��RO� Ұ�E���͐OPsWO�ŀv0���SYSBU�@ʐ$�SOP����#�U<"��pPRUN�I�PA�DH�D����_OU�=��qn�{$}�IMAG��iˀ�0P�qIM��Ơ�IN�q���RGOVRDȡ:���|�aP~���Р�0L_6p0���i��RB���0e��M���EDѐ*F� ��N`M*����鷀˱SL�`ŀw� x $OVS�L�vSDI��DEXm�g�e�9w�����	V� ~�N���w�����Ûǖȳ�M�̐ ���q<��� x �HˁE�F�ATUS
���C�0àǒ�çBTM����If�¿�4����(�ŀy �DˀEz�g���PE��r�����
���EXE��V��E�Y�$Ժ �ŀz @ˁ��UP�{�h�$�p��XN����9�H� ��PG"�{ h �$SUB��c�@_���01\�MPWAI2��P����LO��<��F�p�$RCV?FAIL_C�f��BWD"�F���DE�FSPup | Lˀ`�D�� U�UNI��S���RX`���_L�pP��%�P�ā}��� @B�~���|��`ҲN�`�KET��y���Pԙ $�~���0SI�ZE��ଠ{���S�<�OR��FORMAT/p � F���r�EMR��y�UX8����PLI7�ā�  $�P_SWI������_PL7�AL_ S�ސR�A��B��(0C��Df�$E�h����C_=�U�� � � ���~�J3�0�����TIA4��5��6��MOM������h �B�AD��*��* PU70NARW��W 
R������ A$PI�6���	�� )�4l�}69��Q����c�SPEED�PG q�7�D�>D�� ��>tMt[��SAM�`痰>��MOV���$��p �5��5�D�1�$2�������{�Hip�IN?,{� F(b+=$�H*�(_$�+�+GAMM�f�1{�$GET��ĐH��D����
^pLIB�R�ѝI��$HIB��_��Ȑ*B6E��b*8A$>G086LW= e6\<G9�686��R���ٰV��$PGDCK�Q�H�_����;"��z�.%�7��4*�9� �$IM_SRO��D�s"���H�"�LE��O�0\H��6@�p@�U� �ŀ�P�q?UR_SCR�ӚA�Z��S_SAVEc_D�E��NO��CgA�Ҷ��@�$��� �I��	�I� %Z[�  ��RX" ��m���" �q�'"�8�H ӱt�W�UpS����
T�M��O㵐.'}q ��Cg���@ʣ�ߑ��BM�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PLM���	� 0h�H�{�%X��O��z�Z�eT�M���� pS��C��O__0_B_�a:��_%�� |S��� �@	�v��v �@��ȯw�v��EM��% (-�cu�B�ː��ft�P��PM��QU.� �U�Q��A�f�QTH=�HOLޫ�QHYS�ES��,�UE��B��O.#��  -�P0�|�`gAQ���ʠu�Z���ŀ�ɂv�-�A;ӎ�ROG��a2�D�E�Âv�_�ĀZ�INFO&��+�����b� �킍 =((@SLEQ/�#����@O�o����S`c0O�0�0�1EZ0NUe�_�A�UT�Ab�COPY���Ѓ�{��@M��N@�����1�P�
� ���RGI�����X_�Pl�$�����`�W��P��j@�G����EXT_CYCBtb���p����nh�_NA�!$��\�<�RO�`]��� � m��PO�R�ㅣ���SRV�t�)����DI �T_l���Ѥ{�ۧ��ۧT �ۧ5٩6٩7٩I8����S�B쐒��K$�F6���PqL�A�A^�TAR�@�@E `�Z���9�n�d� ,(@FLq`Lh��@YNL���M�=C���PWRЍ�z쐔e�DELAѰ��Y�pAD#qX� ��QSKIP��� ĕ�x�O�`NT2!� ��P_x�-� ǚ@�b�p1�1� 1Ǹ�?� �?��>���>�&�>�3�>�9��J2R;쐖 46��EX� TQ���� ށ�Q���[�KFд����RDCIf� �U`�X}�R�#%M!�*�0�)��$RGEA�R_0IO�TJBFcLG�igpERa�TC݃������2T�H2N��� 1��b��Gq T�0 �����M���`I�b����REF�1��� l�h��ENsAB��lcTPE?@ ���!(ᭀ����Q �#�~�+2 H�W���2�Қ���"�4�F�X�j�3�қ{��︱����� ��4�Ҝ��
��.�@�R�
j�5�ҝu�������(����j�6�Ҟ���(:Lj�7�ҟ�o�����j�8�Ҡ��"4F^j�SMSK����)�a��E�A����oMOTE�������@ "1��Q�IO��5"%I��P��PO9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C��>%/S232%�Sb�i�DEVICEUS�#�R�RPARIT|�!OPBIT�Q���OWCONT�R��Qⱓ�RCU�� M�SUXTAS�K�3NB��0�$TA;TU�P�"@@R쐦F�6�_�PC}��$FREEFR�OMS]p�ai�GE�TN@S�UPDl�A�RB�#P%0����� !m$USAࢰ�az9�L�ERI��0f��pRY�5~"_ľ@f�P�1�!�6WR	K��D9�F9Х?FRIEND�Q4b�UF��&�A@TOO�LHFMY5�$L�ENGTH_VT��FIR�pqC�@�yE� IUFIN�R:���RGI�1�OAITI:�xGX�l�I�FG2�7G1a�0���3�B�GPRR�DA���O_� o0e�I1R�ER�đ�3&���TCp���AQJV �G|�.2���F��1�!d��9Z�8+5K�+5�� ��y�L0�4�X ��0m�LN�T�3H@z��89��%�4�3G��IW�0�W�RdD� Z��Tܳ�pK�a3d��{$cV 2��`H�1��I1H�02K2sk3K3Jci�a I�i�a�L��SL��RS$Vؠ�BV�EVk���AbQ*R��� � ,6Lc���9V2F{/P�:B��PS_�Et��$rr�C�ѳ$A0��wPR���v�U�cSk�� {�73�1��G� 0���VX`�!�tX`�\`�0P�Ё��
�5SK!� �"-qR��!0���z�MNJ AX�!h�A�@�LlA��A�THIC��1�������1TF�E���q>�IF_C	H�3A�I0�����G1�x������9��Ɇ_JF҇PR|(���RVAT�� �-p��7@�����DO�E��COU�(��AXIg��O�FFSE+�TRIG�SK��c���Ѽ�e��[�K�Hk���8�IG#MAo0�A-��ҙ��ORG_UNEV���� �S�쐮�d �$�������GROU��ݓTqO2��!ݓDSP���JOG'��#	�_P'�2OR���>P67KEPl�IR�0�2PM�RQ�AP�Q���E�0q�e���SYS�G��"��PG��BRAK*Rd�r�3�-���0����ߒ<pAD��ݓ�J�BSOC� N��DUMMY14��pN@SV�PDE_�OP3SFSPD�_OVR��ٰC�O��"�OR-��Nı0.�Fr�.��OV��SFc�2�f��F���!4�S��RA�"L�CHDL�REC�OV��0�W�@M�յ�RO3��9_�0� @�ҹ@�VERE�$OF�S�@CV� 0BWD�G�ѴC��2j�
�T�R�!��E_F�DOj�MB_CM4��U�B �BL=r0�w�=q�tVfQ��x0spd��_�Gxǋ�AM��`k�J0������_M���2{�#�8$CA��{Й���8$HB�K|1c��IO��8.�:!aPPA"�N��3�^�F���:"�DVC_DB�C��d�w"����!��1���ç�y3����ATIO� �q0�UC�&CAB�BS�PⳐ�P�Ȗ��_0c�S�UBCPUq��S �Pa aá�}0�Sb��c���r"ơ$HW_AC���:c��IcA�A~-�l$UNIT��l��ATN�f�����CYCLųNEC�A��[�FLTR_2_FI���(��}&Ɩ�LP&�����_S[CT@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb��r�: _T��PROX��O�� EM�_�r��8u�q u��q��DI�0e�RAOILAC��}RMƐCLOԠdC��:anq���wq����PR��S�LQ�pfC�ѷ 	���FUNCŢ�rRINkP+a�0 ��!3RA� >R 
Я8�ԯWAR�#BLFQ��A�����DA�����LDm0�aB9�2�nqBTIvrb8ؑ���PRIAQ1�"AFS�P�!���𰠓�`%b���M�I1U�DF_j@��y1�°LME�FA�@H�RDY�4��Pn@R�S@Q�0"�MUL�SEj@f�b�q ��X��ȑ���m$.A$�1$c1�Ó���� x~�EG�0ݓ�q!cAR����09LB��%��AXE��RKOB��W�A4�_�-�֣SY���!6��&S&�'WR���-1����STR��5�9�E�� 	5B��=Q�B90�@6������O�T�0o 	$�A�RY8�w20���	�%�FI��;�$LGINK�H��1�aI_63�5�q�2XYZ"��;�q�3@�R�1�2�8{0B�{D��� CFI��6G��
�{��_J��6��3aO�P_O4Y;5�QT�BmA"�BC
�z�D�U"�66CTURN3�vr�E�1�9���GFL�`���~ �@��5<:7�� 1��?0K�Mc�68�Cb�vrb�4�ORQ ��X�>8�#op�������wq�Uf�����TOVE�Q��M;�E# �UK#�UQ"�VW�ZQ �W���Tυ� ;��� �QH�!`�ҽ��U�Q�W`keK#kecXER�
�	GE	0��S�dAWaǢ:D���7!�!AX�rB!{q ��1uy-!y�p z�@z�@z6Pz\P z� z1v�y� y�+y�;y�Ky� [y�ky�{y��y�qޜyDEBU��$ ����L�!º2WG` � AB!�,��SV���� 
w���m� ��w����1���1���A ���A��6Q��\Q���!��m@��2CLAB�3B�U�����S 7 ÐER��
0� � $�@� A6ؑ!p�PO���Z�q0w�^�_MRA�ȑ� d  T�-�ERR��STYz�B�I�V3@��cΑTOQ�d:`L�� �d2�]�X�C�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	�SFZN�_CFG_!� 4 ��?º�|�ų����@��ȲW p ��\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(�����!�s�Q�g�P{RV H�ELLĥ� }56�B_BAS!�GRSR��ԣo �#QS��[��1r�%��U2ݺ3ݺ4ݺ5ݺ�6ݺ7ݺ8ݷ��R�OOI䰝0�0NL�K!�CAB� ��A[CK��IN��T:��1�@�@ z�m�_P�U!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KcARӑ��RE~���P��(��QUE������P
��CST?OPI_AL������0&���㰑�0SE�Ml�b�|�M��d�T�Y|�SOK�}�DI������(���_T}M\�MANRQ���0E+�|�$KEYSWITCH&�	���HE
�BE�AT����E� LE(Ғ���U��FO���|��O_HOM��O�REF�PPR�z��!&0��C+�OA�ECO��B�rIOCM�D8׵��]���8�` � �D�1����U��&�M�H�»P�CFORC<��� �'�����OM�  � @�V��|�U,3P� 1(-�`� 3-�4���NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F��V ��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7s�VP�U�PD��  ���|�԰��YSLO>Ǣ� � z��� ����o�E��`>�^t���АALUץ����C�U���wFOqID_YL�ӿuHI�zI�?$FILE_���tf��$`�JvSA���� h���E_B�LCK�#�C,�D_CPU<�{�<�o�����tJr��R ;��
PW O�[ ��LA��S��8������RUNF�Ɂ ��Ɂ����F�ꁡ�ꁾ���TBCu�C�� �X -$�LENi��v������I��G�LOWo_AXI�F1�
�t2X�M����D�
 ���I�� ��}�T#OR����Dh��� L=��⇒�s���#�_MA`�ޕ���ޑTCV����T ���&��ݡ����J�$����J����Mo����J�Ǜ �������2��� v�����F�JK��VKi�ΡvњΡ3��J0�ңJ�JڣJJ�AAL�ң�ڣ��4�5z�&�N1-�9����J��L~�_Vj������� ` �GGROU�pD��B�NFLIC��R�EQUIREa�E�BUA��p����2�¯�����c��� \��APPR���C���
�EN��CLOe��S_!M v�,ɣ�
���o� ���MC�8&���g�_MG�q��C� �{�9���|�B;RKz�NOL��|�:� R��_LI|���$��k�J����P
��� ڣ�����&���/���Q6��6��8��r�>��� ��8��%�W�2�e�PATHa�z�p�z�=�vӥ��ϰ�x�CN=�CA������p�IN�U�C��bq��CO�UMB��YZ������qE%����2������PAYwLOA��J2L3pOR_AN��<�L���F�B�6�R�{�R_F�2LSHR��|�L�OG��р��ӎ���ACRL_u��������.���H�p�$H�{���FLEX
���J�� : �/����6�2�����;�M�_�F16�����n���������ȟ��E ҟ�����,�>�P� b���d�{������ ������5�T��X��v���Eťm Fѯ������� &�/�A�S�e�+p�x�� � �������j�4pAT����n�EML  �%øJ����ʰJE��CTR,�Ѭ�TN��F&��HAND_VB[q
�pK�� $�F2{�6� �rSW�i��("U��� '$$Mt�h�R��08@��@<b 35��^6A�p 3�k��q{9t�A�̈p
��A��A�ˆ0��U����D��D��P��G��IST��$A��$AN��DYˀ�{�g4 �5D���v�6�v��5� ���^�@��P��� ��#�,�5�>�(#�� &0�_�ER!V<9�SQASYM��] 	�����x��ݑ���_SHl�������sT@�(����(�:�JA����S�cir��_V�I�#Oh9�``V_�UNI��td�~�J ���b�E�b��d��d �f��n���������u�N���(!�H̟�����"CqENL� �pDI��>�Obtq D�Dpx�� �
�2IxQA�q��q���-��s �� s�����{ ��OMME���rr/�TVpP�T�P ���qe�i� ���P�x ��yT�Pj�� $DUMM�Y9�$PS_f��RFq�sp$:�� s���!~q�c X����K�STs��ʰSBR��M2�1_Vt�8$SV_ERt�O��z���WCLRx�A  O�r�?p? Oր � �D $GLOB���#LO��Յ$�po��P�!SYS�ADR�!?p�pTC}HM0 � ,�����W_NA���/�e�os�TSR~��l (: ]8:m�K6�^2m�i7 m�w9m��9���ǳ��� ����ŕߝ�9ŕ�� �i�L���m��_�_��_�TD�XSCRE��ƀ�� ��ST�F���}�pТ6��sq] _v AŁ� 9T����TYP�r�@K��u�!u���-O�@IS�!��tvC�UE{t� �����H�S���!RSM�_�XuUNEXCcEPWv��CpS_�� {ᦵ�ӕ���÷����COU ��� [1�O�UET�փr|���PROGM� {FLn!$CU��cPO*q��c�I_�p}H;� � 8��.N�_HE
p��Q�~�pRY ?����,�J�*��;�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� ��C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!$sqVSHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3��H���w�2u�b�V�rzu��%�DJU��~|#�WAIT�������%ONE���YBOư ?�� $@p%�vC�SBn)TPE��NEC��x"�$t$��.�*B_T��R��% �qR� ���sB�%�tM�+��t�.�F�R!�݀��OPm�MAS��_DOG�OaT	�D����C3S�	�O2DELAY���e2JO��n8E��Ss4'#�J�aP6%�����Y_��O2$��2���5���`? �PZ�ABCS��  �$�2��J�
sp��$$CLAS�����Aspb�'@@VIRT��O.@gABS�$�1 <E�� < *AtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v�p����M@[�AXLրt�&A�dC  ����IN��ā��PRE������LA�RMRECOV c<I䂥�NG��� \K	 A �  J�\�M@PPL�IC�?<E��E�Hand�lingTool� �� 
V7.�50P/28[� � �X0��
��_SW�� UPn*A� ��F0ڑ䢒��A���� 20��*A����:���(<FB 7DA5��� '@Y0�@����None엃���� ���T�K*A4I/Wxl�_��V��t��g�UTOB��ค����HGAPCON8@��LA��U��oD 1<EfA���������� /Q 1שI Ԁ��Ԑ�:�i�n�����#B)B g���\�HE��Z�r�HTTHKY��$BI�[�m��� ��	�c�-�?�Q�o�u� �ϙϫϽ�������� _�)�;�M�k�q߃ߕ� �߹��������[�%� 7�I�g�m����� ��������W�!�3�E� c�i�{����������� ����S/A_e w������� O+=[as� ������K// '/9/W/]/o/�/�/�/ �/�/�/�/G??#?5? S?Y?k?}?�?�?�?�? �?�?COOO1OOOUO gOyO�O�O�O�O�O�O ?_	__-_K_Q_��(��TO4�s���DO_CLEAN��e��S�NM  9� �9oKo]ooo�o�DSPDRYR�_&%�HI��m@&o�o �o#5GYk} ����"���p�Ն# �ǣ�qXՄ���ߢ��g�PLUGGpҠ�Wߣ��PRC�`B`9��o�=��OB��oe�SEGF��K������o%o�����#�5�m���LAP�oݎ���������� џ�����+�=�O�|a���TOTAL�|.���USENUʀ�׫ �X���R(�R�G_STRING� 1��
�kM��Sc�
���_ITEM1 �  nc��.�@�R�d� v���������п������*�<�N�`�r��I/O SIG�NAL��Tr�yout Mod�e�Inp��S�imulated��Out���OVERR�` =� 100�In� cycl����Prog Abo�r�����Sta�tus�	Hea�rtbeat��MH FaulB�K�AlerUم�s� �ߗߩ߻��������� �S���Q� �f�x�������� ������,�>�P�b��t�������,�WOR ������V��
. @Rdv���� ���*<N`PO��6ц�� o�����// '/9/K/]/o/�/�/�/��/�/�/�/�/�DEV�*0�?Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O>�OPALTB��A ���O�O__,_>_P_ b_t_�_�_�_�_�_�_��_oo(o:o�OGRI�p��ra�OLo�o�o �o�o�o�o*< N`r������`o��RB���o� >�P�b�t��������� Ώ�����(�:�L��^�p����PREG �N��.�������� *�<�N�`�r������� ��̯ޯ���&��Ϳ�$ARG_��D ?	���i���  �	$��	[�}�]}���Ǟ�\�S�BN_CONFIOG i��������CII_SA_VE  ��۱�Ҳ\�TCELLSETUP i��%HOME_I�O�͈�%MOVq_�2�8�REP����V�UTOBAC�K
�ƽ�FRA:\�� ��Ϩ���'`!��������  ����$�6�c�Z�lߙ��Ĉ���������� ���!凞��M�_�q� ����2�������� �%�7���[�m���� ����@�������!3E$���Jo��������INI��@��ε��MESSAG����|q��ODE_D$����O,0.��P�AUS�!�i� ((Ol��� ����� /�/ /$/Z/H/~/l/�/�'�akTSK  �q�����UPDT�%�d0;WS�M_CF°i��еU�'1GRP Y2h�93 |�B���A�/S�XSCRDv+11
1; ����/�?�?�? OO $O��߳?lO~O�O�O �O�O1O�OUO_ _2_�D_V_h_�O	_X���G�ROUN0O�SU�P_NAL�h�	��ĠV_ED� 1�1;
 �%-BCKEDT-�_0`�!oEo%���a(��o�����ߨ���e2no_˔o�o�b���ee�o"�o�oED3�o�o ~p[�5GED4� n#�� ~�j���ED5Z��Ǐ6� ~p���}���ED6�� ��k�ڏ ~G���!�3�ED7��Z��~� ~p�V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W��Ư
}3�����CRo�����3�տ@�����P�PNO_D�EL�_�RGE_U�NUSE�_�TLA�L_OUT �q�c�QWD_AB�OR� �΢Q��IT_R_RTN����ONONSe����CAM_PAR�AM 1�U3
� 8
SONY� XC-56 2�34567890��H � @����?���( SАV�|[r؀~�X�HR5k�|U�Q��߿�R57����A�ff��KOW�A SC310M�|[r�̀�d @6�|V��_�X� ����V��� ���$�6���Z�l��CE_R�IA_I857�F�1��R|]]��_LIO4W=V� ��P<~�F<��GP 1�,����_GYk*Cg*  ��C1� �9� @� G� �CVLC]� d� l� Es�R� ��[�Um� v� � �� _�� C�� �"��|W��7�HEӰO�NFI� ��<G_�PRI 1�+ P�m®/���������'CHKPA�US�  1E� ,�>/P/:/t/^/ �/�/�/�/�/�/�/?�(??L?6?\?�?"OƩ����H�1_MkOR�� �0�5 	 �9 O�?�$OOHO6K�2	��H�=9"�Q?55��CR�PK�D3P����>��a�-4�O__|Z
�OG_�7�P O�� ��6_��,xV�A�DB���='�)
�mc:cpmidcbg�_`��S:�)�	���Yp�_)o�S`�BBi�P�_mo8j�)�Koo�oV9i�)��og�o�o�m�of�oGq:�I�ZDEF �f8��)�R6pbuf.txtm�]nd�@����# 	`)н��A=L���zM-C�21�=��9����4�=�n׾�C�z  BHBCCo��C|��Cq�D��C�?��C�{iSZE@�D��F.���F��E⚵F,E�ٙ��E@F�N�IU���I?O�I<�#I6�I�I�SY���vqG����Em�)�.���)�)��<�q�G�)x2��Ң �� a��D�j���E�e��E�X�EQ�E�JP F�E�F� G�ǎ�^F E�� F�B� H,- Ge��H3Y����  >�33 ����xV  n42xQ@��5Y��8B� A�AST<#�
�� �_'�%��wR_SMOFS���~�2�yT1�0DE ��O c
�(�;�"�  <�6�z��R���?�j�C4R��SZm� W���{�m�C��B-G�CR�`@$�q��T{��FPROG %i����c�I��� �����f�KEY_TB�L  �vM�u� ��	
�� �!"#$%&'(�)*+,-./0�1c�:;<=>?�@ABC�pGHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������p���͓���������������������������������耇�������������������s��!j�LCK��x.�j���STAT����_AUTO_D�O���W/�IND�T_ENB߿2R���9�+�T2w�XS�TOP\߿2TRL^l�LETE�����_SCREEN �ikcs�c��U��MMEN�U 1 i  <g\��L�SU+� U��p3g������ ������2�	��A�z� Q�c������������� ��.d;M� q������ N%7]�m ���/��/J/ !/3/�/W/i/�/�/�/ �/�/�/�/4???j? A?S?y?�?�?�?�?�? �?O�?O-OfO=OOO �OsO�O�O�O�O�O_��O_P_Sy�_MA�NUAL��n�DB;COU�RIG��ٟDBNUM�p���<���
�QPXWO_RK 1!R�ү��_oO.o@oRk�Q_�AWAY�S��G�CP ��=��df_CAL�P�db�RY��������X_�p 1">�� , 
�^����o xvf`MT�I�^�rl@�:sONT�IM�������Zv�i
õ�cMOT�NEND���dRECORD 1(R�qa��ua�O��q ��sb�.�@�R��x Z�������ɏۏ� ����#���G���k�}� ����<�ş4��X�� �1�C���g�֟���� ����ӯ�T�	�x�-� ��Q�c�u�������� ��>����)Ϙ�M� ��F�࿕ϧϹ���:� ������%�s`Pn&�]� o��ϓ�~ߌ���8�J� ����5� ��k��� �ߡ��J�����X�� |��C�U�������� ���0�����	��db�TOLERENC�qdBȺb`L����PCS_CFG �)�k)wdM�C:\O L%04�d.CSV
�pcl�)sA �CH� z�p)~���h�MRC_OUT �*�[�`+P S�GN +�e�r���#�10-MA�Y-20 09:�21*V17-FE}Bj19:09�k PQ�8��)~�`pa��m��PJP���VERSIO�N SV�2.0.8.|EF�LOGIC 1,^�[ 	DX�P�7)�PF."PROG�_ENB�o�rj U�LSew �T�"_?WRSTJNEp�V��r`dEMO_OPT_SL ?	�e�s
 	R575)s7)�/??*?�<?'�$TO  ��-��?&V_@pE�X�Wd�u�3PA�TH ASA�\�?�?O/{ICTZ�aFo`-�gd>segM%&A�STBF_TTS��x�Y^C��SqqF��PMAU� t/XrMKSWR.�i6.|S/�Z!D_N�O 0__T_C_x_g_�_�t�SBL_FAUL�"0�[3wTDIAbU 16M6p�A�123456�7890gFP ?BoTofoxo�o�o�o �o�o�o�o,>�Pb�S�pP�_ ���_s�� 0`� ����)�;�M�_� q���������ˏݏ�|)UMP�!� �^�TR�B�#+��=�PMEfEI�Y_�TEMP9 È��3@�3A v�UNI��.(YN_BRK� 2Y)EMG?DI_STA�%W�ЕNC2_SCR 3��1o"�4� F�X�fv���������#��ޑ14���@�)�;�����ݤ5�����x�f	u� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/߭P�b� t�� ��xߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N���r��� ������������ &8J\n��� �����"`� FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/4?,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O?�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�O�O�o �o�o
.@Rd v������� ��*�<�N�`�r��� �o����̏ޏ���� &�8�J�\�n����������ȟڟ����H�E�TMODE 16v��� ���ƨ
R�d�v�נR�ROR_PROG7 %A�%�:߽��  ��TABLE  A�������#�L�RRSEV_?NUM  ��Q���K�S���_�AUTO_ENB�  ��I�Ϥ_N�Oh� 7A�{��R�  *����J��������^�+��pĿֿ迄�HISO����I�}�_ALM �18A� �;�����+�e�wωϐ�ϭϿ��_H���  A���|��4��TCP_VER �!A�!����$E�XTLOG_RE�Q��{�V�SI�Z_�Q�TOL  ���Dz��A= Q�_BWD���иr���n�_DI�� 9��}�z���<m���STEP����|4��OP_DO����ѠFACTO�RY_TUN�d�G�EATURE �:����l��Handlin�gTool �� � - CEn�glish Di�ctionary���ORDEA�A Vis�� M�aster���9�6 H��nalo�g I/O���H�551��uto �Software� Update � ��J��mati�c Backup~��Part&��ground E�dit��  8\�apCame�ra��F��t\j�6R�ell���LwOADR�omm���shq��TI" ��co��
! yo���pane��� 
!��ty�le selec]t��H59��nD�~��onitor��48����tr��R�eliab���a�dinDiagnos"����2��2 ual Che�ck Safet�y UIF lg�\a��hance�d Rob Se�rv q ct\���lUser F�rU��DIF��E�xt. DIO 6��fiA d��wendr Err YL@��IF�r�ನ  �П�90��F�CTN Menu�Z v'��74� T�P In��fac�  SU (�G=�p��k E�xcn g�3��High-Sper wSki+�  sO��H9 � mmuni]c!�onsg�te�ur� ����V��y��conn���2��EN��Inc=rstru����5.fdKA�REL Cmd.� L?uaA� O~�Run-Ti� 'Env����K� ��u+%�s#�S/W���74��Licen�seT�  (A�u* ogBook�(Sy��m)��"�
MACR�Os,V/Off�se��ap��MH�� ����pfa5�M�echStop �Prot��� d��b i�Shif����j545�!x�r ��#��,[>�b ode Swiwtch��m\e�!�o4.�& pr�o�4��g��M?ulti-T7G����net.P{os Regi���z�P��t Fu9n���3 Rz1���Numx �����9�m�1�  Adju<j��1 J7�7�*� ����6tatu�q1EIKRD�Mtot��scove�� ��@By<- }uest1�$G�o� � U5\SNPX b"���<YA�"Libr��㈶�#�� �$~@h�p�d]0�Jts i?n VCCM����ĕ0�  �u!��2 �R�0�/I�08~��TMILIB�M� J92�@P�A�cc>�F�97�TgPTX�+�BRSQselZ0�M8 Rm��q%��692��Unexceptr �motnT  CcVV�P���KC�����+-��~K  I�I)�VSP CSXC�&.c�� e�"��� t�@We�w�AD Q�8bv9r nmen�@�KiP� a0y�0��pfGridAplay !� nh�@*��3R�1M-10iA�(B201 �`2�V"  F���sci�i�load��8�3 M��l����G�uar�d J85��0�mP'�L`���s�tuaPat�&]$C�yc���|0ori�_ x%Data'Pqu���ch�1���g`� j� RLJa�m�5���IMI �De-B(\A�cP"� #^0C  e�tkc^0assw�o%q�)650�Ap�U�Xnt��PvKen�CTqH�5�0�YELLOW� BO?Y��� Arc�0vis��C�h�WeldQci�al4Izt�Op�� ��gs�` 2@�a6��poG yRjcT1 NE�#HTf� xyWb��! �p��`gd`���p\� �=P��JPN ARCP*PR�A�� �OL�pSup̂fil�p��J�� n��cro�670�1�C~E�d��SS�pe.�tex�$ �P� �So7 t� ssa%gN5 <Q�BP:� 2�9 "0�QrtQCr��P�l0dpn������rpf�q�e�ppm�ascbin�4psyn�' pstx]08�HEL�NCL VIS �PKGS �Z@M�B &��B J8�@IPE GET_VAR FI?S_ (Uni� LU��OOL: ADD��@29.FD�TC4m���E�@DVp����`A�ТNO WT?WTEST �� �f�!��c�FOR ^��ECT �a!� �ALSE ALA�`�CPMO-13�0��� b D: H�ANG FROM�g��2��R709� DRAM AV�AILCHECK�S 549��m�V�PCS SU֐L_IMCHK��P�0~x�FF POS� �F�� q8-12 CHARS��ER6�OGRA ���Z@AVEH�AME��.SV��Вאqn$��9�m "y��TRCv� SHA�DP�UPDAT �k�0��STATI���� MUCH ����TIMQ MOTN-003���@OBOGUI�DE DAUGH໱�b��@$tou�� �@C� �0��PA�TH�_�MOVE�T�� R64��V�MXPACK M�AY ASSERyTjS��CYCL`��TA��BE CO�R 71�1-�AN���RC OPTI�ONS  �`��A�PSH-1�`fi	x��2�SO��B��XO򝡞�_T��	�i�j�0j��du�byz �p wa��y�٠H�I������U�pb X?SPD TB/�F�_ \hchΤB0����END�CE�06�\Q�p{ sma'y n@�pk��L} ��traff#��	� ��~1fro�m sysvar/ scr�0R� ��Nd�DJU���H��!A��/��SET GERR�D�P7�����NDANT S�CREEN UNREA VM �P�D�D��PA���R~�IO JNN�0��FI��B��GRwOUNנD Y��Т٠�h�SVIP� 53 QS��DI�GIT VERS���ká�NEW�� �P06�@C�1IMCAG�ͱ���8� �DI`���pSSU�E�5��EPLAN� JON� DELL���157QאD��CALLI���Q��m���IPND}�IMG N9 PZ�{19��MNT/���ES ���`LocR Hol߀=��2�P�n� PG:��=�M��can����С�: 3D mE2view d X���ea1 �0b�po;f Ǡ"HCɰ��ANNOT AC�CESS M c�pie$Et.Qs �a� loMdFle�x)a:��w$qmo+ G�sA9�-'p~0̿�h0pa��eJ AUTO-�0��!�ipu@Т<ᡠIA�BLE+� 7�a F�PLN: L�p�l m� MD<�V�I�и�WIT H�OC�Jo~1Qu�i��"��N��US�B�@�Pt & r�emov���D�vAxis FT_7�PGɰCP:�O�S-144 � h� s 268QՐO�ST�p  CRA�SH DU��$P~��WORD.$��LOGIN�P��P�:	�0�046 i�ssueE�H�:� Slow st�c�`6�����z��IF�IMPR��SPOT:Wh4����N1STY��0V�MGR�b�N�CA�T��4oRRE�� �� 58�1��:N%�RTU!Pe -M .a�SE:�@pp���$AGpL��m@�all��*0a�OC�B WA���"3 �CNT0 T9DW�roO0alarm8�ˀm0d t�M��"0�2|� o�Z@O�ME<�� ��E%  ;#1-�SRE��M��st}0g   �  5KANJI~5no MNS@��INISITA7LIZ'� E�f�cwe��6@� dr�@� fp "��SC�II L�afai�ls w��SY�STE[�i�� � � Mq�1QGro8�m n�@vA�����&��n�0q��R�WRI OF L|k��� \ref"��
�up� de-r�ela�Qd 03�.�0SSchőb�etwe4�INDo ex ɰTPa�#DO� l� �ɰ�GigE�sope�rabil`p l�,��HcB��@]�lye�Q0cflxz�8Ð���OS {�����v4pfigi GL�A�$�c2�7H� wlap�0ASB� �If��g�2 l\�c�0�/�E�� �EXCE 㰁�P����i�� o0��G�d`]Ц�fq�l lsxt��EFal����#0�i�O�Y�n�CL�OS��SRNq1NT^�F�U��FqKP~�ANIO V7/�¥�1�{����DBa �0��ᴥ�ED��DET|�'� �b�F�NLINEb�B�UG�T���C"RL�IB��A��ABC? JARKY@���� rkey�`IL����PR��N��ITG+AR� D$�R �Er *�T��a�U�0��h�[�ZE V�� TASK p7.vr�P2" .�XfJ�srn�S谥d�IBP	c���B/��BUS��UNN�� j0-�{��cR�'���LOE�DIVS�CULs$cb����BW!��R~�W`�P�����IT(঱t�ʠ�OF��UNE�Xڠ+���p�FtE���SVEMG3`N�ML 505� D�*�CC_SAFE��P*� �ꐺ� PE�T��'P�`�F  �!���IR����c Ri S>� K��K��H GUNCHGz��S�MECH��IM��T*�%p6u���tPORY LE�AK�J���SP�EgD��2V 74\GRI��Q�g��oCTLN��TRe `@�_�p ���EN'�IN������$���r��T3)�i�STO��A�s�L��͐X	���q��Y� ��CTO2�J m��0F<�K����DU�S��O���3 9�J F��&���SSVGN�-1#I���RSRwQDAU�Cޱ� �T6��g��� 3�]���BR�KCTR/"� �q\�j5��_�Q�S�qI{NVJ0D ZO�P ݲ���s��г�Ui ɰx̒�a�DUAL�� J50e�x�RV�O117 AW�T�H!Hr%�N�247�%�52��|�&aol� ���R���at�Sd��cU���P,�LER��iԗQ0�ؖ  S!T���Md�Rǰt�_ \fosB�A�0@Np�c����{�U���ROP 2�b�pB>��ITP4M��b !AUt c0< � �plete�N@�� z1^qR635� (AccuCa�l2kA���I) �"�ǰ�1a\�Ps ��ǐ� bЧ0P������ig\cba?cul "A3p_ �1��ն���eta�ca��AT���PC��`�����_p�.�pc!Ɗ��:�cicrcB���5�tl��Bɵ�:�fm+�Ί��V�b�ɦ�r�upf�rm.����ⴊ�x�ed��Ί�~�ped�A�D �}b�ptl�ibB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆Ϙ���c�Ӳ�5�1j>�����tcȐ�Ϣ	�r����mm 1���T�sl^0��T�m�ѡ�#�rm3��u8b Y�q�std}��3pl;�&�ckv�=߆r�vf�䊰��9�v1i����ul�`�04fp�q �.f���� daq; i Da�ta Acqui+si��n�
��4T`��1�89���22 DMCM oRRS2Z�75���9 3 R710,�o59p5\?T "��1 (D�T� nk@���� ����E Ƒȵ��Ӹ��etdmm ��ER�����gE��1�q\mo?۳�=( G���[(

�2�` �! �@JMAC�RO��Skip/Offse:�a���V�4o9� &qR6C62���s�H��
 6Bq8����9~Z�43 J77� =6�J783�o `��n�"v�R5�IKCBq2 PT�LC�Zg R�3; (�s, �������03�	зJ���\sfmnmc? "MNMC�����ҹ�%mnf�FM�C"Ѻ0ª etm�cr� �8����� ,[>D�f>   874\prdq>�,jF0���axi�sHProcess Axes e�wrol^PRA
��Dp� 56 J81�j�59� 56o6�� ���0w�690 998� [!IDV�1��2(x2��2ont �0�
����m2����?C��etis "ISD��9�� F/praxRAM�P�8 D��defB�,��G�isbasicHB�@޲{6�� W708�6��(�Acw:������D
�/,��AMOX�� ��DvE ��?;T��>Pi� RACFM';�]�!PAM�V �W�Ee�U�Q'
bU�75�.�ceN�e� nterfa�ce^�1' 5&!5�4�K��b(Dev am±�/�#���/<�Tazne`"DNEWE����btpdnui� �AI�_s2�d_rsono���bAs�fjN��bdv_arFvf�xhpz�}w��shkH9xstc��gAponlGzv{�ff��r���z��3{q'Td>pcOhampr;e�p� ^5977��	܀�4}0��mɁ�/�����l�f�!�pcchmp�]aMP&B�� �m�pev�����p�cs��YeS�� M/acro�OD��16Q!)*�:$�2U"_,x��Y�(PC ���$_;������o��J�g�egemQ@GEM�SW�~ZG�gesn�dy��OD�ndda��S��syT�Kɓ�Csu^Ҋ���n�m��<�L��  ���9:�p'ѳ޲��spotplusp���`P-�W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\f�eatu 0FEA�WD�oolo�s�rn'!2 p���a؝As3��tT.� (?N. A.)��!�e!�J# (j�,`��oBIB�oD -��.�n��k9�"K���u[-�_���p� "PSEqW����?wop "sEЅ� &�:�J������y�|� �O8��5��Rɺ��� ɰ[��X������ـ%�(
ҭ�q HL �0k�
�z�a!�B�Q�"(g�Q����� ]�'�.�����&���<�0!ҝ_�#��tpJ�H� ~Z��j�����y���� ��2��e������Z�� ��V��!%���=�]�p͂��^2�@iRV� Kon�QYq͋JF0B� 8ހ�`�	(^>�dQueue���X�\1�ʖ`�+F1tpv�tsn��N&��ftupJ0v �RDV�	�f��J1 Q���v��en��kvst�k��mp��btk�clrq���get����r��`kack�XZ��strŬ�%�st0l��~Z�np:!�`����q/�ڡ6!l��/Yr�mc�N+v�3�_� ����.�v�/\jF���� �`Q�΋ܒ�N50 (FRA��+�����fraparm���Ҁ�} 6�J6�43p:V�ELSE�
#�VAR $�SGSYSCFG�.$�`_UNITS 2�DG~°@�4�Jgfr��4A�@FRL-��0ͅ�3ې���L �0NE�:�=�?@�8 �v�9~Qx304��;�BPRSM~QA��5TX.$VNUM_OL��5��DJ�507��l� Functʂ"qwAP��琉�3 H�ƞ�kP	9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TP�PR���QA�prnaSV�ZS��AS8D�j510U�-�`cAr�`8 ��ʇ�DJR`�jYȑH  ��Q �PJ6�a2�1��48AA�VM 5�Q�b0 �lB�`TUP xb?J545 `b�`�616���0V�CAM 9�CwLIO b1�s5 ���`MSC8��
rP R`\s�STYL MNI�N�`J628Q  �`NREd�;@�`�SCH ��9pDCSU Mete�`�ORSR Ԃ�a0�4 kREIO�C �a5�`542�b9vpP<�nP�a�`�R�`7�`�M?ASK Ho�.r�7 �2�`OCO :��r3��p�b�p���r0X��a�`13\�mn�a39 HR�M"�q�q��L�CHK�uOPLG� B��a03 �q.��pHCR Ob�pC�pPosi�`fP6� is[rJ554��òpDSW�bM�D8�pqR�a37 }Rjr30 �1�s4 �R6�m7��52�r5 �2.�r7 1� P6����Regi�@T^�uFRDM�uSaq�%�4�`930�uS�NBA�uSHLB�̀\sf"pM�N{PI�SPVC�oJ520��TC�`�"MNрTMIL��IFV�PAC �W�pTPTXp6�.%�TELN N� Me�09m3�UECK�b�`U�FR�`��VCOR^��VIPLpq89q�SXC�S�`VVF��J�TP �q��Rw626l�u S�`�Gސ�2IGU�I�C��PGSt�\ŀH863�S�q������q34sŁ6�84���a�@b>�3� :B��1 T��9�6 .�+E�51 �y�q53�3�b1 ̛��b1 n�jr9 <���`VAT ߲�q�75 s�F��`�sA�WSM��`TOP u�ŀR52p���a�80 
�ށXY �q���0 ,b�`8855�QXрOLp}��"pE࠱tp�`LCyMD��ETSS�挀6 �V�CPEs oZ1�VRCd3�
�NLH�h��0011m2Ep��3 f��p���4 /165CR��6l���7PR���008 tB��9 o-200�`U0�p�F�1޲1 ��޲2 L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�J�?7 rbcfA�L��8\PC����"�32�m0u�n�K�Rٰn�5� 5EW
n�99 z��40 kB���3 ��6ݲ�`00�iB/��6�u��7�u��8 µ������s�U0�`�t �1 0�5\rb��2 E@���K���j���5˰��60��a�HУ`:Ł63�jAF�_���F�7 ڱ݀H�8�eHЋ�&�cU0��7�p���1u��8u��9 c73������D7� r��5t�97 ��E8U�1��2��1�)1:���h��1np�"���8(�U1��\pyl��,࿱v ��B�854��1V���D�-4��im��1�<����>br�3pr�48@pGPr�6 B����$�p��1����1�`͵�155ض157 �2��62�S����B��1b��2����1Π2"�2���B6`�1<c�4 7B�5i DR��8_�B/���187 uJ�8 ;06�90 rBn��1 (��202 /0EW,ѱ2^��2��90�U2�p�2��S2 b��4��2�a�"RB����9\�U�2�`w�l���4 6	0Mp��7������b�,s
5 ��3����<pB"9 3 ����l�`ڰR,:7 �2��V�2��5���2^H��a^9���qr�����n�5����5᥁""�8a�Ɂ}�5B���5����`UA���� ���86 �6 S�0�5�p�2�#�52�9 �2^�b1
P�5~�2`���&P*5��8��5��u�r!�5��ٵ544��%5��R�ąP nB^,z�c (�4���L���U5J�V�5��1�1^��%�����5 b21��gA���58W82� r�b��5N�E�589�0r� 1�95  �"������c8"a��|�L ���!J"5|6���^!�6��B�"8P�`#��+�8%�6B��AME�"1 iCN��622�Bu�6V���d� 4��84�`A�NRSP�e/S� C�5� �6� ��� \� �6� �V� 3�t��� T20CA�R��8� Hf� 1D�H�� AOE� ��� ,[|�� a�0\�� �!64K���ԓrA� �1 (M{-7�!/50T� [PM��P�Th:1�C��#Pe� �3�0� 5>`M75T"� �D�8p� �0Gc� u�4|��i1-710i�1B� Skd�7j�?6�:-HS,� �RN�@��UB�f�X�=m7C5sA*A6an���!X/CB�B2.6A �0 ;A�CIB�A�2�QF1�U�B2�21� /70�S� �4����Aj1��3p���r#0 B2\m*A@C��;bi"�i1K�u"A~AAU� imm7c7��ZA@HI�@�Df�A�D5*A��E� 0TkdR1�35�Q1�"*�@�Q�1�QC )P�1*A�5*A�EA�5XB�4>\77
B7=Q �D�2�Q$B�E7�C�D%/qAHEE�W7�_|` jz@� 2�0�Ejc�7�`�E"l7�@7@�A
1�E�V~`�W2%Qr�R9ї@0L_�#�����"A���b��H3s=rA/2�R5nR 4�74rNUQ1ZU�A�sw\m9
1M92L2��!F!^Y�ps� 2c1i��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHsXBSt62�q`s������ ��Pxq3530_*A3I)�2�db�u0�@� '4TX�m0�pa3i1A3s0Q25�c��st�r�VR1%e�q0
��j1 ��O2 �A�UEiy�@.�‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?P Q��qA!Pvs� 5	1 5aU���?PŅ���ဝQ9A6�zS*�7�qb5�1����Q��'00P(��V7]u�a itE1���ïp?7� �!?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ�޵y00\ry�"R�2BL�tN  ���� �1DfA>�2�qeR�5���_b�3�X]1m1l�cqP1�a�E�Q� 5�F����!5���@M-16Q�� f���r���Q�e� ��� PN�L�T_�1��i1��945�3��@�e�|�b1l>F1u*AY2�
�R8�Q����RJ�J13�D}T� 85
Qg� /0��*A!P�*A�Ð�d����2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt]1 ^u�ajrI�B����~`�|I�b��yI�\m�Qb�I�uz�A�c3Apa\9q� B6S��S��m���}�85`N�N�  �(M�� �f1���6����161j��5�s`�SC���U��A����5\se�t06c����10��y�h8��a6��6x��9r�2HS �� �Er���W@}�a��IlB���Y�ٖ�m�u �C����5�B��B��h`�F���X0���A :���C�M��AZ��@��4�6i����� e�O�-	���f1��F  �ᱦ�1F�Y	���GT6HL3��U66~`Ȗ��U�dU�9D20Lf0��Qv� ��fjq ��N������0v
� ���i	�	��72l�qQ2������� \�chngmove�.V��d���@2l_arf	�f ~��6������9C��Z���~���kr41@ S���0��V��t�����U�p7nu�qQ%�A]��V�1\"�Qn�BJ�2W� EM!5���)�#:��64��F�e50S �\��0�=�PV�� �e������E������m7shqQSH"U��)��9�!A���(���� �,[>�ॲTR11!��,�60e=��4F�����2��	 R-����������@�Ж��4���LS0R�)"�!lOA��Q�X) %!� 16�
U /��2�"2�E�9p���2>X� SA/i��'�
7F�H�@!B�0�� �D���5V��@2cV E��p��T��pt갖��1L~E�#�F�Q��9�E�#De/��RT��59���	�A�EiR���|����9\m20챃20��+�-u�19r4 �`�E1�=`O9`� �1"ae��O�2��_\$W}am41�4�3��/d1c_std ��1)�!�`_T��r~�_ 4\jdg�a �q�PJ%!~`-�r�+�bgB��#c300D�Y�5j�QpQb1�`bq��vB��v25�Up�����qm43�  �Q<W�"PsA��e ����t�i�P�W .��c�FX.�e4�kE14�44�~o6\j4�443sxj��r�j4up�� �\E19�h�PA�T�= :o�APf��coWol!\�2a��2A;_	2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a�:88J9X�l5�m�1a첚��*���(85�&�������P6���R,52&A����,fA9IfI50\u�z�OV
�v��}E�֖J���Y>� 16�r�C�Y��;��1��L ���Aq�&ŦP1��vB�)e�m�����1pĻ �1Df>�27��F�KAREL �Use S��FC�TN��� J970�FA+�� (�Q޵0�p%�)?�Vj9F?(��j�Rtk208 C"Km�6Q�y�j��iæPr�9�s#��v��krcfp�RCF�t3���Q��kcctme�!ME�g����^6�main�dV�� ��ru��kDº��c���o����J�dt��F �»�.vrT�f�����E%�!��\5�FRj73B�K����UER�HJ�O  �J�� (ڳF���F �q�Y�&T��p�F�z��19�tkvBr���V�Bh�9p�E�y�<�k�������;�v���"CT��f����)�
І ��)�V	�6���!� �qFF��1q���=��� ��O�?�$"���$���je���TCP A�ut�r�<520 �H5�J53E19�3��9��96�!8���9��	 �B574V��52�Je�(�� Se%!Y�����u���ma�Pqtool��ԕ������co�nrel�Ftro�l Reliab�le�RmvCU!��H51����� a�551e"�CNRE¹I�c�&���it�l\sfut?st "UTա��"X�\u��g@�i�D6Q]V0�B,Eѝ6A� �Q�)C���X���Yf�I�1|6s@6i��T6IU��vR��d�
$e%1��2�C58�E6��8�Pv�iV�4OFH58SOeJ� mnvBM6E~O58�I �0�E�#+@�&�F�0 ���F�P6a���)/++��</N)0\tr1x�����P ,[>ɶ��rmaski�ms�k�aA���ky'd�h�	A	�P�sDisp_layIm�`v��~��J887 ("A��+Heůצprd�s��Iϩǅ�h�0p�l�2�R2��:�Gt�@��PRD�TɈ�r��C�@Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��Px^@�P�firmQ� ���Pp�2�=bk�6�r��3��6��tppl��PL���O�p<b�ac�q	��g1J�U�d0�J��gait_9e���Y�&��Q���	�S�hap��erat�ion�0��R6�7451j9(`sGen�ms�42-f�Ár�p�5����2�rsgl�E��p�G���qF�205p�5S���ՁN�retsap�BP�O��\s� "GC�R�ö? �qngda�G��V��st2axU��Aa]��b�ad�_�btpu�tl/�&�e���tp�libB_��=�2.p����5���cird��v�slp��x�hex��v�re?�Ɵx�gkey�v�pm���x�us$�6�gcr��F������[�q27�j92�v�ollismqSk�9O��>�� (pl.���t��p!o��29$Fo8���cg7no@�tptwcls` CLS�o�b�\�km�ai_
�!s>�v�o	�t�b��x�ӿ�E�H��6~�1enu501�[�m��utia|$c�almaUR��Ca�lMateT;R5	1%�i=1]@-��/V�� ��Z�� �fq1�9 "K9E�L����z2m�CLMTq��S#��et �LM�3!} �F�c�ns�pQ�c���c_mo4q��� ��c_e���F��su��ޏ �_ �x@�5�G�join�@i�j��oX���&cW0v	 ���N�ve��C�clm�&Ao# �|$�finde�0�STD ter� FiLANiG���R��
��8n3��z0Cen���r,������J��� �� ���K��Ú�=�К�_Ӛ��r� "FNDR�� 3��}f��tguid��`��N�."��J�tq��  �������������J����_������c���	m�Z��\fndr.��n#>
B2�p��Z�CP Ma�����38A��� c
��6� (���N�B ������� 2�$�	81��m_���"ex�z5�.Ӛ��c���bSа�ef�Q��	��RBT~;�OPTN � +#Q�*$�r*$��*$r *$%/s#C�d/.,P�/|0*ʲDPN���$���$*�Gr�$ko Exc�'IF�$�MASK�%93 {H5�%H558�$_548 H�$4-1��$��#1(�$�0 E�$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3��9j0"M�49�4 � ��4�4tp�sh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E�\���5�A�4��3a�dq\�5K979�":E�ajO l "�DQ^E^�3i�Dq� ��4ҲO ?R�? ��q�5��T��3rAq�O�Lst�5~��7�p�5��REJ#�2�@a�v^Eͱ�F���4��.��5y N� �2il�(in�4��31 aJH1�2Q4�251ݠ��4rmal� �3) �REo�Z_�æOx�����4��^F�?onor Tf��7_ja�UZҒ4l��5rmsAU�Kkg���4�$HCd\�fͲ�e�ڱ�4�REM���4y�ݱ"u@�RER593�2fO��47Z��5lity,�U��e"DGil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe�=$��^�
E��u�IAymptm�U��BU��vste�y\�3��me� b�DvI�[�Qu�:F�U�b�*_�
E,�su$��_ Er��oxx���4huse�E-�?�sn�������FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��� b���(��1�� �c��Y�R�� �>�P� ��W��������'��0ɵ�[��͂����  � ,[N@� �A��bumpšf��B*�Box%��7Aǰ�60�BBw���MC� u(6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`���)���\bbk968� "�4�ω�bb��9va69����etbŠ��X�����#ed	�F��u�f�& �sea"������'�\��,���b�ѽ"�o6�H�
�x�$�f���!y���Q[�!� tperr�f�d� TPl0o� R/ecov,��3D���R642 � 0���C@}s� N@��(NU�rro���yu2�r��  �
�  ����$$�CLe� �������������$~z�_DIGIT��.������ .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ oo$j��+c:PRODUCTM��0\PGSTKD��V&ohozf99���D���$F�EAT_INDE�X��xd���  
�`IL�ECOMP ;����#��`�cS�ETUP2 <��e�b�  �N �a�c_AP2�BCK 1=�i  �)wh0?{%&c����Q� xe%�I�m�� �8��\�n����!� ��ȏW��{��"��� F�Տj���w���/�ğ S���������B�T� �x������=�үa� �����,���P�߯t� �����9�ο�o�� ��(�:�ɿ^���� �ϸ�G���k� �ߡ� 6���Z�l��ϐ�ߴ� ��U���y����D� ��h��ߌ��-���Q� ��������@�R��� v����)�����_��� ��*��N��r� �7��m�@&�3\�i
pP� 2#p*.V1Rc�*��`� /��PC/|1/FR6:/"].��/+T�`�/ �/F%�/�,�`r/?��*.F�8?	�H#&?e<�/�?;STM �2�?�.K �?��=iPen�dant Panel�?;H�?@O�7�.O�?y?�O:GIF �O�O�5�OoO�O_:JPG _J_�56_�O�_�_�	PANE�L1.DT�_@�0�_�_�?O�_2�_�So�WAo�_o�o�Z3 qo�o�W�o�o�o)�Z4�o[�WI���
TPEINSO.XML��0�\���qCust�om Toolb�ar	��PAS�SWORDy�FRS:\L�� �%Passwo�rd Config���֏e�Ϗ�B 0���T�f�������� ��O��s������>� ͟b��[���'���K� �򯁯���:�L�ۯ p�����#�5�ʿY�� }��$ϳ�H�׿l�~� Ϣ�1�����g��ϋ�  ߯���V���z�	�s� ��?���c���
��.� ��R�d��߈���;� M���q������<��� `������%���I��� �����8����n ���!��W�{ "�F�j| �/�Se��/ �/T/�x//�/�/ =/�/a/�/?�/,?�/ P?�/�/�??�?9?�? �?o?O�?(O:O�?^O �?�O�O#O�OGO�OkO }O_�O6_�O/_l_�O �__�_�_U_�_y_o  o�_Do�_ho�_	o�o -o�oQo�o�o�o�o @R�ov��; �_���*��N� �G������7�̏ޏ m����&�8�Ǐ\�� ���!���E�ڟi�ӟ ���4�ßX�j����� ���įS��w�������B�#��$FIL�E_DGBCK �1=��/���� ( ��)
SUMMA�RY.DGL����MD:������Diag Sum�mary��Ϊ
C?ONSLOG������D�ӱCon�sole log�E�ͫ��MEMCHECK:�!ϯ����X�Memory� Data��ѧ��{)��HAD�OW�ϣϵ�J����Shadow C?hangesM�'��-��)	FTAP7Ϥ�3ߨ���Z��mment TB�D��ѧ0=4)�ETHERNET��������T�ӱE�thernet �\�figurat�ionU�ؠ��DCSVRF�߽߫������%�� ve�rify all���'�1PY���DIFF�����[����%��diff]������1R�9�K���� ���X=��CHGD������c��r�����2ZAS� ��GD����k��z��FY�3bI[� �/"GD����s/����/*&UPDATES.� ��/��FRS:\��/�-ԱUpda�tes List��/��PSRBWLOD.CM(?���"�<?�/Y�PS_ROBOWEL��̯�? �?��?&�O-O�?QO �?uOOnO�O:O�O^O �O_�O)_�OM___�O �__�_�_H_�_l_o �_�_7o�_[o�_lo�o  o�oDo�o�ozo�o 3E�oi�o�� �R�v���A� �e�w����*���я `���������O�ޏ s������8�͟\�� ���'���K�]�쟁� ���4���ۯj����� �5�įY��}���� ��B�׿�x�Ϝ�1� ��*�g�����Ϝ��� P���t�	�ߪ�?��� c�u�ߙ�(߽�L߶� �߂���(�M���q�  ���6���Z���� ��%���I���B������2�����h�����$FILE_� P�R� ��������M�DONLY 1=�.�� 
 � ��q��������� �~%�I�m �2��h� �!/�./W/�{/
/ �/�/@/�/d/�/?�/ /?�/S?e?�/�??�? <?�?�?r?O�?+O=O �?aO�?�O�O&O�OJO �O�O�O_�O9_�OF_�o_
VISBCK�L6[*.VD�v_�_.PFR:\��_�^.PVis�ion VD file�_�O4oFo\_ joT_�oo�o�oSo�o wo�oB�of�o �+����� ��+�P��t���� ��9�Ώ]�򏁏��(� ��L�^�������5� ��ܟk� ���$�6�ş�Z��~�����
M�R_GRP 1>�.L��C4 w B���	 W������*u����RHB ���2 ��� ��� ���B� ����Z�l���C���D�ি����Ŀ��K����J�Z�I���T�*�F�?5UP�pE����ֿ E�M.G��E$��;�n߇:G��@�O���@��6�@�O�f���@�T=@�1��*λ� F@ ��������J��N�Jk�H9��Hu��F!��/IP�s�?�����(�9�<9���896C'�6<,6\b��+�&�(�a�L߅�p�A��A��߲�v� ��r������
�C�.� @�y�d�������� ������?�Z�lϖ�;BH�� �Ζ�������
0�PS@�P�J���ܿ�� �B���/ ��@�33:��.�gN��UUU�U��q	>u.�?!r�X��	�-=�[z�=�̽=�V6<�=�=�=$q������@8�i7�G��8�D�8@9!�7��:����D�@ D�� Cϥ�V�C������'/ 0-��P/����/N��/ r��/���/�??;? &?_?J?\?�?�?�?�? �?�?O�?O7O"O[O FOOjO�O�O�O�O�� �ߵ��O$_�OH_3_l_ W_�_{_�_�_�_�_�_ o�_2ooVohoSo�o wo�o�i��o�o�o ��);�o_J�j �������%� �5�[�F��j����� Ǐ���֏�!��E� 0�i�{�B/��f/�/�/ �/���/��/A�\�e� P���t��������ί ��+��O�:�s�^� p�����Ϳ���ܿ�  ��OH��o�
ϓ�~� �Ϣ����������5�  �Y�D�}�hߍ߳ߞ� �������o�1�C�U� y��߉������ ������-��Q�<�u� `��������������� ;&_J\� ���������ڟ �F�j4���� �����!//1/ W/B/{/f/�/�/�/�/ �/�/�/??A?,?e? ,φ?P�q?�?�?�?�? O�?+OOOO:OLO�O pO�O�O�O�O�O�O_ '__K_�o_�_�_�_ l��_0_�_�_�_#o
o Go.okoVoho�o�o�o �o�o�o�oC. gR�v���� �	���<�`�* <��`�����ޏ ��)��M�8�q�\��� ����˟���ڟ��� 7�"�[�F�X���|��� |?֯�?�����3�� W�B�{�f�����ÿ�� �������A�,�e� P�uϛ�b_�����Ϫ_ ��߀�=�(�a�s�Z� ��~߻ߦ��������  �9�$�]�H��l�� �����������#�� G�Y� �B�������z� ������
ԏ:�C. gRd����� �	�?*cN �r�����/ ̯&/�M/�q/\/�/ �/�/�/�/�/�/?�/ 7?"?4?m?X?�?|?�? �?�?�?��O!O3O�� WOiO�?�OxO�O�O�O �O�O_�O/__S_>_ P_�_t_�_�_�_�_�_ �_o+ooOo:oso^o �o�op��o�� �� $��o�o�~ �������5�  �Y�D�}�h������� ׏����
�C�.� /v�<���8������ П����?�*�c�N� ��r��������̯� �)��?9�_�q���JO �����ݿȿ��%� 7��[�F��jϣώ� �ϲ�������!��E� 0�i�T�yߟߊ��߮� �߮o�o��o>� t�>��b�������� ���+��O�:�L��� p������������� 'K6oZ�Z� |�~�����5  YDi�z�� ����/
//U/ @/y/@��/�/�/�/�� �/^/???Q?8?u? \?�?�?�?�?�?�?�? OO;O&O8OqO\O�O �O�O�O�O�O�O_�O�7_��$FNO ����VQ��
F0�fQ kP FLAG�8�(LRRM_C�HKTYP  rWP��^P�WP��{QOM�P_MI�N�P����P��  XNPSSB_CFG ?VU ���_���S ooIUTP�_DEF_OW � ��R&hIR�COM�P8o�$G�ENOVRD_D�O�V�6�flTH�R�V d�edkd_�ENBWo k`R�AVC_GRP s1@�WCa X"_ �o_1U<y �r�����	� �-��=�c�J���n� �������ȏ�����;�"�_�F�X���ibR�OU�`FVX�P��&�<b&�8�?��埘���|����  D?��јs���@@g�B��7�p�)�ԙ���`SMT�cG�mM����| �LQHOSTC�Rs1H���P��a�t�SM��f��\���	127�.0��1��  e��ٿ�����ǿ�@�R�d�vϙ�0�*�	�anonymou�s�����������0Qu[�� � ��� ��r����ߨߺ����� -���&�8�[�I�� �������1� C��W�y���`�r��� ���ߺ�������%� c�u�J\n���� �����M�"4 FX��i���� ��7//0/B/T/ ���m/��/�/ �/??,?�/P?b?t? �?�/�?��?�?�?O Oe/w/�/�/�?�O�/ �O�O�O�O�O=?_$_ 6_H_kOY_�?�_�_�_ �_�_'O9OKO]O__Do �Ohozo�o�o�o�O�o �o�o
?o}_Rd v���_�_oo! �Uo*�<�N�`�r��o ������̏ޏ�?Q�&�8�J�\���>�EN�T 1I�� P�!􏪟  �� ��՟ğ�������A� �M�(�v���^����� 㯦��ʯ+�� �a� $���H���l�Ϳ���� �ƿ'��K��o�2� hϥϔ��ό��ϰ�� �����F�k�.ߏ�R� ��v��ߚ��߾���1����U��y�<�QUICC0��b�t���1�����%���2�&���u�!ROUTERv�R�d���!PCJOG�����!192.�168.0.10���w�NAME �!��!ROBO�Tp�S_CFG� 1H�� ��Auto-started�t/FTP��� ���� 2D ��hz����U ��
//./�v�� �/���/�/�/�/ �/�!?3?E?W?i?�/ ?�?�?�?�?�?�?� ��AO�?eO�/�O�O �O�O�?�O�O__+_ NO�OJ_s_�_�_�_�_ 
OO.OoB_'ovOKo ]ooo�oP_>o�o�o�o �oo�o5GYk }�_�_�_��8o ��1�C�U�$y��� �����ӏf���	�� -�?�����Ə�� �ϟ�����;� M�_�q���.�(���˯ ݯ��P�b�t����� m���������ǿٿ�� ���!�3�E�h��{� �ϟϱ����$�6�H� J�/�~�S�e�w߉ߛ� jϿ��������*߬��=�O�a�s��YT_?ERR J5
�����PDUSIZ � ��^J�����>��WRD ?�t��  ?guest}���%�7�I�[�m�$SC�DMNGRP 2�Kt�������V$�K�� �	P01.14� 8��   �y����B  _  ;������ ���������
 �������������~�����C.gR|����  i  ��  
��������� +��������
����l .r���"B�l��� m
d�������_GROuU��L�� ��	����07EQU�PD  	պ��J�TYa �����TTP_AUT�H 1M�� <�!iPenda�ny��6�Y!�KAREL:*8��
-KC///�A/ VISION SETT�/v/�"�/�/�/#�/ �/
??Q?(?:?�?^?�p>�CTRL �N����5�
�FFF9E3�?��FRS:DE�FAULT�<�FANUC We�b Server�:
�����<kO}O��O�O�O�O��WR_�CONFIG �O�� �?��I�DL_CPU_P5C@�B��7Pw�BHUMIN(\���<TGNR_IO������PNPT_SIM_DOmV�w[TPMODN�TOLmV �]_P�RTY�X7RTOL_NK 1P��� �_o!o3oEoWoio�RMASTElP��R>�O_CFG�o�i�UO��o�bCYC�LE�o�d@_AS�G 1Q����
 ko,>Pbt� ��������\sk�bNUM����<K@�`IPCH�o���`RTRY_CN�@oR��bSCRN(����Q��� �b�`��bR���Տ���$J23_DSP_EN	����?OBPROC�Un�iJOGP1SY�@��8�?��!�T�!�?*�POS�RE�zVKANJI_�`��o_�� ���T�L�6͕����C�L_LGP<�_���EYLOGGIN�`���LANGUAGE YF�7RD w���LeG��U�?⧈�x� �����=P�V�'0��$ N�MC:\RSC�H\00\��LN�_DISP V���
��������OC��R.RDzVTA{�O�GBOOK W�
{��i��ii��X�����ǿٿ���b��"��6	h������e�?�G_B�UFF 1X�]��2	աϸ���� �������!�N�E� W߄�{ߍߺ߱����߀�����J���D�CS Zr� =����^�+�ZE���������a�IO 1[
{ ُ!� �!�1�C�U�i�y��� ������������	 -AQcu�������EfPTM  �d�2/AS ew������ �//+/=/O/a/s/p�/�/��SEV�����TYP��/??y͒�RS�@"��×�FL 1\
������?�?��?�?�?�?�?/?TP�6��">�NG�NAM�ե�U`�UPS��GI}�𑪅}mA_LOAD��G %�%D?F_MOTN���O��@MAXUALRM<��J��@sA�Q�����WS ��@C �]�m�-_���MP2�7�^�
{ ر�	�!P�+ʠ�;_/��Rcr�W�_�WU�W �_��R	o�_o?o"o coNoso�o�o�o�o�o �o�o�o;&Kq \�x����� ��#�I�4�m�P��� |���Ǐ���֏��!� �E�(�i�T�f����� ß��ӟ���� �A� ,�>�w�Z�������ѯ ����د���O�2� s�^�������Ϳ����ܿ�'��BD_LDXDISAX@	��MEMO_APR@�E ?�+
 � *�~ϐϢϴ�����������@ISC ;1_�+ ��I� �T��Q�c�Ϝ߇��� ������w����>�)� b�t�[����{��� �������:���I�[� /������������o� ����6!ZlS� �s���� 2�AS'�w� ���g��.//�R/d/�_MSTR� `�-w%SCD 1am͠L/�/H/ �/�/?�/2??/?h? S?�?w?�?�?�?�?�? 
O�?.OORO=OvOaO �O�O�O�O�O�O�O_ _<_'_L_r_]_�_�_ �_�_�_�_o�_�_8o #o\oGo�oko�o�o�o �o�o�o�o"F1 jUg����� ����B�-�f�Q����u�����ҏh/MK�CFG b�-�㏕"LTARM_���cL��� σQ�N�<�ME�TPUI�ǂ����)NDSP_CM�NTh���|�  d�.��ς�ҟ|ܔ|�POSCF�����PSTOL �1e'�4@�<#�
5�́5�E�S�1� S�U�g�������߯�� ӯ���	�K�-�?����c�u�����|�SIN�G_CHK  ���;�ODAQ,�f���Ç��DEV �	L�	MC:>!�HSIZEh��-���TASK �%6�%$1234?56789 �Ϡ���TRIG 1g.�+ l6�%����ǃ�����8�p�YP�[� ��EM_IN�F 1h3�� `)AT?&FV0E0"ߙ��)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ������H�����A���AI�q�,��|���� ���ߵ����� J���n������W��� ��������"����X ��/����e�� ����0�T;x �=�as��/ �,/c=/b/�/A/ �/�/�/�/��?� ��^?p?#/�?�/�? s?}/�?�?O�?6OHO �/lO?1?C?U?�Oy? �O�O3O _�?D_�OU_�z_a_�_�ONIT�OR��G ?5� �  	EXESC1Ƀ�R2�X3�XE4�X5�X���V7�X8�X9Ƀ�RhBLd �RLd�RLd�RLd
bLd bLd"bLd.bLd:bLdTFbLc2Sh2_h2khU2wh2�h2�h2�hU2�h2�h2�h3Sh�3_h3�R�R_G�RP_SV 1i�n���(����C�?BPP�A4��>%��gY��>r��x�_D�=R^��PL_NA_ME !6��p��!Defau�lt Perso�nality (�from FD)� �RR2eq 1�j)TUX)TX9��q��X dϏ8� J�\�n���������ȏ ڏ����"�4�F�X� j�|������2'�П �����*�<�N�`�r��<��������ү �����,�>�P�b�: �Rdr 1o�y �{\�, �3����� @D� M ��?�����?�<���A'�6�����;�	lʲ	 ��x�J����� �< �"��� �(pK���K ��K=*��J���J���JV���Z��ƌ��rτ́p@j��@T;f����f��ұ]�l��I����������������b��3���´  ��`��>����bϸ�z���Ꜧ���Jm��
� B�H�˱`]���q�	� p��  P�pQ��p��p|  ���g���c�	'� �� ��I� �  �����:�È
�È=G���"�nÿ�	����I  �n @B�cΤ�\��ۤ�!�q�y�o�N���  '�����@2��@����¬��/�C��C�C��@ C�������
�A�W�@�<�P�R�
h�BD�b�A��j�����:��Dz۩���������j��(� �� -���C���'�7������q�Y����� �??�ff ��g|y �����o�:a��
>+�  PƱj�(�����7	���|�?˙���xZ�p<
�6b<߈;����<�ê<�? <�&Jσ��AI�ɳ+���?offf?I�?&��k�@�.��J<?�`�q�.� �˴fɺ�/��5/� ���j/U/�/y/�/�/ �/�/�/?�/0?q��F�?l??�?/�?+)�?�?�E��� E�I�G+� F��?)O�?9O_O`JO�OnO�Of�BL޳B�?_h�.��O�O�� %_�OL_�?m_�?�__�_�_�_�_�
�h�yÎg>��_�Co�_goRodo�o�GA�ds�q�C�o�o�o|����$]�Hq���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?��$�?�K/����
=ç>�����3�W
=�s#�W��e��9������{�����<��(��B�u���=B0�������	L��H�F��G���G���H�U`E����C�+���I�#�I��H�D�F��E���RC�j=��
�I��@H��!H�( E<YD0q�$� �H�3�l�W���{��� �����՟���2�� V�A�z���w�����ԯ ��������R�=� v�a������������ ߿��<�'�`�Kτ� oρϺϥ�������� &��J�\�G߀�kߤ� ���߳�������"�� F�1�j�U��y���� ���������0��T��?�Q����(��ٙ3/E����u�������q3��8�����q4Mgqs&IB+2�D�a���{�^^	�������uP2P7Q 4_A��M0bt��R������/   �/�b/ P/�/t/�/ *a)_3/�/�/�%1a?�/�?;?M?_?q?   �?�/�?�?�?�?O �2 F�$�vGb�/�A��@�a�`�qC��C@�o�Ot����KF� Dz�H@�� F�P �D���O�O�ys�<O!_3_E_W_i_s?_���@@pZ�4�22!2~
 p_�_�_�_ 	oo-o?oQocouo�o��o�o�o��Q ���+��1��$M�SKCFMAP � �5�� �6�Q�Q"~�cONREL  
�q3�bEXC/FENB?w
s1u�XqFNC_QtJO�GOVLIM?wdtIpMrd�bKEY?wu�u�bRUN�|��u�bSFSP�DTY�avJu3sS�IGN?QtT1M�OT�Nq�b_C�E_GRP 1p�5s\r���j� ����T��⏙���� ��<��`��U���M� ��̟��🧟�&�ݟ J��C���7������� گ�������4�V�`�TCOM_CFG 1q}�Vp������
P�_ARC_�\r
jyUAP_�CPL��ntNOCHECK ?{ 	r�� 1�C�U�g�yϋϝϯπ��������	��({N�O_WAIT_L��	uM�NTX�r�{�[m�_ERR�Y�2sy3�  &�������r�c� ��T_MO��t>��, �A$�k�3�PARAM��u{�	�[����u?�� =9@345?678901�� &���E�W�3�c�����`{�������������=�UM_RSPACE �Vv���$ODRDS�P���jxOFFSET_CARTܿαDIS��PE?N_FILE� �q���c֮�OPTIO�N_IO��PW�ORK v_�ms �P(�R�Qp
�j.j	 ��H�j&6$� RG_DSBL  �5�Js�\��RIE�NTTO>p9!CᴧPqfA� UT__SIM_D
r��b� V� LCT ww�bc��U)+$�_PEXE�d&R�ATp �vju�p��2�X�j)TUX)T�X�##X d -�/�/�/??1?C? U?g?y?�?�?�?�?�?��?�?	OO-O?O�H2 �/oO�O�O�O�O�O�O�O�O_]�<^O;_M_ __q_�_�_�_�_�_�_`�_o���X�OU[��o(��(����$o�, ���IpB` @D��  Ua?�[cAa?p]a]�DWcUa쪞�l;�	lmb�`�xJ�`�p���a�<� ��`� ���b��H(��H3�k7HSM5G��22G���Gpc
��
���,'|��CR�>�>q��GsuaT�3���  �4spBpyr�  ]o�*SB_�����j]��t3�q� ��r�na �,���6 W ��PQ�|N�M�,k����	'� � ���I� � � ��%�=�̡ͭ���ba	����I  �n �@��~���p��������N	 W�  �'!o�:q�pC	 C��@@sBq�|��� Nm�
�!�h@ߐE�n����*�B	 ��A���p� �-�qbz��P��t��_������( �� -��@恊�n�ڥ[A]Ѻ�b�4�'!5�(p �?�ff� ��
����!OZ�R*�85�z�:��>΁  Pia��(5���@���ک�a�c��dF#?��5�x���*�<
6b<�߈;܍�<��ê<� <�#&�o&�)�A�lc�ΐI�*�?fff?��?&c���@�.�uJ<?�`��Yђ^�nd��]e ��[g��Gǡd<���� 1��U�@�y�dߝ߯� �����߼�	���-�������&��"�E��� E��G+� Fþ������������&��J�5��bB��AT�8�ђ��0�6� ��>���J�n�7���[m�0��h�y�1��>�M��I
�@��A�[��C-�)<��?����( /�YĒ��Jp���vav`CH/����x��}!@I�Y��'�3A�A�A�R1AO�^??�$�?�����±
=ç>�����3�W
=�#����+e���ܒ�����{�����<��.�(�B�u���=B0�������	�*H��F�G���G���H�U`E����C�+�-I�#�I��H�D�F��E��RC�j=U>�
I��@H��!H�( E?<YD0/�? �?�?�?�?O�?3OO WOBOTO�OxO�O�O�O �O�O�O_/__S_>_ w_b_�_�_�_�_�_�_ �_oo=o(oaoLo�o �o�o�o�o�o�o�o '$]H�l� ������#�� G�2�k�V���z���ŏ ���ԏ���1��U� g�R���v�����ӟ��������-��(��3������a�����Q�c�,!3ǭ8�}���,!4M�gs����ɢIB+�կ篴a���{���A�/�e�S�(��w��P!�P�������7��ӯ����R9�Kτ�oχ�,�ϥ�  ���χ� ���)��M������ z���{߉ߛ������ߤ�������  )�G�q�_����~��2 F�$�&'Gb���n�[Z,jM!C�s�@j/��A�S�=�F� D�z��� F�P D��W����)�����������x�?���@@
J9�=�=��=��
 v� �������*<N`�*P ����˨�1��$�PARAM_ME�NU ?-���  �DEFPULS�El	WAIT�TMOUT�R�CV� SH�ELL_WRK.�$CUR_STY�L�,OPT��/PTB./("C��R_DECSN ���,y/�/�/�/�/ �/�/?	??-?V?Q?�c?u?�?�USE_PROG %�q%�?�?�3CCR������7_HOSoT !�!�44O�:T̰�?PCO)A�RC�O�;_TIMqE�XB�  �?GDEBUGV@���3GINP_FL'MSK�O�IT`��O��EPGAP �L̳�#[CH�O�HTY+PE����?�? �_�_�_�_�_oo'o 9obo]ooo�o�o�o�o �o�o�o�o:5G Y�}����������1�Z��EW�ORD ?	7]�	RS`�	P�NS�$��JO�E!>�TEs@WVT�RACECTL �1x-�� �����Ɇ_DT Qy-��~�D � ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�T�(�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_j��_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ�_��� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��������//"#��$PGTRACE�LEN  #! � ���" �8&_UP _z���g!o �S!h 8!_CFoG {g%Q#�"!x!�$J �#|"D�EFSPD |��,!!J �8 I�N TRL }ʇ-" 8�%�!PE�_CONFI� ~>g%�g!�$��%�$LID�#��-74GRP 1��7Q!�#!A ���&ff"!�A+33D�� �D]� CÀ SA@+6�!�" d�$�9�9*1*0� 	� +9�(�&�"�? #´	C�?�;B@3A�O�?OIO3OmO"!>�T?�
5�O��O�N�O =��=#�
�O_�O_ J_5_n_Y_�O}_�_y_x�_�_�_  Dzco" 
oBo�_Roxo co�o�o�o�o�o�o �o>)bM��;�
V7.10b�eta1�$ � A�E�r�ϻ�A " �p?!{G��q>���r���0�q�ͻqB7Q��qA\�p�q��4�q�p�"�B�@�2�D�V�h�w��p�?�?)2{ȏw� ׏���4��1�j�U� ��y�����֟���� ��0��T�?�x�c��� ����ү����!o�,� ۯP�;�M���q����� ο���ݿ�(��L��7�p�+9��sF@ �ɣͷϥ�g%��� ���+�!6I�[߆��� ���ߵߠ��������� !��E�0�B�{�f�� ������������ A�,�e�P���t����� �������=( aL^����� ��'9$]�� ���ϖ������� /<�5/`�r߄ߖߏ/ >�/�/�/�/�/?�/ 1??U?@?R?�?v?�? �?�?�?�?�?O-OO QO<OuO`O�O�O�O�O ���O_�O)__M_8_ q_\_n_�_�_�_�_�_ �_o�_7oIot�� �o�o���o�o�o(/ !L/^/p/�/{*o� �������� A�,�e�P�b������� ���Ώ��+�=�(� a�L���p������Oߟ 񟠟� �9�$�]�H� ��l�~�����ۯƯ�� �#�No`oro�on��o �o�o�oԿ���8 J\ng����vϯ� ��������	���-�� Q�<�u�`�r߫ߖ��� ��������;�M�8� q�\��������z��� ���%��I�4�m�X� ��|����������� :�L�^���Z������ �����$�6�H� Swb��� ����//=/(/ a/L/�/p/�/�/�/�/ �/?�/'??K?]?H? �?��?�?f?�?�?�? O�?5O OYODO}OhO �O�O�O�O�O�O&8 J4_F_����_�_ ��_�_"4-o�O *ocoNo�oro�o�o�o �o�o�o)M8 q\������ ���7�"�[�m��? ����R�Ǐ���֏� !��E�0�i�T���x� �������_$_V_ ��2�l_~_�_�����R��$PLID_KNOW_M  �T?������SV ��U.͠�U��
� �.�ǟR�=�O������mӣM_GRP S1��!`0u��T�@ٰo�ҵ�
 ���Pзj��`��� !�J�_�W�i�{ύϟπ����������߱�MR�����T��s�w� s��ߠ޴߯߅� �ߩ߻�����A��� '��������� ������=���#��� ������}������S��{ST��1 1��U�# ���0�_ A .��,>Pb �������� 3(iL^p������2�*���<-/3 /)/;/M/4f/x/�/�/5�/�/�/�/�6??(?:?7 S?e?w?�?8�?�?��?�?MAD  �d#`PARNUM  qw�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a�OT>_CMP_��B@��P@'˥TER�_CHK'U��0˪?R$_6[RSl�¯���_MOA@�_�U_��_RE_RES_G ��>�oo8o +o\oOo�oso�o�o�o �o�o�o�o�W �\�_%�Ue Baf �S� ����S0� ���SR0��#��S �0>�]�b��S�0}���<���RV 1�����^rB@c]��t�_(@c\����_D@c[�$���RTHR_INRl��DA��˥d,�MASmS9� ZM�MN8��k�MON_QUEUE ���˦��Vx� RDNPUbQqN{�P[��END���_ڙEXE�ڕ�@�BE�ʟ��OPT�IOǗ�[��PROGRAM %���%��ۏ�O��TA�SK_IAD0�OCFG ���tO��^ŠDATA���Ϋ@��27�>�P� b�t���,�����ɿۿ������#�5�G���IWNFOUӌ���� ���ϭϿ�������� �+�=�O�a�s߅ߗ� �߻��������^�jč�� yġ?PDIT �ίc���WERFL
��
�RGADJ �&n�A����?�����@���IORITY�{�QV���MPDSQPH�����Uz��ޝ�OTOEy�1��R� (!AF�4�E�P]���!�tcph���!�ud��!icqm��ݏ6�XY_ȡ��R��ۡ)�� *+/ ۠� W:F�j�� ����%7�[B�*��POSRT#�BC۠�����_CARTR�EP
�R� SKS�TAz��ZSSAV����n�	2500H863���r�T$!�R���Áq�n�}/�/�'� U�RGE�B��rYW�F� DO{�rUVW�V��$�A�WRUP�_DELAY ��R��$R_HOT�k��%O]?�$R_?NORMALk�L?<�?p6SEMI?�?|�?3AQSKIP!��n�l#x 	 1/+O+ OROdOvO9H n��O�G�O�O�O�O�O _�O_D_V_h_._�_ z_�_�_�_�_�_
o�_ .o@oRoovodo�o�o �o�o�o�o�o*< Lr`���n��$RCVTM�v����pDCR!��LЈqB���C*J�C$��>�$ >5?�-;��04M¹��O��ǃ���?����~��9O�n�Y�<
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E/� ATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960/�W+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�M�A�%aR  ��ϰ�P{_��P_INTVAL��@����JR_OPoTION�V �E�BpVAT_GR�P 2�����(y_Ho � e_vo�o�oYo�o�o�o �o�o*<�bOo NDpw����� �	���?�Q�c�u� ����/���ϏᏣ��� �)�;���_�q����� ����O�ɟ���՟ 7�I�[�m�/������� ǯٯ믁��!�3��� C�i�{���O���ÿտ ���ϡ�/�A�S�e� 'ωϛϭ�oρ����� ��+�=���a�s߅� Gߕ߻����ߡ��� '�9�K�]��߁��� ��y����������5��G�Y��E�$SCAN_TIM�AYue�w�R �(ӿ#((�<0.a�aPaP
Tq>��Q��oa�����OOE2/��:	d/"JaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>7��̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:��_O�UT",REC 1�Z� d w   	�    �� @������A�����
 ��PSD#6 rT��O� �� �� �`�� �Z�{�� �� *�  �+X- � I- �*- !- � �X��YZ�PSJ;4� �?  (�  � ���R ��� E*- � �/e/��l4�/��� X� (,/>/P/��/�/�""4� =T�!� � ؀  ?�"S1��'!�/���("- ��\?�? $=�=�?�?�?"OOFO 4OjO|O^O�O�O�O�O �O�O�O_ __T_B_ x_f_�_�_�_�_�_�_ �_oooPo>oto�o ho�o�o�o�o�o�o (
L:\�p���w,��� �4�"�X�F�|���p� ����֏ď����0� �@�f�T���x����� ҟ�Ɵ���,��<� b�P���h�z������ ί��(�:��^�L� n�p�������ܿ�п � �6�$�Z�H�jϐ� rϴϢ���������� 2�D�&�h�Vߌ�z߰� ������������
�@��.�d�R��ZjV 1�w P�����j 
�� ���
TYPE�VFZN_CF�G ��5�d�4�GRP �1�A�c ,B� A� D;� �B���  B4~RB21/HELL:�(
���?���<%RS'!��H3l W�{�������2Vh������%w����#!�1���S��7�2�0d�|���HK 1��� �k/f/x/�/ �/�/�/�/�/�/?? C?>?P?b?�?�?�?�?~��OMM �����?��FTOV_E�NB ���+�HOW_REG_UIO~��IMWAITB��JKOUT;Fܻ�LITIM;E����OVAL[OMC_�UNITC�F+�M�ON_ALIAS� ?e�9 ( he��_&_8_J_\_ B_�_�_�_�_j_�_ �_oo+o�_Ooaoso �o�oBo�o�o�o�o �o'9K]n� ���t���#� 5��Y�k�}�����L� ŏ׏������1�C� U�g����������ӟ ~���	��-�?��c� u�������V�ϯ�� ����;�M�_�q�� ������˿ݿ���� %�7�I���m�ϑϣ� ��`�������ߺ�3� E�W�i�{�&ߟ߱��� ���ߒ���/�A�S� ��w����X���� ������=�O�a�s� ��0������������� '9K]�� ��b���# �GYk}�:� �����/1/C/ U/ /f/�/�/�/�/l/ �/�/	??-?�/Q?c? u?�?�?D?�?�?�?�? O�?)O;OMO_O
O�O �O�O�O�OvO�O__�%_7_�C�$SMO�N_DEFPRO ���`Q� *�SYSTEM* � d=OUREC�ALL ?}`Y� ( �}4xc�opy fr:\�*.* virt�:\tmpbac�k�Q=>192.�168.4�P46?:7924 �R�_X�_�_�K}5�Ua�_��_�V�_goyo�o}
�xyzrate 61 +o=oOo�o�o�e�g�n6580 �o�ocu�b�9�Ts:orde�rfil.dat��l*<q���l0�Rmdb:�o�<q �b�t���c6��x�emp:�1652� W������.��*.d��ƎϏ`�r����o1 +�=�O���� �)Ғ��ҟc�u� ����5�͇ٯ��� �"���̈ѯb�t��� c�_�o?�U����
� o����=�׿h�z�� ����:�տ����
�� ��A���d�v߈ߛ�.� ;�ѿ�����Ϫ߼� O�`�r��ϩ�2��� ������'���K�\� n����ߥ�8������� ���#��G�j| ���o3EW���<��W5012?� bt����4�5� ���"��5�b/�t/�/������P8188 W/�/�/�/� �/�)�/`?r?�?��� ;?M?�?�?O'�4 �?�?cOuO�O��5/ �'�O�O�O/"/�O�) �Oc_u_�_����RB U_�_�_
o�_�_TA �_hozoo�O�O:_�_ �o�o
_�oA_�od v��_.o;�_�� �o��Oo`�r��� �o�o2�oޏ����'K\�n�������$SNPX_AS�G 1�������� P� 0 '%�R[1]@1.1,����?���%֟� �&�	��\�?�f��� u��������ϯ��"� �F�)�;�|�_����� ��ֿ��˿���B� %�f�I�[Ϝ�Ϧ��� ��������,��6�b� E߆�i�{߼ߟ����� ������L�/�V�� e���������� ��6��+�l�O�v��� ������������2 V9K�o�� �����&R 5vYk���� �/��<//F/r/ U/�/y/�/�/�/�/? �/&?	??\???f?�? u?�?�?�?�?�?�?"O OFO)O;O|O_O�O�O �O�O�O�O_�O_B_ %_f_I_[_�__�_�_ �_�_�_�_,oo6obo Eo�oio{o�o�o�o�o �o�oL/V� e������� �6��+�l�O�v��������PARAM ������ W�	��P�����OFT_KB_CFG  ������PIN_SI/M  ���C��U�g�����RVQS�TP_DSB,��򂣟����SR ��/�� &  �AR�����TOP_ON_ERސ����PTN� /�@��A	�RING_�PRM� ��V�DT_GRP 1y�ˉ�  	�� ����������Я��� ��*�Q�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߣߠ߲��� ��������0�B�i� f�x���������� ���/�,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZ�~��� ����/ /G/D/ V/h/z/�/�/�/�/�/ �/?
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8___\_��VPRG_COUNT���@���RENB�U��UM�S��__U�PD 1�/�8  
s_�oo*o SoNo`oro�o�o�o�o �o�o�o+&8J sn������ ���"�K�F�X�j� ��������ۏ֏��� #��0�B�k�f�x��� ������ҟ������ C�>�P�b����������ӯί�����UY?SDEBUG�P�P��)�d�YH�SP_�PASS�UB?~Z�LOG ��U+�S)�#�0��  ��Q)�
M�C:\��6���_M�PC���U���Q�ñ8� �Q�SAV �����ǲ%��ηSV;�TE�M_TIME 1]��[ (�P�T�y�ؿT1SVGgUNS�P�U'�U����ASK_OPTION�P�U�Q�Q���BCCFG 3��[u� n�X�G�`a�gZo��߃� ���߹�������:� %�^�p�[����� ���� �����6�!�Z� E�~�i���������%�������&8�� nY�}�?��� � ��(L: p^������ �/ /6/$/F/l/Z/ �/~/�/�/�/�/�/�/ �/2?8 F?X?v?�? �??�?�?�?�?�?O *O<O
O`ONO�OrO�O �O�O�O�O_�O&__ J_8_n_\_~_�_�_�_ �_�_�_o�_ o"o4o joXo�oD?�o�o�o�o �oxo.TBx ��j����� ���,�b�P���t� ����Ώ��ޏ��(� �L�:�p�^������� ʟ��o��6�H� Z�؟~�l�������د ���ʯ ��D�2�h� V�x�z���¿���Կ 
���.��>�d�Rψ� vϬϚ��Ͼ������� *��N��f�xߖߨ� ��8���������8� J�\�*��n����� ��������"��F�4� j�X���|��������� ����0@BT �x�d���� �>,Ntb� �����/�(/ /8/:/L/�/p/�/�/ �/�/�/�/�/$??H? 6?l?Z?�?~?�?�?�? �?�?O�&O8OVOhO zO�?�O�O�O�O�O�O 
__�O@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<o^o�oro�o �o�o�o�o�o  J8n$O���� �X���4�"�X��B�v��$TBCS�G_GRP 2��B�� � �v� 
 ?�  ������׏�� �����1��U�g�z����ƈ�d, ����?v�	 HC{��d�>����~e�CL  B����Пܘ������\)��Y  A��ܟ$�B�g�B�Bl��i�X�ɼ���X��  D	J���r������C����үܬ���D�@v�=�W�j�}� H�Z���ſ���������v�	V�3.00��	mw61c�	*X�0P�u�g�p�>���v�(:�� ��p͟�w  O����p������z�JCFG [�B��� ���������=��=�c�q�K�q� �߂߻ߦ�������� '��$�]�H��l�� �����������#�� G�2�k�V���z����� ���������p* <N���l��� ����#5GY }h����v� b��>�// /V/D/ z/h/�/�/�/�/�/�/ �/?
?@?.?d?R?t? v?�?�?�?�?�?O�? *OO:O`ONO�OrO�O �O��O�O�O_&__ J_8_n_\_�_�_�_�_ �_�_�_�_�_oFo4o jo|o�o�oZo�o�o�o �o�o�oB0fT �x������ �,��P�>�`�b�t� ����Ώ������� &�L��Od�v���2��� ��ȟʟܟ� �6�$� Z�l�~���N�����د Ư�� �2��B�h� V���z�����Կ¿� ���.��R�@�v�d� �ψϪ��Ͼ������ �<�*�L�N�`ߖ߄� �ߨ����ߚ����� ��\�J��n���� �������"���2�X� F�|�j����������� ����.TBx f������� >,bP�t �����/�(/ /8/:/L/�/�ߚ/�/ �/h/�/�/�/$??H? 6?l?Z?�?�?�?�?�? �?�?O�?ODOVOhO "O4O�O�O�O�O�O�O 
_�O_@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<oro`o�o�o �o�o�o�o�o&�/ >P�/���� �����4�F�X� �(���|�����֏� ���Ə0��@�B�T� ��x�����ҟ����� �,��P�>�t�b��� ������������ :�(�^�L�n������� 2d�����̿�$� Z�H�~�lϢϐ����� ���Ϻ� ��0�2�D� zߌߞ߰�j������� ���
�,�.�@�v�d� ������������ �<�*�`�N���r��� ����������& J\�t��B� �����F4 j|��^���8�/�  2 6#� 6&J/6"�$�TBJOP_GR�P 2����  ?��X,i#�p,� ��xJ� �6$�  �<� �� �6$� @2 �"	 ��C�� �&b  �Cق'�!�!>��1�
559>�0+1��33=�C�L� fff?+0?�ffB� J1�%Y?�d7�.��/>���2\)?0�5����;��hCY�� �  @� �!B�  A�P?�?�3~EC�  D�!8�,�0*BOߦ?�3�JB��
:���Bl�0��0�$�1�?�O6!Aə�A�̔C�1D�G6�=qq�E6O0�p��B��Q�;�A}�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH�1�ts�A@33@?1� C�� �@�_x�_&_8_>��D�U�V_0�LP�Q30<{�zR� @�0�V�P !o3o�_<oRifoPo^o �o�o�oRo�o�o�o�o M(�ol�p~(��p4�6&�q5	V3.00�#�m61c�$*�(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I�R�CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;S@;Q��|8�`rz@/&�8�6&<��1�w�^$�ESTPARS c *({ _#HR��ABLE 1�p+IZ�6#|�Q� � 1�|�|�|�5'=!*|�	|�
|�|�˕�6!|�|�|�N��RDI��z!ʟ@ܟ� ��$���O�������¯ԯ�����S��x# V���˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� U-����ĜP�9�K�]� o��-�?�Q�c�u���~6�NUM  ��z!� >  �Ȑ����_CFG ������!@b IMEBF_TT��p��x#��a�VER���b�w�a�R 1Ξp+
 (3�6"1 ��  6!������ ���� �9�$�:�H�Z� l�~����������������^$��_��@�x�
b MI_CH�ANm� x� kDOBGLV;0o�x��a!n ETHERA�D ?�� ��y�$"�\&n R�OUT��!p*!�*�SNMA�SK�x#�25�5.h�fx^$O�OLOFS_DI�[ՠ	ORQC?TRL �p+;/ ���/+/=/O/a/ s/�/�/�/�/�/��/��/�/!?��PE_D�ETAI��PON_SVOFF��33P_MON ��H�v�2-9STRTCHK ����42VTCOM�PATa8�24:0FPROG %��%CA)&O�3I�SPLAY��L:_�INST_MP 2GL7YDUS���?��2LCK�LPKQUICKMEt �O�2oSCRE�@�
tps��2�A�@�I��@_Y���9��	SR_GRP �1�� ���\�l_zZg_�_�_�_�_�_�^�^�oj �Q'ODo/ohoSe��o o�o�o�o�o�o�o !WE{i�������	1234567��!�ڎ�X�E1�V[
 ��}ipnl/�a�gen.htm�no��������ȏ~��Panel s/etup̌}�?�`�0�B�T�f� �� 񏞟��ԟ���o� ���@�R�d�v����� �#�Я�����*� ��ϯůr��������� ̿C��g��&�8�J� \�n�����϶����� ����uϣϙ�F�X�j� |ߎߠ����;��������0�B��*NUA�LRMb@G ?�� [������ ������ ��%�C�I��z�m�������v�SEoV  �����t�ECFG �Ё=]/BaA$  w B�/D
 �� /C�Wi{��� ���� PRց; �To\o�eI�6?K0(%�� ��0�����/ /;/&/L/q/\/�/�/�/l�D �Q�/�I_�@HIST �1ׁ9  (�  ��(/S�OFTPART/�GENLINK?�current=�menupage?,153,1?v?8�?�?�?�� >?P=962c?�?
OO.O�?�?�136�?|O�O �O�OAOSOeO�O__ 0_�HM___q_�_�_�_ �_H_�_�_oo%o7o �_[omoo�o�o�oDo �o�o�o!3E ��a81�ou��� ���o���)�;� M��q���������ˏ Z�l���%�7�I�[� ��������ǟٟh� ���!�3�E�W���� ������ïկ�v�� �/�A�S�e�Pb�� ����ѿ������+� =�O�a�s�ϗϩϻ� ������ߒ�'�9�K� ]�o߁�ߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y��� v�����������	 �?Qcu��( ����)� M_q���6� ��//%/�I/[/ m//�/�/�/D/�/�/ �/?!?3?�/W?i?{? �?�?�?�����?�?O O/OAOD?eOwO�O�O �O�ONO`O�O__+_ =_O_�Os_�_�_�_�_ �_\_�_oo'o9oKo �_�_�o�o�o�o�o�o jo�o#5GY�o�}������?���$UI_PAN�EDATA 1������  	�}��0�B�T�f�x��� ) ����mt�ۏ���� #�5���Y�@�}���v� ����ן�������1���U�g�N������ �1��Ïȯگ� ���"�u�F���X�|� ������Ŀֿ=���� ��0�T�;�x�_Ϝ� �ϕ��Ϲ������,���M��j�o߁ߓ� �߷������`��#� 5�G�Y�k��ߏ��� �����������C� *�g�y�`��������� F�X�	-?Qc ����߫���� ~;"_F� �|�����/ �7/I/0/m/�����/ �/�/�/�/�/P/!?3? �W?i?{?�?�?�?? �?�?�?O�?/OOSO eOLO�OpO�O�O�O�O �O_z/�/J?O_a_s_ �_�_�_�O�_@?�_o o'o9oKo�_oo�oho �o�o�o�o�o�o�o# 
GY@}d�� &_8_����1�C� �g��_��������ӏ ���^���?�&�c� u�\�������ϟ��� ڟ�)��M����� ������˯ݯ0��� ��7�I�[�m������ ����ٿ�ҿ���3� E�,�i�Pύϟφ���0����Z�l�}���1� C�U�g�yߋ�)߰� #������� ��$�6� ��Z�A�~�e�w��� ��������2��V��h�O�����v�p��$�UI_PANEL�INK 1�v��  ��  ��}12�34567890 ����	-?G � ��o�����a ��#5G�	�����p&���   R�����Z� �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?.O@O ROdOvO�O O�O�O�O �O�O_�O�O<_N_`_0r_�_�_�0,���_ �X�_�_�_ o2ooVo hoKo�ooo�o�o�o�o �o�o��,>r} ��������� ���/�A�S�e�w� �������я���t v�z����=�O�a� s�������0S��ӟ� ��	��-���Q�c�u� ������:�ϯ��� �)���M�_�q����� ����H�ݿ���%� 7�ƿ[�m�ϑϣϵ� D��������!�3�E� �_i�{�
�߂����� �������/��S�e� H���~��R~'�'� a��:�L�^�p��� ������������  ��6HZl~�� �#�5��� 2 D��hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?�/ �?�?�?�?�?�?m?O O&O8OJO\O�?�O�O �O�O�O�O�O[�_�� 4_F_)_j_|___�_�_ �_�_�_�_o�_0oo Tofo��o��o��o �o�o,>1b t����K�� ��(�:����{O ������ʏ܏�uO� $�6�H�Z�l������� ��Ɵ؟����� �2� D�V�h�z�	�����¯ ԯ������.�@�R� d�v��������п� ��ϕ�*�<�N�`�r� ���O�Ϻ�Io������ ���8�J�-�n߀�c� �߇����߽����o 1�oX��o|���� ���������0�B� T�f������������ ��S�e�w�,>Pb t��'���� �:L^p� �#���� // $/�H/Z/l/~/�/�/ 1/�/�/�/�/? ?�/ D?V?h?z?�?�?�??? �?�?�?
OO.O��RO dO�߈OkO�O�O�O�O �O�O_�O<_N_1_r_ �_g_�_7OM�m��$UI_QUI�CKMEN  >��_Ao�bRESTORE� 1�?  �|��Rto�o�im�o�o�o�o �o:L^p� %������o� ���Z�l�~����� E�Ə؏���� �Ï D�V�h�z���7����� ��/���
��.�@�� d�v�������O�Я� ����ßͯ7�I��� m�������̿޿��� �&�8�J��nπϒ� �϶�a�������Y�"� 4�F�X�j�ߎߠ߲� �����ߋ���0�B�T�gSCRE`?�#mu1s]co`u2��3��U4��5��6��7��y8��bUSERq�dv��Tp���ks����4��5��6��7���8��`NDO_�CFG �#k � n` `PDA�TE ����NonebSE�UFRAME  ��TA�n�RTO?L_ABRTy�l�Α�ENB����GR�P 1�ci/aCz  A�����Q@�� $6HR�d��`U�����MSK  �����MNv�%�U�%����bVISCAN�D_MAX�I���FAIL_�IMG� �PݗP#���IMREGN�UM�
,[SI�Z�n`�A�,~VONTMOU��@���2���a��a��~��FR:\� � MC{:\�\LOG�7B@F� !�'/�!+/O/�Uz �MCV�8#U�D1r&EX{+�S|�PPO64_���0'fn6PO��LIb�*�#9V���,f@�'�/�� =	�(SZV��.����'WAI��/STAT 	����P@/�?�?�:�$�?�?��2DW�P  ��P yG@+b=��� H��O_JMPE�RR 1�#k
 � �2345678901dF�ψO{O �O�O�O�O�O_�O*_�_N_A_S_�_
� M�LOWc>
 �_�TI�=�'M�PHASE  ���F��PSHI[FT�1 9�]@<�\�Do�U#oIo �oYoko�o�o�o�o�o �o�o6lCU �y����� �@�	�V�-�e2����	VSFT1�2�	VM�� ��5�1G� ���%A_�  B8̀̀E�@ pكӁ˂�у���z�ME@�?��{��!c>&%�aM�1��k�0�{ �$�`0TDINEND��\�O� �z���S��w��P��=�ϜRELE�Q���Y���\�_ACT�IV��:�R�A ���e���e�:�R�D� ���YBOX� �9�د�6���02���1�90.0.�83v��254�:�QF�	 �X��j��1�ro�bot���  � p�૿�5pc��̿������7�����-�f�ZABC�����,]@U��2 ʿ�eϢωϛϭϿ� ���� ���V�=�zߐa�s߰�E�Z��1� Ѧ