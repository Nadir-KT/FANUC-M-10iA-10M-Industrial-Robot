��   9�A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT�
&F/�d $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STPS_L�OG_P N��$��T�N�  �6 COUNT_D�OWN�$EN�B_PCMPWD� � DV�I�N!$C� C{RE�PARM:z� T:DIAG:�)�LVCHK|!FULLM0�YXT�CNTyD�MENU!�AUTO,��$$CL(   O������	���	�VIRTUA�� ��$DCS_7COD@������  W'_S+  *�! T&��A91&"!=. 
 $��� ~-�/�/�/�/�/�/�/ ??0?>?T?b?x?�?��?�?�?��`#SUP�� l+�?�?`#F��?OFO�� C sLpA���O z ��� V�[t�&��j�� mB@O�O��G�O��XU 