��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �
  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"'�ASB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�:�OFF_ N�3D;ELHLOGn25Aa2?i1@N�?�� -M�H W�+0�$Y $DB\� 6COMW!2�MO� 21\D.	� \rVE�1$qF��A{$O���D�B�CTMP1_5F�E2�G1_�3�B��2GXD�#�
 d $CA�RD_EXIST�4$FSSB_�TYPuAHKBgD_S�B�1AGN �Gn $SL?OT_NUMJQoPREV,DBU� �g1G ;1_EDIT�1 � 1G�=� S�0%$�EP�$OP��AETE_�OKRUS�P_CRQ$;4�V� ^0LACIw1`�RAPk �1x@ME@$D�V�Q�P�v�A{oQL� OUzR ,mA�0��!� B� LM_O��^eR�"CAM_�;1 xr$ATTR4NP� �ANN�@5IMG?_HEIGHQ�c�WIDTH4VT�� �UU0F_ASwPECQ$M�0gEXP��@AX�f��CFT X O$GR� � S�!z�@B@NFLI�`<t� UIRE 3dT�uGITCHC�`N�� S�d_L�`�C��"�`EDlpE� J�4S�0� �zsa4 hq�;G0 � 
?$WARNM�0f�!,P� �s�pNST�� CORN�"a1F�LTR�uTRAT�� T�p H0AC�Ca1���{�OcRI
`"S={RT0�_S�B�qHG,I.1 [ Tp�"3I9�TY�D,P*
2 �`w@� �!R*HD�cJ* C��U2��3��4��5��U6��7��8��94u�qO�$ <� �$6xK3 1w`O_�M�@�C t 2� E#6NGP�ABA� �c��ZQ���`���@nr��� ��aP�0����x�p�PzPb26����"MJ�_R��BC�1J��3�JVP���tBS��}Aw��"�tP�_*0OFSzR @� RO_K8���a�IT�3��NOM_��0�1ĥ3�ACPT �� $���2AxP��K}EX�� ��0g0I01��p�
$�TFa��C$MD3&��TO�3�0U� ��/ �Hw2�C%1|�EΡg0wE{`vF�vF�40CPp@��a2 
P$A`PqU�3N)#��dR*�AX�!sDET;AI�3BUFV��p@1 |�p۶�pkPIdT� PP[�EMZ�Mg�Ͱj�F[�SIMQSI�"0��A.���:�kx T�p|zM��P�B�F�ACTrbHPEW�7�P1Ӡ��v��MC�d� �$*1JqB�p<�*1DECH����H��(�c� �� +PNS_EMP��$GP���,P!_��3�p�@Pܤ��TC��|r��0�s�� b�0�� �B���!
����JR� ��SEGF�R��Iv �aR�TrkpN&S,�PVF4|��� &k� Bv�u�cu��aE�� !2���+�MQ��E�SIZ�3����T��P���|��aRSINF� ����kq���������LX�����F�CRCMu�3CClpG�� p���O}���b�1����P���2�V�DxIC��C���r����P��{�� EV �zF_J��F�pNB0�?�������A�! � r�Rx����V�lp�2���aR�t�,�g�R>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!��$SK��2��P� �"�"@�P�R8� 
 �D8���# >�q1�$��$��E�L9$?(�V�y%@?�Ai�PC9&_?R4ENE��c'~?(�� RE�p�Y2(H �O�S��#$L�3$$@3R��;3�MVOks_D@!V�ROScr�r�w�S���CRIG7GER2FPA�S��>7�ETURN0B�c�MR_��TUː\[��0EWM%���cGN>`��RLA���Eݡ�P�&$�P�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWA�YRMO#�aw!��DCS_)7  `IS#�  �� �s3S�AQ汯 4Rx�ZSW�AQ�p�@r1UW��cTNTV)�5RV
a���|c�éW�ƃ��JB��x0��S�AFEۥ�V_SV>�bEXCLUU�;���ONL��cY�g�~az�OT�a{�HI_V? ��R, M��_ *�0� ��_�z�2� CdSGO  +�rƐm@��A�c~b���w@��V��i�b�fANNUNXx0�$�dIDY�UABc�@Sp�i�a+ �j��f�"�pOGIx2,���$F�b�$ѐO�T�@A $DUMMY��Ft��Ft�±� 6U- ` !�HE�|s���~bc�B@ SUFFmI��4PCA��Gs5Cw6Cq����DMSWU.{ 8!�KEYI��5�TM�1�s�qoA�v�INޱE��!, /{ D��HOST�P!4���<���<�°<��p<�EM'���Z�n� SBL� UL��0  �	�����DT�01 ϴ $��9USAMPLо�/����ĺ�$ I@갯 $SUBӄ��w0QS��8���#��SAV������c�S< 9�`�fP�$�0E!� YN_�B�#2 0�`DI��d�pO|�m��#$�F�R_IC� �?ENC2_Sd�3  ��< 3�9����� cgp����4��"��2�A��ޖ5���`ǻ�@Q@�K&D-!�a�AVE�R�q����DSP
���PC_�q��"�x|�ܣ�VALU3��HE�(�M�IP\)���OPPm �CTH�*��S" $T�/�Fb�;�d�����d D�.'��ET�6 H(rLL_DUǀ�a�@��k����֠OT�"U�/���o�@@NOAUT5O70�$}�x�~�@s��|�C� ���C� 2iaz�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|�pw�����9 <���z�ΓKI����H猡�BaFEq@{@:� ,��&a? �P_P?��>�����E�@��iaQQ���;fp$TP�$VARI����,�7UP2Q`< W�߃TD��g���`�������!��BAC�"=# T2����$)�,+r8³�p IFI��p�� q M�P"�l@|``>t ;��46����ST����T��M ����0	 ��i���F����������kRt ����FORC�EUP�b܂FLUS
pH(N��� ��^6bD_CM�@E��7N� (�v�P��REM� Fa��@Pj���
K�	N����EFF/���@I�N�QOV��O{VA�	TROV� DT)��DTMX:e �P:/��P`q�vXpCLN A_�p��@ ��	_|�F�_T: �|�&P%A�QDI���`1��0�Y0RQ"m�_+qH���M���sCL�d#�RIV{��ϓN"EAR/�IOF�PCP��BR���CM�@N 1b �3GCLF��!DaY�(��a�#5T�CDG���� �%,��FSS� )�? PP(q1�1�`_1�"811�EC13zD;5D6�GRA�J��@�����PW��ON2EBUG��S�2�C`gϐ_E� A ��?�q��TERM�5�B�5$Z �OR�Iw�0C�5.TP��SM_-`���0DV�5���0A�9E�5�LD1�UP��F�� -QϒA��P�3�@B$SEG�GJ� EL�UUSE.PNFI��pBx���1@��4>DC$UF�P��$���Q�@"C���G�0T������SNSTj�PATxۡg��APTHJ�A�E*�Z%qB\`F�{E��F�q�pARxPY�aSHFT͢qA�AX_SHOR$�>��6% @$GqPE���GOVR���aZPI@P�@$U?r *aAYLO���j�I�"��A8ؠ��ؠERV��Q i�[Y)��G�@R��i�e��i�R�!P�uA�SYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C��%UP���P���WORڒ@M��k0SM5T��G��GR��3�aPA�@��p5�'�_H � j�A�'TOCjA7pP]Pp$OPd�O��C��%�p�O!��R%E.pR�C�AO�?��Be5pR�EruIx|'QG�e$PWR) �IMdu�RR_$s �PT�b�B I�z2H8�=�_ADD�RH�H_LENG��B�q�q:�x�R��S�o�J.�SS��SK������� ��-�S�E*����HSN�M-N1K	�j�5�@r�֣OL��\�WpxW�Q�>pACRO�p ���@H ����Q� N��OUPW3�b_>�I��!q�a1����� ���|��������`-���:���iIOX2S=�D�e��]���L $��p�!_�OFF[r_�PRM�_��aTTPu_�H��M (�p�OBJ�"�pG�$�H�LE�C��ٰN� � 9�*�AB%_�T��
�S�`�S6��LV��KRW"du�HITCOU?B-Gi�LO�q�����d� Fpk�GpSS� ���HWh�wA���O.��`INCP}UX2VISIO�� !��¢.�á<�á-¿ �IOLN)�P� 87�R'�[p$�SL�bd PUTM_��$dp�Pz x�� F_AS2Q/�$LD���D�DaQT U�0]P�A������PHYG灱Z�̵�5�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp���x�X�ٶ%�UJ��S��v��NE�WJOG�GN �DIS��&�KĠL��3T |��AV���`_�CTR!S^�FgLAGf2&�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_H��Dq��N?���V��EE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�B�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S Sxn��I�BUFF1�XY��PT�$��� �v��f���װA
�rYY��P ������pOS1�2�3�K�0Z � � ��aiE�*��IKDX�dP�RhrO�X+��A&ST��R���Yz�<! Y$EK&CK+���Z&m&pFp�5�0[ L�� o�0��]PL�6pwq�t�^����t�7�_ \ �`��瀰�7�t�#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3�1DM�R7��LDR5<4R5ORG.���e2(` ���V�8.��T<�4�d^ �q�<4��-4R5�S�`T00m��0D>FRCLMC!D�?0�?3I@��MIC��dg_ d���RQm�=q�DSTB	� c �Fg�HAX;b� �H�LEXCE�SZrBPqCMup�a`Z��B;d�oE`��`5a��F_A�J���$[�O�H0K�db q\��ӂS�$MB���LIБ}SREQU�IR�R>q�\Á�XD�EBU��oAL� MP�c�ba��P؃ӂ!B�oAND���`�`d0�҆�c�cDC1��IN�����`@�(h?�Nz�@q��o��UP�ST8� e�rL�OC�RI�p�E�X�fA�p��AoAOwDAQP�f X��3ON��[rMF���� �f)�"I��%�e��T�vQFX�@IGG� g �q��"E��0��#���$R�a% ;#7y��Gx��VvCPi�ODATAw�pE:��y��RFЭ�NVh �t $MD�qI�ё)�v+�tń�tH��`�P�u�|��sAN�SW}��t�?�uD��)�b�	@Ði -�@CU��V�T0�eRR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2N�RIN��v�<��'NTE���kE����,��b����_Nl@��ڂ��kDׄRm�7DIViFDH�@ـ:n�$V��'cv!$��$Z������~�[��o�H �$BEL�Tb��!ACCEL�+��ҡ��IRC��t����T/!���$PS�@#2L�@ q�Ɣ83������� ��PATH��������3̒Vp�A_�Q�.��4�B�Cᐈ�_M=Gh�$DDQ���G�$FWh��p���m�����b�DE��P�PABNԗROTSPEED����00�J�Я8��@���@�$USE_��P���s�SY��c�A �>qYNu@Ag��OsFF�q�MOUN�3NGg�K�OL�H�INC*��a��q��Bxj�L@�BENCS���q�Bđ���D��IN�#"I̒��4�\BݠV�EO�w�Ͳ23_UyPE�߳LOWLA���00����D��@�Bp��� �1RCʀ�ƶMOSIV�JRM�O���@GPERC7H  �OV�� ^��i�<!�ZD<!�c@��d@�P��V1�#P͑��L���EW�ĆĸUP������T�RKr�"AYLOA�!�� Q-�̒<�1�8�`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H�����b�DUM2(�S_�BCKLSH_C ̒��>�=�q�#�U��������2�t�]ACLA�LvŲ�1n�P�C�HK00'%SD�RT�Y4�k��y�1�q_�6#2�_UM$Pj�C�w�_�SCL��ƠLMT_J1_LO�"�@���q��E������๕�幘SPC`��7������PCo�B��H� �PU�m�C/@��"XT_�c�CN_b��N��e���SFu���V�&#����9�̒d��=�C�u�SH6# ��c����1�Ѩ�o�0�0͑
��_�PAt�h�_Ps�W�_10��4֠R�01D�VG�J� L��@J�OGW���ToORQU��ON*ɀMٙ�sRHљ��_	W��-�_=��C��TI��I�I�II�	F�`�JLA.�1[��VC��0�D�BO1�U�@i�B\JRK�U��	@DBL_�SMd�BM%`_D9LC�BGRV��0C��I��H_� �*COS+\�(LN�7+X>$C�9)�I�9)u*c,)�Z2 HƺMY@!�( "�TH&-�)THET=0�NK23I��"l=�A CB6CB=�C�A�B(261C�61�6SBC�T25GT	S QơC��aS$�" �4c#�7r#$DUD�EX�1s�t��B�6䆱�AQ|r�f$NE�DpIB U�\B5��	$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2��&�C�J�&!�VAHV�6H3�YLVhJVuKV��KV�KV�KV�KV�IHAHZF`RXM��wX�uKH�KH�KH�KH��KH�IO2LOAHOT�YWNOhJOuKO�KUO�KO�KO�KO�&�F�2#1ic%�d4GS�PBALANCE�_�!�cLEk0H_�%SP��T&�bc&�b>r&PFULC�hr��grr%Ċ1ky�U�TO_?�jT1T2Cy��2N&�v�ϰ ctw�g�p�0Ӓ~����T��O���� IN�SEGv�!�REV8�v!���DIF�鉳1l�w�1m
�OaB�q
����MIϰ�1��LCHWAR̭���AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|�n��ROBR�CR�����N�'�MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD���ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDX�Р  ��MOR^��t $-�U�� )��r�B���������Gؒu � $SIMULT ��~�x�� ���OBJE�`> �ADJUS>�1�OAY_Ik��D_�����C�_FIF�=�T� ��Ұ��{���p� �����p�@��DN�FRI��ӥT�ՓRO� ��E����͐OPWO�ŀv�0��SYSBU<�@ʐ$SOP�����#�U"��pPRUYN�I�PA�DH��D����_OU��=��qn�$}�IMKAG��ˀ�0P�q3IM����IN�q�~��RGOVRDȡ:���|�P~���Р�0�L_6p���i��R)B������M���SEDѐF� ��N`�M*�����̰SL��`ŀw x $�OVSL�vSDI��DEXm�g�e�9Hw�����V� ~�N����w����Ûǖȳ�M��͐�q<��� �x HˁE�F�AWTUS���C�08àǒ��BTM����If���4����(�.ŀy DˀEz�g���PE�r�����
���EXE��V��E�pY�$Ժ ŀz @ˁf��UP{�h�$�p��XN���9�H�� �PG"�{ h $SUB���c�@_��01\�MP�WAI��P����L�O��-�F�p�$�RCVFAIL_9C�-�BWD"�F����DEFSPup | Lˀ`�D��8� U�UNI���S���R`���_L��pP��̐���ā} ��� B�~���|��`Ҳ�N�`KET��y�R��P� $�~���0SIZE�ଠ{����S<�OR��FORMAT/p � F�,��rEMR��y�cUX���LI7�~ā  $�P_SWI���@��_PL7�AL_� �ސR�A��B��(0C��Df�$mEh����C_=��U� � � 1���~�J3�0��^��TIA4��5��6��MOM������� �B�AD`��*��* PU70�NRW��W �R����� A$PI�6���	�� )�4l�}69��Q�|��c�SPEED�PGq�7�D�>D�� ���>tMt[��SAM�`痰>��MOV���$�@�p�5��5�D�1�$2�������{�2��Hip�IN?,{� �F(b+=$�H*�(_$<�+�+GAMM�f�1>{�$GET��Đ�H�D����
^pLI�BR�ѝI��$H�I��_��Ȑ*B6Eď�*8A$>G086LW =e6\<G9�686��R���ٰV��$�PDCK�Q�H�_����;"��z�.%��7�4*�9� ��$IM_SR�O�D�s"���H�"�L	E�O�0\H��6@Á��U� �ŀ��P�qUR_SCR�ӚAZ��S_SA�VE_D�E��NO��CgA�Ҷ��@�$ ����I��	�I� %Z [� ��RX" ��m� ��"�q�'"�8 �Hӱt�W�UpS�*��R�M��O㵐 .'}q��Cg���@ʣȳߑ��BM�AÂ� ?� $PY��g$WH`'�NGp� ��H`��Fb��Fb��Fb��PLM���	� 0h�H�{�X��O��z�Zp�eT�M���� pS��C��O__0_�B_�a��_%�� | S����@	�v��v  �@���w�v��EM��%(O�fr�B�ː��ft�P��PM��QU.� �U�Q��A�-�QTH=�HOLޫ�QHYS�ES��,�UE��B��O.#��  -�P0�|��gAQ���ʠu���O��ŀ�ɂv�-�A;ӎ�ROG��a2�D�E�Âv�_�ĀZ�INFO&��+�����bȜ�OI킍 =((@SLEQ/��#������o���DS`c0O�0�01�EZ0NUe�_�AUyT�Ab�COPY�P�Ѓ�{��@M��N������1�P�
� ��RiGI�����X_�P�l�$�����`�W��P��j@�G���EXT_CYCtb!���p����h�7_NA�!$�\��<�RO�`]�� � m��PORp�ㅣ���SRVt��)����DI �T_ l���Ѥ{�ۧ��ۧ Ъۧ5٩6٩7٩8����AS�B쐒���$�F6���PL8�A�A^�TAR��@ E `�Z�����<��d7� ,(@FLq`hѦ�@YNL���M�C���PWRЍ��=�e�DELAѰ��Y�pAD#q��Q�SKIP�� Ĵ��x�O�`NT!� ��P_x���ǚ@ �b�p1�1�1Ǹ� ?� �?��>��>�&��>�3�>�9�J2�R;쐖 4��EX� TQ����ށ�Q����[�KFд��@R;DCIf� �U`�X}�R�#%M!*�0��)��$RGEAR_�0IO�TJBFLG��igpERa��TC�݃������2TH2yN��� 1�b���Gq T�0 �$���M���`Ib�����REF�1��� l�h��ENAB��lcTPE?@��� !(ᭀ����Q�#�@~�+2 H�W���2������"�4�F�X���
��3�қ{����(����j�4�Ҝ��
���.�@�R�j�5�ҝ�u�����������j�6�Ҟ��(:L
j�7�ҟo���(��j�8�Ҡ���"4Fj�SMS�K�����a��E��A��MOTE������@ "1�L�Q�IO�5"%I���P�ARd�Wi@쐣  �����X�gpi��쐤��Y"$DSB_SIGN4A�Qi��̰C�ШP��S23�2%�Sb�iDEVICEUS#�R�R�PARIT�!O�PBIT�Q��O?WCONTR��QXⱓ�RCU� M�S�UXTASK�3NxB��0�$TATU�P#�#@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�U�PDl�ARB^�� P|%0���� !m$USA���az9�L�ERI�0f��p�RY�5~"_�@f�P8�1�!�6WRK���D9�F9ХFRIgEND�Q4bUF���&�A@TOOLHFM�Y5�$LENG�TH_VT��FI!R�pqC�@�E� IOUFIN�R����RGI�1�AIT�I:�xGX��I�FG2�7G1a����3�B��GPRR�DA��O_0� o0e�I1RER�đ�3&���TC���AQ�JV �G|�.2���F��1�!d�9Z�8+5�K�+5��E�y�L0�4�OX �0m�LN�T�3Hz��89��%�4J�3G��W�0�W�RdD�Z��Tܳ��K��a3d��$cV C2���1��I1H��02K2sk3K3 Jci�aI�i�a�L���SL��R$Vؠ�BVB�EVk�]V*R��� �,6Lc���9V2F{X/P:B��PS_�E���$rr�C�ѳ$A0��wPR���v�Ub�cSk�� {���2��� 0���VX`�!�tX`��0P��Ё�
�!�1SK!� �-qR��!0�i��z�NJ AX�!�h�A�@LlA��A�THIC�1��������1TFE���q>�IOF_CH�3A�I0�����G1�x����豉9�Ɇ_JF�҇PR(���RV{AT�� �-p0��7@����DO�E���COU(��AXI|g��OFFSE+�TRIG�SK��c�� �Ѽ�e�[�K�Hk���8�IGMAo0�A-���ҙ�ORG_U�NEV��� �S��쐮d �$�������GROU���ݓTO2��!ݓD;SP��JOG'��#&	�_P'�2OR�㵸�>P6KEPl�I�R�0�PM�RQ�A	P�Q��E�0q�e����SYSG��"��PG��BRK*Rd�r�3��-�������ߒ<pA�D�ݓJ�BSOC�� N�DUMMgY14�pN@SV�P�DE_OP3SFSPD_OVR���ٰCO��"�OR$-��N�0.�Fr�.�6�OV�SFc�2�f��F��!4�S��|RA�"LCHDL�RECOV��0��W�@M�յ�RO�3��_�0� �@�ҹ@VERE�o$OFS�@CV� 0BWDG�ѴC��2,j�
�TR�!���E_FDOj�MB�_CM��U�B �BAL=r0�w�=q�tVfQ ��x0sp��_�Gxǋ�AM��k�J0�����σ_M��2{�#�8�$CA�{Й���8�$HBK|1c��I�O��.�:!aPPA"�N�3�^�F���:"~�DVC_DB�C���d�w"����!��1ȯ��ç�3����AT�IO� �q0�U8C�&CAB�B�S�PⳍP�Ȗ��_�0c�SUBCPUq��S�Pa aá�}0��Sb��c��r"ơ$HW_C���:c���IcA�A-�l$UNkIT��l��ATN�xf����CYCLų�NECA��[�FLTR_2_FI��0�(��}&��LP&���ނ�_SCT@SF_´�F����G���FS8|!�¹�CHAA/�p���2��RSD�`x"ѡb�r�: _T���PRO��O�� EM��_��8u�qc u�q��DI�0~e�RAILAC��}RMƐLOԠdC���:anq��wq����P�R��SLQ�pfC�ѷ 	��FUNCŢ�rRINkP+a�0� ��!RA� >R �
Я�ԯWAR�BLFQ��aA�����DA��0���LDm0��aB9��nqBT�Ivrbؑ���PRIYAQ1�"AFS�P�! �����`%b����M�I1U�DF_�j@��y1°LME�F=A�@HRDY�4��Pn@RS@Q�0"�MULSEj@f�b�q �X��ȑm���$.A$�1�$c1Ó���o� x~�EGvpݓ�q!AR�����09LB�%��AX]E��ROB��W�A24�_�-֣SY���!46��&S�'WR���-91���STR��t5�9�E�� 	5B��=QB90�@6��������0X1?0�A�RY8�w20���	�%�FI��;�$LGINK�H��1�aI_63�5�q�2XYZ"��;�q�3@�R�1�2�8{0B�{D��� CFI��6G��
�{��_J��6��3aO�P_O4Y;5�QT�BmA"�BC
�z�D�U"�66CTURN3�vr�E�1�9���GFL�`���~ �@��5<:7�� 1��?0K�Mc�68�Cb�vrb�4�ORQ ��X�>8�#op�������wq�Uf�����TOVE�Q��M;�E# �UK#�UQ"�VW�ZQ �W���Tυ� ;��� �QH�!`�ҽ��U�Q�W`keK#kecXER�
�	GE	0��S�dAWaǢ:D���7!�!AX�rB!{q ��1uy-!y�p z�@z�@z6Pz\P z� z1v�y� y�+y�;y�Ky� [y�ky�{y��y�qޜyDEBU��$ ����L�!º2WG` � AB!�,��SV���� 
w���m� ��w����1���1���A ���A��6Q��\Q���!��m@��2CLAB�3B�U�����S 7� ÐER����� � $�@� A6ؑ!p�PO���Z�q0w�_�_MR}Aȑ� d  9T�-�ERR��æ�TYz�B�I�V83@�cΑTOQ�d:`L� �d2ᕴP��˰�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	V FZN_C;FG_!� 4��?� ��|�ų����@�ȲW� �&����\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(�����!�s�Q�g�P{RV H�ELLĥ� }56�B_BAS!�GRSR��ԣo �#QS��[��1r�%��U2ݺ3ݺ4ݺ5ݺ�6ݺ7ݺ8ݷ��R�OOI䰝0�0NL�K!�CAB� ��A[CK��IN��T:��1�@�@ z�m�_P�U!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KcARӑ�@��RE~���P��(�QUE������P
��CST?OPI_AL������0&���㰑�0SE�Ml�b�|�M��d�T�Y|�SOK�}�DI������(���_T}M\�MANRQ���0E+�|�$KEYSWITCH&�	���HE
�BE�AT��cE� LE(Ғ���U��FO���|��O_HOM��O�REF�PPR�z��!&0��C+�OA�ECO��B�rIOCM�D8׵�����8�` � �D�1����U��&�M�H�»P�CFORC���� ��OM>�  � @V��*|�U,3P� 1-�`ʀ 3-�4��NP�X_ASǢ� 0�ȰADD����$�SIZ��$VA�Rݷ TIP]�\�2�A򻡐��Ȑ]�_� �"S꣩!C<ΐ��FRIF⢞�aS�"�c���NF���T�S��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7s��VP�U�PD��  ���|�԰��YSLO>Ǣ� � z��� ����o�E��`>�^t���АALUץ����C�U���wFOqID_YL�ӿuHI�zI�?$FILE_���tf��$`�JvSA���� h���E_B�LCK�#�C,�D_CPU<�{�<�o�����tJr��R ;��
PW O�[ ��LA��S��8������RUNF�Ɂ ��Ɂ����F�ꁡ�ꁾ���TBCu�C�� �X -$�LENi��v������I��G�LOWo_AXI�F1�
�t2X�M����D�
 ���I�� ��}�T#OR����Dh��� L=��⇒�s���#�_MA`�ޕ���ޑTCV����T ���&��ݡ����J�$����J����Mo����J�Ǜ �������2��� v�����F�JK��VKi�ΡvњΡ3��J0�ңJ�JڣJJ�AAL�ң�ڣ��4�5z�&�N1-�9����J��L~�_Vj�ϱ����� ` �GGROU�pD��B�NFLIC��R�EQUIREa�E�BUA��p����2�¯�����c��� \��APPR���C���
�EN��CLOe��S_!M v�,ɣ�
���o� ��MC�8&���g�_MG�q��C� �{�9���|�B;RKz�NOL��|�:� R��_LI|���$��k�J����P
��� ڣ�����&���/���6��6��8��q���� ��8�%��W�2�e�PATH a�z�p�z�=�vӥ�ϰm�x�CN=�CA������p�IN�UCh��bq��CO�UM��!YZ������qE%����2������PAYL�OA��J2L3pR'_AN��<�L��F��B�6�R�{�R_F2�LSHR��|�LO�G��р��ӎ���ACRL_u�������.�r��H�p�$H{�^��FLEX
��}J�� :� /����6�2�����;�M�_�F16����n�@��������ȟ��Eҟ �����,�>�P�b� ��d�{�������������5�T��X ��v���EťmF ѯ�������&��/�A�S�e�&	�x�� � ������j��4pAT����n�EL�  �%øJ���vʰJE��CTR�і��TN��F&��H�AND_VB[�
�pK�� $Fa2{�6� �rSW	��D�U��� $$	Mt�h�R��08��@<b 35��^6A�p3�kƈ�q{9t�A�̈p��A���A�ˆ0��U���D*��D��P��G��ICST��$A��$AN��DYˀ�{�g4�5D� ��v�6�v��5缧�^�@��P����ՠ#�,�5�>�D�J�� &0�_�ER!V9��SQASYM��] ������x��ݑ���_SHl�������sT�( ����(�:�JA����S�cir��_VI��#Oh9�``V_UCNI��td�~�J�� �b�E�b��d��d�f ��n���������uNI����D��H��f����"CqEN� &a�DI��>�Obt2�Dpx�� ��2IxQA����q��-��s� �� s����� �^�OMME�h�rr�QTVpPT�P  ���qe�i����P��x ��yT�Pj� �$DUMMY9��$PS_��R�Fq�0$:� �s���!~q� XX����K�STs�ʰ�SBR��M21_�Vt�8$SV_E�Rt�O��z���CLRx�A  O�r?p? �Oր � D ?$GLOB���#LO��Յ$�o���P�!SYSADqR�!?p�pTCHM0 � ,����oW_NA��/��e�os�TSR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T>D�XSCRE�ƀ5�� ��STF���#}�pТ6�1] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��t<qUE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$1VSHIF��|s�P�p�6��s���R���OSU�RW�pRADIz��2�_�q�h�g!� �q)�LUza�$OUTPUT_3BM��IML�oRp6(`)�@TIL<'SCO�@Ce�; ��9��F��T��a ��o�>�3�����w�2u�<qV�zu✫�%�DJU��|#_�WAIT������%ONE���YBOư ��� $@p%�C�S�Bn)TPE��NE�C��x"�$t$���*B_T��R��%�qRH� ���sB�%�tM�+ Z�t�.�F�R!݀���OPm�MAS�_�DOG�OaT	�D�����C3S�	�O2DE�LAY���e2JO ��n8E��Ss4'#J�aP`6%�����Y_��O2� �2���5��`?� �&�Z�ABCS��  �$�2��J�
 � �$$CLAS>�����A��x@'@@VIRT��O.@ABS�$�1� <E� < *A tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R��d�v�����M@[�AX�Lր�&A�dC  ����IN��ā��P#RE������LARMRECO�V <I䂥�N�G�� \K	 �A   J�\�M@PoPLIC�?<E��E�Ha�ndlingTo�ol �� 
V�7.50P/28~[�  ��o���
�_SW�� �UP*A� ��F�0ڑ����A@��� 20��*A��:���X{�FB 7DA�5�� '@ωo@����No�ne������ ���T�*A4_ynxl�_���V����g�UT�OB�ค����HGAPON8@��LA�ѽU��D 1<EfA����������� Q 1שI Ԁ��Ԑ�:��i�n����#B�)B ���\��HE�Z�r�HTTHKY��$BI�[�m� ����	�c�-�?�Q� o�uχϙϫϽ����� ���_�)�;�M�k�q� �ߕߧ߹�������� [�%�7�I�g�m��� �����������W�!� 3�E�c�i�{������� ��������S/A _ew����� ��O+=[a s������� K//'/9/W/]/o/�/ �/�/�/�/�/�/G?? #?5?S?Y?k?}?�?�? �?�?�?�?COOO1O OOUOgOyO�O�O�O�O �O�O?_	__-_K_Q_���(�TO4�s���DO_CLEAN��|e��SNM  9� �9oKo]ooo��o�DSPDRY�R�_%�HI��m@ &o�o�o#5GY k}����"����p�Ն �ǣ�qX�Մ��ߢ��g�PLU�GGҠ�Wߣ��PRUC�`B`9��o��=�OB��oe�SEGF��K������o %o����#�5�m���LAP�oݎ������ ����џ�����+��=�O�a���TOTA�L�.���USENUʀ׫ �X���R�(�RG_STRI�NG 1��
��M��Sc��
��_ITEM1 �  nc��.�@� R�d�v���������п �����*�<�N�`��r�I/O S�IGNAL���Tryout M�ode�Inp���Simulat{ed�Out��OVERR�`� = 100�In cycl����Prog A�bor�����S�tatus�	H�eartbeat���MH FauylB�K�AlerU� ��s߅ߗߩ߻�����8���� �S�� �Q��f�x���� ����������,�>��P�b�t�������,�WOR������V��
 .@Rdv�� �����*8<N`PO��6� ���o����� //'/9/K/]/o/�/ �/�/�/�/�/�/�/�DEV�*0�?Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO��O�O�OPALT B��A���O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:o�OGRI�p��ra�OLo �o�o�o�o�o�o *<N`r��� ���`o��RB�� �o�>�P�b�t����� ����Ώ�����(��:�L�^�p����PREG�N��.������ ��*�<�N�`�r��� ������̯ޯ����&����$ARG_���D ?	����i�� � 	$��	+[}�]}���Ǟ��\�SBN_CON?FIG i��������CII_SAVE  ���۱Ҳ\�TCEL�LSETUP �i�%HOME�_IO�͈�%M�OV_�2�8�RE�P���V�UTOB�ACK
�ƽFRA:\��� �Ϩ���'`�!��������� ����$�6�c�Z�8lߙ��Ĉ������ �������!凞��M� _�q����2����� ����%�7���[�m� �������@�������`!3E$���J�o�������I�NI�@��ε~��MESSAG�����q��ODE_!D$���O,0.ޜ�PAUS�!�~i� ((Ol� ������� / �//$/Z/H/~/l/�/�'akTSK � q�����UP3DT%�d0;�WSM_CF°�i�еU�'1GRgP 2h�93 |��B��A�/S�XSC�RD+11
1; 	����/�?�?�?  OO$O��߳?lO~O �O�O�O�O1O�OUO_  _2_D_V_h_�O	_X�>��GROUN0O��SUP_NAL��h�	�ĠV_ED�� 11;
 �%�-BCKEDT�-�_`�!oEo%����a��o����,�ߨ���e2no_��o�o�b���ee�o"�o�oED3�o��o ~[�5GED4�n#�� ~�j���ED5Z��Ǐ�6� ~���}���ED6����k�ڏ ~G���!�3�ED7��Z���~� ~�V�şןEDa8F�&o��Ů}p����i�{�ED9���W�Ư
}3�����CRo�����3��տ@ϯ����P�PNO�_DEL�_�RGE?_UNUSE�_�T�LAL_OUT �q�c�QWD_ABOR� �΢Q��ITR_RTN�=���NONSe����CAM_PARAM 1�U�3
 8
SO�NY XC-56� 2345678�90�H � �@���?���(O АV�|[r�u�~�X�HR5k�p|U�Q�߿�R57�����Aff��K�OWA SC31�0M|[r�̀�d @6�|V�� _�Xϸ���V��� ����$�6��Z�l��CE�_RIA_I8j57�F�1��tR|]��_LIO4YW=� ��P<~��F<�GP 1�,���_GYk�*C*  ��CU1� 9� @� G� Z�CLC]� d� l� s�R� ��U[�m� v� � }�� �� C�� ő"�|W��7�HEӰONFI� ��<�G_PRI 1�+P�m®/���������'CHK�PAUS�  1E� ,�>/P/:/ t/^/�/�/�/�/�/�/ �/?(??L?6?\?�?"O�����H�1�_MOR�� =�XaBiq-���5 	 �9 O�?$O@OHOZK�2	���=$9"�Q?55��C�P)K�D3P������a�-4�O__|Z
�OG_�7�PO��� ��6_��,xV�AD�B���='�)
m�c:cpmidb�g�_`��S:�)�����Yp�_)o�S`	�BBi�P�_mo8j�)�Koo�o9i+�)��og�o�o
�m�of�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`)ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCPU�eB�_B�y�;��>C����CnSZE@E�?{hD]^Dْ?r�����D��^��G	���F��F���Cm	fF�O��F�ΫSY����vqG���Em�J)�.���1)��<�Lq�G�x2��Ң ��� a�D�j���E��e��X�EQ��EJP F�E��F� G����F^F E��� FB� H,�- Ge��H3�Y���  >�?33 ���xV�  n2xQ@��5�Y��8B� A�AST<7#�
� �_'��%��wRSMOFSb���~2�yT1�0�DE �O c
��(�;�"�  (<�6�z�R���?��j�C4��SZm� �W��{�m�C��B�-G�C�`@$�q���T{�FPROG� %i����c�I���� �Ɯ�f�KEY?_TBL  �vM��u� �	
��� !"#$%�&'()*+,-�./01c�:;<=>?@ABC�p�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������p��������������������������������������������������������������!j�L�CK��.�j���ST�AT���_AUT/O_DO���W/��INDT_ENB�߿2R��9�+�T2<w�XSTOP\߿2�TRLl�LETE�����_SCRE�EN i�kcsc��U��MMENU 1 i?  <g\�� L�SU+�U��p3g�� ����������2�	� �A�z�Q�c������� ��������.d ;M�q���� ��N%7] �m���/� �/J/!/3/�/W/i/ �/�/�/�/�/�/�/4? ??j?A?S?y?�?�? �?�?�?�?O�?O-O fO=OOO�OsO�O�O�O �O�O_�O_P_Sy�_MANUAL���n�DBCOU�RI�G���DBNUM��p��<���
�QP�XWORK 1!R�ү�_oO.o@o|Rk�Q_AWAY�S���GCP ��=��df_AL�P�dbB�RY�������X_�p� 1"�� , 
�^���o xvJf`MT�I^�rl@��:sONTIM��M����Zv�i
õ��cMOTNEND����dRECORD 1(R�a��ua�O��q��sb� .�@�R��xZ������ �ɏۏ폄���#��� G���k�}�����<�ş 4��X���1�C��� g�֟��������ӯ� T�	�x�-���Q�c�u� ���������>��� �)Ϙ�Mϼ�F�࿕� �Ϲ���:�������%� s`Pn&�]�o��ϓ�~� ����8�J�����5�  ��k����ߡ��J� ����X��|��C�U� ���������0������	��dbTOLEoRENCqdBȺb�`L�͐PCS_?CFG )�k)wdMC:\O �L%04d.CS�V
�`c�)sA V�CH� z�`�)~���hMRC_�OUT *�[��nSGN +��e�r��#�10�-MAY-20 �10:37*V15o-JANj51�k P/Vt��)~�`pa��m��PJP���VERSIO�N SV�2.0.8.|EF�LOGIC 1,^�[ 	DX�P�7)�PF."PROG�_ENB�o�rj U�LSew �T�"_?WRSTJNEp�V��r`dEMO_OPT_SL ?	�e�s
 	R575)s7)�/??*?�<?'�$TO  ��-��?&V_@pE�X�Wd�u�3PA�TH ASA�\�?�?O/{ICTZ�aFo`-�gd>segM%&A�STBF_TTS��x�Y^C��SqqF��PMAU� t/XrMKSWR.�i�a.|S/�Z!D_N�O 0__T_C_x_g_�_�t�SBL_FAUL�"0�[3wTDIAbU 16M�ap�A�123456�7890gFP ?BoTofoxo�o�o�o �o�o�o�o,>�Pb�S�pP�_ ���_s�� 0`� ����)�;�M�_� q���������ˏݏ�|)UMP�!� �^�TR�B�#+��=�PMEfEI�Y_�TEMP9 È��3@�3A v�UNI��.(YN_BRK� 2Y)EMG?DI_STA�%W�ЕNC2_SCR 3��1o"�4� F�X�fv���������#��ޑ14���@�)�;�����ݤ5�����x�f	u� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/߭P�b� t�� ��xߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N���r��� ������������ &8J\n��� �����"`� FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/4?,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O?�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�O�O�o �o�o
.@Rd v������� ��*�<�N�`�r��� �o����̏ޏ���� &�8�J�\�n����������ȟڟ����H�E�TMODE 16v��� ���ƨ
R�d�v�נR�ROR_PROG7 %A�%�:߽��  ��TABLE  A�������#�L�RRSEV_?NUM  ��Q���K�S���_�AUTO_ENB�  ��I�Ϥ_N�Oh� 7A�{��R�  *����J��������^�+��pĿֿ迄�HISO����I�}�_ALM �18A� �;�����+�e�wωϐ�ϭϿ��_H���  A���|��4��TCP_VER �!A�!����$E�XTLOG_RE�Q��{�V�SI�Z_�Q�TOL  ���Dz��A= Q�_BWD���иr���n�_DI�� 9��}�z���<m���STEP����|4��OP_DO����ѠFACTO�RY_TUN�d�G�EATURE �:����l��Handlin�gTool �� � - CEn�glish Di�ctionary���ORDEA�A Vis�� M�aster���9�6 H��nalo�g I/O���H�551��uto �Software� Update � ��J��mati�c Backup~��Part&��ground E�dit��  8\�apCame�ra��F��t\j�6R�ell���LwOADR�omm���shq��TI" ��co��
! yo���pane��� 
!��ty�le selec]t��H59��nD�~��onitor��48����tr��R�eliab���a�dinDiagnos"����2��2 ual Che�ck Safet�y UIF lg�\a��hance�d Rob Se�rv q ct\���lUser F�rU��DIF��E�xt. DIO 6��fiA d��wendr Err YL@��IF�r�ನ  �П�90��F�CTN Menu�Z v'��74� T�P In��fac�  SU (�G=�p��k E�xcn g�3��High-Sper wSki+�  sO��H9 � mmuni]c!�onsg�te�ur� ����V��y��conn���2��EN��Inc=rstru����5.fdKA�REL Cmd.� L?uaA� O~�Run-Ti� 'Env����K� ��u+%�s#�S/W���74��Licen�seT�  (A�u* ogBook�(Sy��m)��"�
MACR�Os,V/Off�se��ap��MH�� ����pfa5�M�echStop �Prot��� d��b i�Shif����j545�!x�r ��#��,�}�b ode Swiwtch��m\e�!�o4.�& pr�o�4��g��M?ulti-T7G����net.P{os Regi���z�P��t Fu9n���3 Rz1���Numx �����9�m�1�  Adju<j��1 J7�7�*� ����6tatu�q1EIKRD�Mtot��scove�� ��@By<- }uest1�$G�o� � U5\SNPX b"���<YA�"Libr��㈶�#�� �$~@h�p�d]0�Jts i?n VCCM����ĕ0�  �u!��2 �R�0�/I�08~��TMILIB�M� J92�@P�A�cc>�F�97�TgPTX�+�BRSQselZ0�M8 Rm��q%��692��Unexceptr �motnT  CcVV�P���KC�����+-��~K  I�I)�VSP CSXC�&.c�� e�"��� t�@We�w�AD Q�8bv9r nmen�@�KiP� a0y�0��pfGridAplay !� nh�@*��3R�1M-10iA�(B201 �`2�V"  F���sci�i�load��8�3 M��l����G�uar�d J85��0�mP'�L`���s�tuaPat�&]$C�yc���|0ori�_ x%Data'Pqu���ch�1���g`� j� RLJa�m�5���IMI �De-B(\A�cP"� #^0C  e�tkc^0assw�o%q�)650�Ap�U�Xnt��PvKen�CTqH�5�0�YELLOW� BO?Y��� Arc�0vis��C�h�WeldQci�al4Izt�Op�� ��gs�` 2@�a6��poG yRjcT1 NE�#HTf� xyWb��! �p��`gd`���p\� �=P��JPN ARCP*PR�A�� �OL�pSup̂fil�p��J�� n��cro�670�1�C~E�d��SS�pe.�tex�$ �P� �So7 t� ssa%gN5 <Q�BP:� 2�9 "0�QrtQCr��P�l0dpn������rpf�q�e�ppm�ascbin�4psyn�' pstx]08�HEL�NCL VIS �PKGS �Z@M�B &��B J8�@IPE GET_VAR FI?S_ (Uni� LU��OOL: ADD��@29.FD�TC4m���E�@DVp����`A�ТNO WT?WTEST �� ��!��c�FOR ^��ECT �a!� �ALSE ALA�`�CPMO-13�0��� b D: H�ANG FROM�g��2��R709� DRAM AV�AILCHECK�S 549��m�V�PCS SU֐L_IMCHK��P�0~x�FF POS� �F�� q8-12 CHARS��ER6�OGRA ���Z@AVEH�AME��.SV��Вאqn$��9�m "y��TRCv� SHA�DP�UPDAT �k�0��STATI���� MUCH ����TIMQ MOTN-003���@OBOGUI�DE DAUGH໱�b��@$tou�� �@C� �0��PA�TH�_�MOVE�T�� R64��V�MXPACK M�AY ASSERyTjS��CYCL`��TA��BE CO�R 71�1-�AN���RC OPTI�ONS  �`��A�PSH-1�`fi	x��2�SO��B��XO򝡞�_T��	�i�j�0j��du�byz �p wa��y�٠H�I������U�pb X?SPD TB/�F�_ \hchΤB0����END�CE�06�\Q�p{ sma'y n@�pk��L} ��traff#��	� ��~1fro�m sysvar/ scr�0R� ��Nd�DJU���H��!A��/��SET GERR�D�P7�����NDANT S�CREEN UNREA VM �P�D�D��PA���R~�IO JNN�0��FI��B��GRwOUNנD Y��Т٠�h�SVIP� 53 QS��DI�GIT VERS���ká�NEW�� �P06�@C�1IMCAG�ͱ���8� �DI`���pSSU�E�5��EPLAN� JON� DELL���157QאD��CALLI���Q��m���IPND}�IMG N9 PZ�{19��MNT/���ES ���`LocR Hol߀=��2�P�n� PG:��=�M��can����С�: 3D mE2view d X���ea1 �0b�po;f Ǡ"HCɰ��ANNOT AC�CESS M c�pie$Et.Qs �a� loMdFle�x)a:��w$qmo+ G�sA9�-'p~0̿�h0pa��eJ AUTO-�0��!�ipu@Т<ᡠIA�BLE+� 7�a F�PLN: L�p�l m� MD<�V�I�и�WIT H�OC�Jo~1Qu�i��"��N��US�B�@�Pt & r�emov���D�vAxis FT_7�PGɰCP:�O�S-144 � h� s 268QՐO�ST�p  CRA�SH DU��$P~��WORD.$��LOGIN�P��P�:	�0�046 i�ssueE�H�:� Slow st�c�`6�����z��IF�IMPR��SPOT:Wh4����N1STY��0V�MGR�b�N�CA�T��4oRRE�� �� 58�1��:N%�RTU!Pe -M .a�SE:�@pp���$AGpL��m@�all��*0a�OC�B WA���"3 �CNT0 T9DW�roO0alarm8�ˀm0d t�M��"0�2|� o�Z@O�ME<�� ��E%  ;#1-�SRE��M��st}0g   �  5KANJI~5no MNS@��INISITA7LIZ'� E�f�cwe��6@� dr�@� fp "��SC�II L�afai�ls w��SY�STE[�i�� � � Mq�1QGro8�m n�@vA�����&��n�0q��R�WRI OF L|k��� \ref"��
�up� de-r�ela�Qd 03�.�0SSchőb�etwe4�INDo ex ɰTPa�#DO� l� �ɰ�GigE�sope�rabil`p l�,��HcB��@]�lye�Q0cflxz�8Ð���OS {�����v4pfigi GL�A�$�c2�7H� wlap�0ASB� �If��g�2 l\�c�0�/�E�� �EXCE 㰁�P����i�� o0��G�d`]Ц�fq�l lsxt��EFal����#0�i�O�Y�n�CL�OS��SRNq1NT^�F�U��FqKP~�ANIO V7/�¥�1�{����DBa �0��ᴥ�ED��DET|�'� �b�F�NLINEb�B�UG�T���C"RL�IB��A��ABC? JARKY@���� rkey�`IL����PR��N��ITG+AR� D$�R �Er *�T��a�U�0��h�[�ZE V�� TASK p7.vr�P2" .�XfJ�srn�S谥d�IBP	c���B/��BUS��UNN�� j0-�{��cR�'���LOE�DIVS�CULs$cb����BW!��R~�W`�P�����IT(঱t�ʠ�OF��UNE�Xڠ+���p�FtE���SVEMG3`N�ML 505� D�*�CC_SAFE��P*� �ꐺ� PE�T��'P�`�F  �!���IR����c Ri S>� K��K��H GUNCHGz��S�MECH��IM��T*�%p6u���tPORY LE�AK�J���SP�EgD��2V 74\GRI��Q�g��oCTLN��TRe `@�_�p ���EN'�IN������$���r��T3)�i�STO��A�s�L��͐X	���q��Y� ��CTO2�J m��0F<�K����DU�S��O���3 9�J F��&���SSVGN�-1#I���RSRwQDAU�Cޱ� �T6��g��� 3�]���BR�KCTR/"� �q\�j5��_�Q�S�qI{NVJ0D ZO�P ݲ���s��г�Ui ɰx̒�a�DUAL�� J50e�x�RV�O117 AW�T�H!Hr%�N�247�%�52��|�&aol� ���R���at�Sd��cU���P,�LER��iԗQ0�ؖ  S!T���Md�Rǰt�_ \fosB�A�0@Np�c����{�U���ROP 2�b�pB>��ITP4M��b !AUt c0< � �plete�N@�� z1^qR635� (AccuCa�l2kA���I) �"�ǰ�1a\�Ps ��ǐ� bЧ0P������ig\cba?cul "A3p_ �1��ն���eta�ca��AT���PC��`�����_p�.�pc!Ɗ��:�cicrcB���5�tl��Bɵ�:�fm+�Ί��V�b�ɦ�r�upf�rm.����ⴊ�x�ed��Ί�~�ped�A�D �}b�ptl�ibB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆Ϙ���c�Ӳ�5�1j>�����tcȐ�Ϣ	�r����mm 1���T�sl^0��T�m�ѡ�#�rm3��u8b Y�q�std}��3pl;�&�ckv�=߆r�vf�䊰��9�v1i����ul�`�04fp�q �.f���� daq; i Da�ta Acqui+si��n�
��4T`��1�89���22 DMCM oRRS2Z�75���9 3 R710,�o59p5\?T "��1 (D�T� nk@���� ����E Ƒȵ��Ӹ��etdmm ��ER�����gE��1�q\mo?۳�=( G���[(

�2�` �! �@JMAC�RO��Skip/Offse:�a���V�4o9� &qR6C62���s�H��
 6Bq8����9~Z�43 J77� =6�J783�o `��n�"v�R5�IKCBq2 PT�LC�Zg R�3; (�s, �������03�	зJ���\sfmnmc? "MNMC�����ҹ�%mnf�FM�C"Ѻ0ª etm�cr� �8����� ,�}D��}   874\prdq>�,jF0���axi�sHProcess Axes e�wrol^PRA
��Dp� 56 J81�j�59� 56o6�� ���0w�690 998� [!IDV�1��2(x2��2ont �0�
����m2����?C��etis "ISD��9�� F/praxRAM�P�8 D��defB�,��G�isbasicHB�@޲{6�� W708�6��(�Acw:������D
�/,��AMOX�� ��DvE ��?;T��>Pi� RACFM';�]�!PAM�V �W�Ee�U�Q'
bU�75�.�ceN�e� nterfa�ce^�1' 5&!5�4�K��b(Dev am±�/�#���/<�Tazne`"DNEWE����btpdnui� �AI�_s2�d_rsono���bAs�fjN��bdv_arFvf�xhpz�}w��shkH9xstc��gAponlGzv{�ff��r���z��3{q'Td>pcOhampr;e�p� ^5977��	܀�4}0��mɁ�/�����l�f�!�pcchmp�]aMP&B�� �m�pev�����p�cs��YeS�� M/acro�OD��16Q!)*�:$�2U"_,x��Y�(PC ���$_;������o��J�g�egemQ@GEM�SW�~ZG�gesn�dy��OD�ndda��S��syT�Kɓ�Csu^Ҋ���n�m��<�L��  ���9:�p'ѳ޲��spotplusp���`P-�W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\f�eatu 0FEA�WD�oolo�s�rn'!2 p���a؝As3��tT.� (?N. A.)��!�e!�J# (j�,`��oBIB�oD -��.�n��k9�"K���u[-�_���p� "PSEqW����?wop "sEЅ� &�:�J������y�|� �O8��5��Rɺ��� ɰ[��X������ـ%�(
ҭ�q HL �0k�
�z�a!�B�Q�"(g�Q����� ]�'�.�����&���<�0!ҝ_�#��tpJ�H� ~Z��j�����y���� ��2��e������Z�� ��V��!%���=�]�p͂��^2�@iRV� Kon�QYq͋JF0B� 8ހ�`�	(^>�dQueue���X�\1�ʖ`�+F1tpv�tsn��N&��ftupJ0v �RDV�	�f��J1 Q���v��en��kvst�k��mp��btk�clrq���get����r��`kack�XZ��strŬ�%�st0l��~Z�np:!�`����q/�ڡ6!l��/Yr�mc�N+v�3�_� ����.�v�/\jF���� �`Q�΋ܒ�N50 (FRA��+�����fraparm���Ҁ�} 6�J6�43p:V�ELSE�
#�VAR $�SGSYSCFG�.$�`_UNITS 2�DG~°@�4�Jgfr��4A�@FRL-��0ͅ�3ې���L �0NE�:�=�?@�8 �v�9~Qx304��;�BPRSM~QA��5TX.$VNUM_OL��5��DJ�507��l� Functʂ"qwAP��琉�3 H�ƞ�kP	9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TP�PR���QA�prnaSV�ZS��AS8D�j510U�-�`cAr�`8 ��ʇ�DJR`�jYȑH  ��Q �PJ6�a2�1��48AA�VM 5�Q�b0 �lB�`TUP xb?J545 `b�`�616���0V�CAM 9�CwLIO b1�s5 ���`MSC8��
rP R`\s�STYL MNI�N�`J628Q  �`NREd�;@�`�SCH ��9pDCSU Mete�`�ORSR Ԃ�a0�4 kREIO�C �a5�`542�b9vpP<�nP�a�`�R�`7�`�M?ASK Ho�.r�7 �2�`OCO :��r3��p�b�p���r0X��a�`13\�mn�a39 HR�M"�q�q��L�CHK�uOPLG� B��a03 �q.��pHCR Ob�pC�pPosi�`fP6� is[rJ554��òpDSW�bM�D8�pqR�a37 }Rjr30 �1�s4 �R6�m7��52�r5 �2.�r7 1� P6����Regi�@T^�uFRDM�uSaq�%�4�`930�uS�NBA�uSHLB�̀\sf"pM�N{PI�SPVC�oJ520��TC�`�"MNрTMIL��IFV�PAC �W�pTPTXp6�.%�TELN N� Me�09m3�UECK�b�`U�FR�`��VCOR^��VIPLpq89q�SXC�S�`VVF��J�TP �q��Rw626l�u S�`�Gސ�2IGU�I�C��PGSt�\ŀH863�S�q������q34sŁ6�84���a�@b>�3� :B��1 T��9�6 .�+E�51 �y�q53�3�b1 ̛��b1 n�jr9 <���`VAT ߲�q�75 s�F��`�sA�WSM��`TOP u�ŀR52p���a�80 
�ށXY �q���0 ,b�`8855�QXрOLp}��"pE࠱tp�`LCyMD��ETSS�挀6 �V�CPEs oZ1�VRCd3�
�NLH�h��0011m2Ep��3 f��p���4 /165CR��6l���7PR���008 tB��9 o-200�`U0�p�F�1޲1 ��޲2 L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�J�?7 rbcfA�L��8\PC����"�32�m0u�n�K�Rٰn�5� 5EW
n�99 z��40 kB���3 ��6ݲ�`00�iB/��6�u��7�u��8 µ������s�U0�`�t �1 0�5\rb��2 E@���K���j���5˰��60��a�HУ`:Ł63�jAF�_���F�7 ڱ݀H�8�eHЋ�&�cU0��7�p���1u��8u��9 c73������D7� r��5t�97 ��E8U�1��2��1�)1:���h��1np�"���8(�U1��\pyl��,࿱v ��B�854��1V���D�-4��im��1�<����>br�3pr�48@pGPr�6 B����$�p��1����1�`͵�155ض157 �2��62�S����B��1b��2����1Π2"�2���B6`�1<c�4 7B�5i DR��8_�B/���187 uJ�8 ;06�90 rBn��1 (��202 /0EW,ѱ2^��2��90�U2�p�2��S2 b��4��2�a�"RB����9\�U�2�`w�l���4 6	0Mp��7������b�,s
5 ��3����<pB"9 3 ����l�`ڰR,:7 �2��V�2��5���2^H��a^9���qr�����n�5����5᥁""�8a�Ɂ}�5B���5����`UA���� ���86 �6 S�0�5�p�2�#�52�9 �2^�b1
P�5~�2`���&P*5��8��5��u�r!�5��ٵ544��%5��R�ąP nB^,z�c (�4���L���U5J�V�5��1�1^��%�����5 b21��gA���58W82� r�b��5N�E�589�0r� 1�95  �"������c8"a��|�L ���!J"5|6���^!�6��B�"8P�`#��+�8%�6B��AME�"1 iCN��622�Bu�6V���d� 4��84�`A�NRSP�e/S� C�5� �6� ��� \� �6� �V� 3�t��� T20CA�R��8� Hf� 1D�H�� AOE� ��� ,�|�� a�0\�� �!64K���ԓrA� �1 (M{-7�!/50T� [PM��P�Th:1�C��#Pe� �3�0� 5>`M75T"� �D�8p� �0Gc� u�4|��i1-710i�1B� Skd�7j�?6�:-HS,� �RN�@��UB�f�X�=m7C5sA*A6an���!X/CB�B2.6A �0 ;A�CIB�A�2�QF1�U�B2�21� /70�S� �4����Aj1��3p���r#0 B2\m*A@C��;bi"�i1K�u"A~AAU� imm7c7��ZA@HI�@�Df�A�D5*A��E� 0TkdR1�35�Q1�"*�@�Q�1�QC )P�1*A�5*A�EA�5XB�4>\77
B7=Q �D�2�Q$B�E7�C�D%/qAHEE�W7�_|` jz@� 2�0�Ejc�7�`�E"l7�@7@�A
1�E�V~`�W2%Qr�R9ї@0L_�#�����"A���b��H3s=rA/2�R5nR 4�74rNUQ1ZU�A�sw\m9
1M92L2��!F!^Y�ps� 2c1i��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHsXBSt62�q`s������ ��Pxq3530_*A3I)�2�db�u0�@� '4TX�m0�pa3i1A3s0Q25�c��st�r�VR1%e�q0
��j1 ��O2 �A�UEiy�@.�‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?P Q��qA!Pvs� 5	1 5aU���?PŅ���ဝQ9A6�zS*�7�qb5�1����Q��'00P(��V7]u�a itE1���ïp?7� �!?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ�޵y00\ry�"R�2BL�tN  ���� �1D�A}�2�qeR�5���_b�3�X]1m1l�cqP1�a�E�Q� 5�F����!5���@M-16Q�� f���r���Q�e� ��� PN�L�T_�1��i1��945�3��@�e�|�b1l>F1u*AY2�
�R8�Q����RJ�J13�D}T� 85
Qg� /0��*A!P�*A�Ð�d����2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt]1 ^u�ajrI�B����~`�|I�b��yI�\m�Qb�I�uz�A�c3Apa\9q� B6S��S��m���}�85`N�N�  �(M�� �f1���6����161j��5�s`�SC���U��A����5\se�t06c����10��y�h8��a6��6x��9r�2HS �� �Er���W@}�a��IlB���Y�ٖ�m�u �C����5�B��B��h`�F���X0���A :���C�M��AZ��@��4�6i����� e�O�-	���f1��F  �ᱦ�1F�Y	���GT6HL3��U66~`Ȗ��U�dU�9D20Lf0��Qv� ��fjq ��N������0v
� ���i	�	��72l�qQ2������� \�chngmove�.V��d���@2l_arf	�f ~��6������9C��Z���~���kr41@ S���0��V��t�����U�p7nu�qQ%�A]��V�1\"�Qn�BJ�2W� EM!5���)�#:��64��F�e50S �\��0�=�PV�� �e������E������m7shqQSH"U��)��9�!A���(���� �,�}�ॲTR11!��,�60e=��4F�����2��	 R-����������@�Ж��4���LS0R�)"�!lOA��Q�X) %!� 16�
U /��2�"2�E�9p���2>X� SA/i��'�
7F�H�@!B�0�� �D���5V��@2cV E��p��T��pt갖��1L~E�#�F�Q��9�E�#De/��RT��59���	�A�EiR���|����9\m20챃20��+�-u�19r4 �`�E1�=`O9`� �1"ae��O�2��_\$W}am41�4�3��/d1c_std ��1)�!�`_T��r~�_ 4\jdg�a �q�PJ%!~`-�r�+�bgB��#c300D�Y�5j�QpQb1�`bq��vB��v25�Up�����qm43�  �Q<W�"PsA��e ����t�i�P�W .��c�FX.�e4�kE14�44�~o6\j4�443sxj��r�j4up�� �\E19�h�PA�T�= :o�APf��coWol!\�2a��2A;_	2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a�:88J9X�l5�m�1a첚��*���(85�&�������P6���R,52&A����,fA9IfI50\u�z�OV
�v��}E�֖J���Y>� 16�r�C�Y��;��1��L ���Aq�&ŦP1��vB�)e�m�����1pĻ �1D�}�27��F�KAREL �Use S��FC�TN��� J970�FA+�� (�Q޵0�p%�)?�Vj9F?(��j�Rtk208 C"Km�6Q�y�j��iæPr�9�s#��v��krcfp�RCF�t3���Q��kcctme�!ME�g����^6�main�dV�� ��ru��kDº��c���o����J�dt��F �»�.vrT�f�����E%�!��\5�FRj73B�K����UER�HJ�O  �J�� (ڳF���F �q�Y�&T��p�F�z��19�tkvBr���V�Bh�9p�E�y�<�k�������;�v���"CT��f����)�
І ��)�V	�6���!� �qFF��1q���=��� ��O�?�$"���$���je���TCP A�ut�r�<520 �H5�J53E19�3��9��96�!8���9��	 �B574V��52�Je�(�� Se%!Y�����u���ma�Pqtool��ԕ������co�nrel�Ftro�l Reliab�le�RmvCU!��H51����� a�551e"�CNRE¹I�c�&���it�l\sfut?st "UTա��"X�\u��g@�i�D6Q]V0�B,Eѝ6A� �Q�)C���X���Yf�I�1|6s@6i��T6IU��vR��d�
$e%1��2�C58�E6��8�Pv�iV�4OFH58SOeJ� mnvBM6E~O58�I �0�E�#+@�&�F�0 ���F�P6a���)/++��</N)0\tr1x�����P ,�}ɶ��rmaski�ms�k�aA���ky'd�h�	A	�P�sDisp_layIm�`v��~��J887 ("A��+Heůצprd�s��Iϩǅ�h�0p�l�2�R2��:�Gt�@��PRD�TɈ�r��C�@Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��Px^@�P�firmQ� ���Pp�2�=bk�6�r��3��6��tppl��PL���O�p<b�ac�q	��g1J�U�d0�J��gait_9e���Y�&��Q���	�S�hap��erat�ion�0��R6�7451j9(`sGen�ms�42-f�Ár�p�5����2�rsgl�E��p�G���qF�205p�5S���ՁN�retsap�BP�O��\s� "GC�R�ö? �qngda�G��V��st2axU��Aa]��b�ad�_�btpu�tl/�&�e���tp�libB_��=�2.p����5���cird��v�slp��x�hex��v�re?�Ɵx�gkey�v�pm���x�us$�6�gcr��F������[�q27�j92�v�ollismqSk�9O��>�� (pl.���t��p!o��29$Fo8���cg7no@�tptwcls` CLS�o�b�\�km�ai_
�!s>�v�o	�t�b��x�ӿ�E�H��6~�1enu501�[�m��utia|$c�almaUR��Ca�lMateT;R5	1%�i=1]@-��/V�� ��Z�� �fq1�9 "K9E�L����z2m�CLMTq��S#��et �LM�3!} �F�c�ns�pQ�c���c_mo4q��� ��c_e���F��su��ޏ �_ �x@�5�G�join�@i�j��oX���&cW0v	 ���N�ve��C�clm�&Ao# �|$�finde�0�STD ter� FiLANiG���R��
��8n3��z0Cen���r,������J��� �� ���K��Ú�=�К�_Ӛ��r� "FNDR�� 3��}f��tguid��`��N�."��J�tq��  �������������J����_������c���	m�Z��\fndr.��n#>
B2�p��Z�CP Ma�����38A��� c
��6� (���N�B ������� 2�$�	81��m_���"ex�z5�.Ӛ��c���bSа�ef�Q��	��RBT~;�OPTN � +#Q�*$�r*$��*$r *$%/s#C�d/.,P�/|0*ʲDPN���$���$*�Gr�$ko Exc�'IF�$�MASK�%93 {H5�%H558�$_548 H�$4-1��$��#1(�$�0 E�$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3��9j0"M�49�4 � ��4�4tp�sh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E�\���5�A�4��3a�dq\�5K979�":E�ajO l "�DQ^E^�3i�Dq� ��4ҲO ?R�? ��q�5��T��3rAq�O�Lst�5~��7�p�5��REJ#�2�@a�v^Eͱ�F���4��.��5y N� �2il�(in�4��31 aJH1�2Q4�251ݠ��4rmal� �3) �REo�Z_�æOx�����4��^F�?onor Tf��7_ja�UZҒ4l��5rmsAU�Kkg���4�$HCd\�fͲ�e�ڱ�4�REM���4y�ݱ"u@�RER593�2fO��47Z��5lity,�U��e"DGil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe�=$��^�
E��u�IAymptm�U��BU��vste�y\�3��me� b�DvI�[�Qu�:F�U�b�*_�
E,�su$��_ Er��oxx���4huse�E-�?�sn�������FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��� b���(��1�� �c��Y�R�� �>�P� ��W��������'��0ɵ�[��͂����  � ,�N@� �A��bumpšf��B*�Box%��7Aǰ�60�BBw���MC� u(6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`���)���\bbk968� "�4�ω�bb��9va69����etbŠ��X�����#ed	�F��u�f�& �sea"������'�\��,���b�ѽ"�o6�H�
�x�$�f���!y���Q[�!� tperr�f�d� TPl0o� R/ecov,��3D���R642 � 0���C@}s� N@��(NU�rro���yu2�r��  �
�  ����$$�CLe� �������������$~z�_DIGIT��.������ .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ oo$j��+c:PRODUCTM��0\PGSTKD��V&ohozf99���D���$F�EAT_INDE�X��xd���  
�`IL�ECOMP ;����#��`�cS�ETUP2 <��e�b�  �N �a�c_AP2�BCK 1=�i  �)wh0?{%&c����Q� xe%�I�m�� �8��\�n����!� ��ȏW��{��"��� F�Տj���w���/�ğ S���������B�T� �x������=�үa� �����,���P�߯t� �����9�ο�o�� ��(�:�ɿ^���� �ϸ�G���k� �ߡ� 6���Z�l��ϐ�ߴ� ��U���y����D� ��h��ߌ��-���Q� ��������@�R��� v����)�����_��� ��*��N��r� �7��m�@&�3\�i
pP� 2#p*.V1Rc�*��`� /��PC/|1/FR6:/"].��/+T�`�/ �/F%�/�,�`r/?��*.F�8?	�H#&?e<�/�?;STM �2�?�.K �?��=iPen�dant Panel�?;H�?@O�7�.O�?y?�O:GIF �O�O�5�OoO�O_:JPG _J_�56_�O�_�_�	PANE�L1.DT�_@�0�_�_�?O�_2�_�So�WAo�_o�o�Z3 qo�o�W�o�o�o)�Z4�o[�WI���
TPEINSO.XML��0�\���qCust�om Toolb�ar	��PAS�SWORDy�FRS:\L�� �%Passwo�rd Config���֏e�Ϗ�B 0���T�f�������� ��O��s������>� ͟b��[���'���K� �򯁯���:�L�ۯ p�����#�5�ʿY�� }��$ϳ�H�׿l�~� Ϣ�1�����g��ϋ�  ߯���V���z�	�s� ��?���c���
��.� ��R�d��߈���;� M���q������<��� `������%���I��� �����8����n ���!��W�{ "�F�j| �/�Se��/ �/T/�x//�/�/ =/�/a/�/?�/,?�/ P?�/�/�??�?9?�? �?o?O�?(O:O�?^O �?�O�O#O�OGO�OkO }O_�O6_�O/_l_�O �__�_�_U_�_y_o  o�_Do�_ho�_	o�o -o�oQo�o�o�o�o @R�ov��; �_���*��N� �G������7�̏ޏ m����&�8�Ǐ\�� ���!���E�ڟi�ӟ ���4�ßX�j����� ���įS��w�������B�#��$FIL�E_DGBCK �1=��/���� ( ��)
SUMMA�RY.DGL����MD:������Diag Sum�mary��Ϊ
C?ONSLOG������D�ӱCon�sole log�E�ͫ��MEMCHECK:�!ϯ����X�Memory� Data��ѧ��{)��HAD�OW�ϣϵ�J����Shadow C?hangesM�'��-��)	FTAP7Ϥ�3ߨ���Z��mment TB�D��ѧ0=4)�ETHERNET��������T�ӱE�thernet �\�figurat�ionU�ؠ��DCSVRF�߽߫������%�� ve�rify all���'�1PY���DIFF�����[����%��diff]������1R�9�K���� ���X=��CHGD������c��r�����2ZAS� ��GD����k��z��FY�3bI[� �/"GD����s/����/*&UPDATES.� ��/��FRS:\��/�-ԱUpda�tes List��/��PSRBWLOD.CM(?���"�<?�/Y�PS_ROBOWEL��̯�? �?��?&�O-O�?QO �?uOOnO�O:O�O^O �O_�O)_�OM___�O �__�_�_H_�_l_o �_�_7o�_[o�_lo�o  o�oDo�o�ozo�o 3E�oi�o�� �R�v���A� �e�w����*���я `���������O�ޏ s������8�͟\�� ���'���K�]�쟁� ���4���ۯj����� �5�įY��}���� ��B�׿�x�Ϝ�1� ��*�g�����Ϝ��� P���t�	�ߪ�?��� c�u�ߙ�(߽�L߶� �߂���(�M���q�  ���6���Z���� ��%���I���B������2�����h�����$FILE_� P�R� ��������M�DONLY 1=�.�� 
 � ��q��������� �~%�I�m �2��h� �!/�./W/�{/
/ �/�/@/�/d/�/?�/ /?�/S?e?�/�??�? <?�?�?r?O�?+O=O �?aO�?�O�O&O�OJO �O�O�O_�O9_�OF_�o_
VISBCK�L6[*.VD�v_�_.PFR:\��_�^.PVis�ion VD file�_�O4oFo\_ joT_�oo�o�oSo�o wo�oB�of�o �+����� ��+�P��t���� ��9�Ώ]�򏁏��(� ��L�^�������5� ��ܟk� ���$�6�ş�Z��~�����
M�R_GRP 1>�.L��C4 w B���	 W������*u����RHB ���2 ��� ��� ���B� ����Z�l���C���D�ি����Ŀ��K���L6��J���F�5UT?w�Q�0!����ֿ G,�F�I�/E���.���9:�]�@��'�A&�#�A�|f�?�f��A��r��E�� F@ ��������J��NJ�k�H9�H�u��F!��IP�s�?����(��9�<9��896C'�6<,6\b� �+�&�(�a�L߅�X���A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�P=��P��T���ܿ� �B���/ ��@�33�:��.�g&�@U�UU�U��q	>u?.�?!rX���	�-=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7��:����D�@ ?D�� Cϥ��C������Q�,/� �����/M��/q��/ �/�/�??:?%?^? p?[?�??�?�?�?�?  O�?�?6O!OZOEO~O iO�O�O�O�OW�ߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������X[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U�� 
//./�v���/ ���/�/�/�/�/� !?3?E?W?i?�/?�? �?�?�?�?�?��� AO�?eO�/�O�O�O�O �?�O�O__+_NO�O J_s_�_�_�_�_
OO .OoB_'ovOKo]ooo �oP_>o�o�o�o�oo �o5GYk}�_ �_�_��8o�� 1�C�U�$y������� �ӏf���	��-�?� ����Ə���ϟ �����;�M�_� q���.�(���˯ݯ� �P�b�t�����m��� ������ǿٿ����� !�3�E�h��{ύϟ� �����$�6�H�J�/� ~�S�e�w߉ߛ�jϿ� �������*߬�=�O��a�s��YT_ER�R J5
���P�DUSIZ  j��^J����>��?WRD ?t���  guest}��%�7��I�[�m�$SCDMNGRP 2Ktw�������V$�K�� 	�P01.14 8~��   y�����B   � ;����� ����������
 �������?�����~����C.gR|����  i  ��  
��������� +�������
���l �.r���"�l��� m
d����|��_GROU��]L�� �	�����07EQUPD'  	պ�J��TYa ����T�TP_AUTH �1M�� <!iPendany���6�Y!K?AREL:*��
-KC///A/ �VISION �SETT�/v/� "�/�/�/#�/�/
? ?Q?(?:?�?^?p>�CTRL N�����5�
�.?FFF9E3�?��FRS:DEF�AULT�<F�ANUC Web Server�:
�����<kO}O�O�O�O�O��WR_C�ONFIG OΡ� �?��ID�L_CPU_PC�@�B��7P�;BHUMIN(\��~<TGNR_IO�������PNPT_�SIM_DOmV�w[TPMODNT�OLmV �]_PR�TY�X7RTOLN/K 1P����_�o!o3oEoWoio�RMASTElP��R��O_CFG�o�iU�O��o�bCYCL�E�o�d@_ASG� 1Q����
  ko,>Pbt�� �������sk.�bNUM����K@�`IPCH�o��`RTRY_CN@xoR��bSCRN����Q��� �b�`�b�R���Տ��$�J23_DSP_�EN	����OBPROC�U�i�JOGP1SY@~��8�?�!��T�!�?*�POSR�E�zVKANJI�_�`��o_�� ��T��L�6͕����CL�_LGP<�_���EY�LOGGIN�`���LANG?UAGE YF7R�D w���LG���U�?⧈�xR� �����=P��'0��$ N�MC:\RSCH�\00\��LN_DISP V��`
��������OC�R�.RDzVTA{�OGBOOK W
{���i��ii��X �����ǿٿ����1�"��6	h������e�?�G_BU_FF 1X�]��2	աϸ����� ������!�N�E�W� ��{ߍߺ߱�����������J���DC�S Zr� =����^�+�ZE���������a�IO 1[�
{ ُ!� � !�1�C�U�i�y����� ����������	- AQcu��������EfPTM  �d�2/ASe w������� //+/=/O/a/s/�/8�/��SEV���]�TYP`�/??y͒�RS@�"��×�FL 1\
������?�?�?`�?�?�?�?/?TP6���">�NGN�AM�ե�U`�UP�S��GI}�𑪅�mA_LOAD�G� %�%DF_MOTN���O�@�MAXUALRM <��J��@sA�Q����QWS ��@C �]m�@-_���MP2�7�^
{� ر�	�!�P�+ʠ�;_/��R1r�W�_�WU�W�_ ��R	o�_o?o"oco Noso�o�o�o�o�o�o �o�o;&Kq\ �x������ �#�I�4�m�P���|� ��Ǐ���֏��!�� E�(�i�T�f�����ß ��ӟ���� �A�,� >�w�Z�������ѯ�� ��د���O�2�s� ^�������Ϳ���ܿ��'��BD_LDX�DISAX@	��M�EMO_APR@E� ?�+
  � *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT ��Q�c�Ϝ߇��ߧ� ����w����>�)�b� t�[����{����� �����:���I�[�/� �����������o��� ��6!ZlS� �s����2 �AS'�w�� ��g��.//R/�d/�_MSTR �`�-w%SCD 1am͠L/�/H/�/ �/?�/2??/?h?S? �?w?�?�?�?�?�?
O �?.OORO=OvOaO�O �O�O�O�O�O�O__ <_'_L_r_]_�_�_�_ �_�_�_o�_�_8o#o \oGo�oko�o�o�o�o �o�o�o"F1j Ug������ ���B�-�f�Q����u�����ҏh/MKC_FG b�-�~�"LTARM_���cL�� �σQ�N�<�METsPUI�ǂ���)�NDSP_CMN�Th���|�  	d�.��ς�ҟܔ�|�POSCF�����PSTOL 1�e'�4@�<#�
5�́5�E�S�1�S� U�g�������߯��ӯ ���	�K�-�?���c��u�����|�SING_CHK  ��^;�ODAQ,�f���Ç��DEV }	L�	MC:!̟HSIZEh��-���TASK %�6�%$123456789 �Ϡ��TRIG 1g�+ l6�%���ǃ`�����8�p�YP[�� ��EM_INF� 1h3� �`)AT&�FV0E0"ߙ�)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ������H�����A���AI�q�,��|���� ���ߵ�����J� ��n������W����� ������"����X� �/����e��� ���0�T;x� =�as��/� ,/c=/b/�/A/�/ �/�/�/��?�� �^?p?#/�?�/�?s? }/�?�?O�?6OHO�/ lO?1?C?U?�Oy?�O �O3O _�?D_�OU_z_�a_�_�ONITO�R��G ?5�  � 	EXEC�1Ƀ�R2�X3�X4��X5�X���V7�X8
�X9Ƀ�RhBLd�R Ld�RLd�RLd
bLdb Ld"bLd.bLd:bLdFb�Lc2Sh2_h2kh2�wh2�h2�h2�h2��h2�h2�h3Sh3�_h3�R�R_GRP_SV 1in����(ͅ�
�3w�8��r�ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A��W�@<�P�R�
h�B�b�A��j���a��:��Dzۀ���߹�����j���( �� -��C���'�7��&���q�Y������ �?�ff ���gy ������q+q��
>N+�  PƱj�(�� ��7	���|�/?����xZ�p�<
6b<߈�;܍�<�ê�<� <�&Jσ�AI�ɳ+����?fff?I�?y&�k�@�.��J<?�`� q�.�˴fɺ�/�� 5/����j/U/�/y/ �/�/�/�/�/?�/0?q��F�?l??��?/�?+)�?�?�E��� E�I�G+� F��?)O�?�9O_OJO�OnO�Of�BL޳B�?_h�.��O �O��%_�OL_�?m_�?��__�_�_�_�_�
��h�Îg>��_Co�_goRodo�oF�GA�ds�q�C�op�o�o|�����$]Hq���D��fpC���pCHm�ZZ7t���6q�q�����N'�3A�A��AR1AO�^?�$�?�K��0±
=ç>�����3�W
�=�#�W��e���9�����{����<���(�B�u�����=B0�������	L��H��F�G���G���H�U`E���C�+����I#�I���HD�F���E��RC�j=���
I��@�H�!H�( E<YD0q �$��H�3�l�W��� {��������՟��� 2��V�A�z���w��� ��ԯ�������� R�=�v�a��������� ���߿��<�'�`� Kτ�oρϺϥ����� ���&��J�\�G߀� kߤߏ��߳������� "��F�1�j�U��y� ������������0�@�T�?�Q����(�1g��3/E�����5������q�3�8�����q4�Mgs&IB�+2D�a���{�^^	���P���uP2P7Q4_A��M0bt��R����X��/   �/ �b/P/�/t/�/ *a@)_3/�/�/�%1a�?�/?;?M?_?q?  �?�/�?�?�?�?�O 2 F�$N�vGb�/�A��@X�a�`�qC��C@�o��O2���OF� �DzH@�� F�P D���O�O�ys<O!_3_E_W_i_~s?���@@pZ�.t22!:2~
 p_�_ �_�_	oo-o?oQoco�uo�o�o�o�o��Q ���+��1���$MSKCFMA�P  �5� �6�Q�Q"~��cONREL  �
q3�bE�XCFENB?w
8s1uXqFNC_Qt�JOGOVLIM�?wdIpMrd�bKE�Y?w�u�bRU�N�|�u�bSFSPDTY�avJu�3sSIGN?QtTO1MOT�Nq�b�_CE_GRP [1p�5s\r� ��j�����T��⏙� �����<��`��U� ��M���̟��🧟� &�ݟJ��C���7��� ����گ�������4��V�`TCOM_C_FG 1q}�V�p�����
P�_AR�C_\r
jyUA�P_CPL��ntN�OCHECK ?={ 	r ��1�C�U�g�yϋ� �ϯ���������	���({NO_WAITc_L�	uM�NTX��r{�[m�_E�RRY�2sy3�� &�������r��c� ��T_MO���t��, K��$�k�3�PARAM:��u{��V[ﰽ�!�u?�� =9@3�45678901 ��&���E�W�3�c������{������� �����=�UM_RSPACE ��Vv��$ODR�DSP���jxOF�FSET_CAR9Tܿ�DIS���PEN_FILE�� �q��c֮�OPT?ION_IO���PWORK v_�ms �P(��R�Q
�j.j	 ���Hj&6$� R�G_DSBL  ��5Js�\��R�IENTTO>p�9!C��PqfA� UT_SIM_D�
r�b� V� LCT ww�bc��|U)+$_PEXE�d&RATp �vju�p���2X�j)TUX�)TX�##X d-�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O�H2�/oO�O�O�O�O@�O�O�O�O_]�<^O ;_M___q_�_�_�_�_��_�_�_o���X�O�U[�o(��(����$o�,� ��IpB` @oD�  Ua?�[cbAa?��]a]�DWcxUa쪋l;�	lmb��`�x�J�`�����a�< ��`�� ��b, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�"���� �N	 W��  '!o�:q�pC	 C�@@sBq�|�:�� m�
�!�h@ߐ�n����Z��B	 �A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�'!��(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��W ��Ӱ�|�ɆDT Qy-����D � ��,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�T�(�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_j��_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ�_ ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������//�"#�$PGTRA�CELEN  �#!  ���" �8&_UP z���g!�o S!h 8!_�CFG {g%Q#"!x!�$J �"� |"DEFSPD� |�,!!J ��8 IN TRLW }�-" 8�(�IPE_CONF�I� ~g%��g!�$�$�"8 L�ID�#�-74G�RP 1�7Q!��#!A ����&ff"!A+33�D�� D]� ?CÀ A@+6�!�" d�$�9�9*1*0?� 	 +9�-+6�? ´	C�?�;B@3AO�?OIO3O�mO"!>�T?��
5�O�O�N�O =��=#�
�O _�O_J_5_n_Y_�O�}_�_y_�_�_�_  #Dzco" 
oBo �_Roxoco�o�o�o�o �o�o�o>)b�M��;
V7.10beta1�$�  A�E}�rӻ�A " ޼p?!G��q>˙��r��0�q̽ͻqBQ��qAA\�p�q�4�q�p�"�BȔ2�D�V�h�Bw��p�?�?)2{ ȏw�׏���4�� 1�j�U���y�����֟ ������0��T�?� x�c�������ү���� !o�,�ۯP�;�M��� q�����ο���ݿ� (��L�7�p�+9��sF@ �ɣͷϥ� g%������+�!6I� [߆������ߵߠ��� ������!��E�0�B� {�f���������� ���A�,�e�P��� t���������� ��=(aL^�� �����'9 $]�Ϛ��ϖ��� ����/<�5/`�r� �ߖߏ/>�/�/�/�/ �/?�/1??U?@?R? �?v?�?�?�?�?�?�? O-OOQO<OuO`O�O �O�O�O���O_�O)_ _M_8_q_\_n_�_�_ �_�_�_�_o�_7oIo t���o�o���o �o�o(/!L/^/p/�/ {*o������ ���A�,�e�P�b� ���������Ώ�� +�=�(�a�L���p��� ���Oߟ񟠟� �9� $�]�H���l�~����� ۯƯ���#�No`oro �on��o�o�o�oԿ ���8J\ng�� ��vϯϚ�������	� ��-��Q�<�u�`�r� �ߖ��ߺ������� ;�M�8�q�\������ ��z������%��I� 4�m�X���|������� ����:�L�^���Z ����������� $�6�H�Swb �������/ /=/(/a/L/�/p/�/ �/�/�/�/?�/'?? K?]?H?�?��?�?f? �?�?�?O�?5O OYO DO}OhO�O�O�O�O�O �O&8J4_F_�� ��_�_��_�_" 4-o�O*ocoNo�oro �o�o�o�o�o�o) M8q\��� ������7�"� [�m��?����R�Ǐ�� �֏�!��E�0�i� T���x��������_ $_V_ �2�l_~_�_������R�$PLID�_KNOW_M � �T������SV �v�U͠�U��
��.�ǟR�=��O�����mӣM_G�RP 1��!`0*u��T@ٰo�ҵ�
���Pзj�� `���!�J�_�W�i� {ύϟϱ��������Ϭ߱�MR�����T��s�w� s��ߠ� �߯߅��ߩ߻����� A���'����� ����������=�� �#���������}���ء��S��ST��1 �1��U# ���0�_ A .��, >Pb����� ���3(iL ^p������2*���<-/3/)/;/M/A4f/x/�/�/5�/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?MA/D  d#`�PARNUM � w�%OS+CH?J ME
�G`A8�Iͣ�EUPD`OrE�
a�OT_CMPa_��B@�P@'˥~TER_CHK'U���˪?R$_6[RqSl�¯��_MOA@�_�U_�_RE_RES_G ��>� oo8o+o\oOo�oso �o�o�o�o�o�o�o�W �\�_%�Ue  Baf�S� ��� �S0����SR0� �#��S�0>�]�b��S��0}������RV 1񈟥��rB@c]���t�(@c\�����D@c[��$���RTHR_ICNRl�DA��˥d,�oMASS9� ZM��MN8�k�MON_�QUEUE ����˦��x� RDN�PUbQN{�P[��E�ND���_ڙEXE�ڕ�@BE�ʟ��OPTIOǗ�[���PROGRAM %��%��ۏ�O~��TASK_IAD�0�OCFG ��tO��ŠDATA����Ϋ@��2 7�>�P�b�t���,��� ��ɿۿ�����#�5ϼG���INFOUӌ�������ϭϿ��� ������+�=�O�a� s߅ߗߩ߻�������h�^�jč� y�ġ?PDIT ��ίc���WERFL�
��
RGADJ7 �n�A�����?����@���IOR�ITY{�QV���M�PDSPH�����U�z����OTOE�y�1�R� (!AF4�E�P]���?!tcph����!ud��!�icm��ݏ6�X�Y_ȡ�R��ۡ)� *+/ ۠�W:F� j�������%7[B�*���PORT#�BC�۠����_CARTREP
�R� �SKSTAz��ZS�SAV���n�	�2500H863����r�$!�R�
���q�n�}/�/��'� URGE�Bl��rYWF� DO{��rUVWV��$�A�W�RUP_DELA�Y �R��$R_'HOTk��%O]?��$R_NORMA�Lk�L?�?p6SEM�I?�?�?3AQSKkIP!�n�l#x 	1/+O+ ORO dOvO9Hn��O�G�O�O �O�O�O_�O_D_V_ h_._�_z_�_�_�_�_ �_
o�_.o@oRoovo do�o�o�o�o�o�o�o *<Lr`����n��$RCV�TM�����pDkCR!�LЈq�Cl�fC���C��>?�A��>:��<l���4M�b�����O
�n��������{��4Oi��O <
�6b<߈;����>u.�??!<�&{�b� ˏݏ��8�����,� >�P�b�t��������� Ο���ݟ��:�%� 7�p�S������ʯܯ � ��$�6�H�Z�l� ~�������ƿ���տ ���2�D�'�h�zϽ� �ϰ���������
�� .�@�R�d�Oψߚ߅� �ߩ���������<� N��r������� ������&�8�#�\� G�����}��������� ��S�4FXj| ������� ��0T?x�u ����'//,/ >/P/b/t/�/�/�/�/ �/�/�?�/(??L? 7?p?�?e?�?�?��? �? OO$O6OHOZOlO ~O�O�O�?�?�O�O�O �O __D_V_9_z_�_ �?�_�_�_�_�_
oo�.o@oRodovo�X�qG�N_ATC 1��� AT�&FV0E0�k�ATDP/6/�9/2/9�hA�TA�n,A�T%G1%B96}0�i+++�o�,�aH,�qIO�_TYPE  �u�sn_�oREFPOS1 1�P{� x�o�X h_�d_����� K�6�o�
���.���R�x���{{2 1�P{���؏V�ԏz����q3 1��$�6��p��ٟ���S4 1�����˟���n�|��%�S5 1�<��N�`�����<���S6 1�ѯ���/�𭿘�ѿO�S7 1�f�x���ĿB�-�f�>�S8 1������Y�������y�SM�ASK 1�P � 
9�G��XNO�M���a~߈ӁqMOTE  h�~t��_CFG �������рrPL_RA�NG�ћQ��POW_ER ��e����SM_DRYP_RG %i�%���J��TART ��
�X�UME_P�RO'�9��~t_E�XEC_ENB � �e��GSPD�������c��TDB����RM��MT�_!�T���`O�BOT_NAME� i���iO�B_ORD_NU�M ?
�\q�H863  a�T��������b�PC_TIMEO�UT�� x�`S2�32��1��k �LTEACH PENDAN ��ǅ�}���`�Maintena�nce ConsțR}�m
"{�dKCL/Cg��Z ���n� No Use}�	���*NPO��х����(CH_�L�������	��mMAVAILȰ�{��ՙ�SPACE1 2��| d��(>���&���p��M,8�?�ep/eT/ �/�/�/�/�W//,/ >/�/b/�/v?�?Z?�/ �?�9�e�a�=??,? >?�?b?�?vO�OZO�?��O�O�Os�2� /O*O<O�O`O�O�_��_u_�_�_�_�_[3 _#_5_G_Y_o}_�_ �o�o�o�o�o[4.o@oRodovo$�o �o����"�	�7�[5K]o��A� ���	�̏�?�&�T�[6h�z������� ^�ԏ���&��;�\�C�q�[7�������� ͟{���"�C��X�y�`���[8����Ư دꯘ��0�?�`�#��uϖ�}ϫ�[G ��i� �ϋ
G� ����$�6� H�Z�l�~ߐ��8 ǳ�@����߈��d(� ��M�_�q���� ��������?���2� %�7�e�w��������� �����������!�R E�W�����������?Q; `�� @0�@�ߖrz	�V_ �����
/L/^/ |/2/d/�/�/�/�/�/ �/?�/�/�/*?l?~? �?R?�?�?�?�?�?�?�?2O�?
��O[�_MODE  ��˝IS ���vO,*ϲ�O-_���	M_v_#dCWO�RK_AD�M9{�P%aR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/$��:	d/JaR��WY��^���^R�^	r  P��� �  8��P�	�D��GYk}�� ������Qp/@/R//)P;�o\T��Q�pg-�t�_�DiKT��[  � lv%������/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OWW�#�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_olO~O d+No`oro�o�o�o�o �o�o�o&8J \n������u�  0�"0g�/� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q�����$o��˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�����Do ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������w
�  58�J�\�n߀� �ߜկ���������	� �-�?�Q�c�u������ ��-�� ��� �2�D�V�h�z���������������v���& ���%	12345�678�" 	�
�/� `r�������� (:L^p�� ����� //$/ 6/H/Z/l/~/��/�/ �/�/�/�/? ?2?D? V?h?�/�?�?�?�?�? �?�?
OO.O@Oo?dO vO�O�O�O�O�O�O�O __*_YON_`_r_�_ �_�_�_�_�_�_oo C_8oJo\ono�o�o�o �o�o�o�oo"4 FXj|���������	��s�3�E�W�{�Cz � Bp��   ��2���z�$S�CR_GRP 1��(�U8(�\�x^ @�  �	!�	 ׃���"� $� ��-��+��R�nw����D~������#����O����M-10iA 78909905 Ŗ~5 M61C >P4��Jׁ
� ���0�����#�1�	"�z�������4¯Ҭ ���c� ��O�8�J��� ����!�����ֿ��B�y�������r��A��$�  @���<� �R�?��d���H�y�u�O���F@ F�`�§�ʿ�϶� ������%��I�4�m� �<�l߃ߕߧ߹�B���\����1�� U�@�R��v����� �������;���*<=�
F���?�d�<��>m���@��:��� B����ЗЙ���EL_D�EFAULT  ������B�MIPOWERFL  �x$1 WFDO� $��ERVE�NT 1������"�pL!D?UM_EIP��8���j!AF_I�NE �=�!FIT���!���4 ��[!�RPC_MAIN�\>�J�nVI�Sw=���!�TP�PU��	d��?/!
PMON?_PROXY@/�Ae./�/"Y/�fz/��/!RDM_S�RV�/�	g�/#?!#R C?�h?o?K!
pM�/�i^?��?!RLSYN�C�?8�8�?O!�ROS�.L�4 �?SO"wO�#DOVO�O �O�O�O�O_�O1_�O U__._@_�_d_v_�_ �_�_�_o�_?ooco�iICE_KL �?%y (%SVCPRG1ho 8��e���o�m3�o�o"�`4 �`5(-"�`6PU�`7x}��`���l9��{ �d:?��a�o��a�o E��a�om��a���a B���aj叟a�� �a�5��a�]��a� ���a3����a[�՟�a �����a��%��aӏM� �a��u��a#����aK� ů�as���a��mob �`�o�`8�}�w����� ��ɿ���ؿ���5� G�2�k�VϏ�zϳϞ� ���������1��U� @�y�dߝ߯ߚ��߾� ������?�*�Q�u� `���������� ��;�&�_�J���n������������sj_�DEV y	��MC:Pϻ_OUT"�,REC 1q�Z� d  / 	 	�������
� �PJ�%6 (�&�[w֍,�*  �T - �- �A�- c|�P�� ���//B/0/f/ x/Z/�/�/�/�/�/�/ �/?�/?P?>?t?b? �?�?�?�?�?�?�?O OOLO:OpO�OdO�O �O�O�O�O�O�O$__ H_6_X_~_l_�_�_�_ �_�_�_�_ ooDo2o Tozo\o�o�o�o�o�o �o�o.R@v d����},� ���4�"�X�F�|� ��p�����֏ď�� ��0��@�f�T���x� ����ҟ�Ɵ���,� �<�b�P���h�z��� ���ί��(�:�� ^�L�n�p�������ܿ �п� �6�$�Z�H� jϐ�rϴϢ������� ���2�D�&�h�Vߌ� z߰ߞ����������� 
�@�.�d�R��ZjoV 1�w P��m��	>  � ��
T�YPEVFZN_CFG ��'d7�?GRP 1�A�c/ ,B� A� �D;� B����  B4R�B21HELL�:�(
� �X����%RSR ����E0iT� x�������/Sew�  ��%w��(���#��������2#�d�����HK 1��� �k/f/x/ �/�/�/�/�/�/�/? ?C?>?P?b?�?�?�?��?��OMM �����?��FTOV_�ENB ���+�HO�W_REG_UI�O��IMWAITrB�JKOUT;F���LITIM;E;���OVAL[OMC_UNITC�F+��MON_ALIA�S ?e�9 ( he��_&_8_J_ \_��_�_�_�_�_j_ �_�_oo+o�_Ooao so�o�oBo�o�o�o�o �o'9K]n ����t��� #�5��Y�k�}����� L�ŏ׏������1� C�U�g���������� ӟ~���	��-�?�� c�u�������V�ϯ� �����;�M�_�q� �������˿ݿ��� �%�7�I���m�ϑ� �ϵ�`�������ߺ� 3�E�W�i�{�&ߟ߱� �����ߒ���/�A� S���w����X�� ��������=�O�a� s���0����������� ��'9K]� ���b��� #�GYk}�: ������/1/ C/U/ /f/�/�/�/�/ l/�/�/	??-?�/Q? c?u?�?�?D?�?�?�? �?O�?)O;OMO_O
O �O�O�O�O�OvO�O_�_%_7_�C�$SM�ON_DEFPR�O ����`Q �*SYSTEM*�  d=OURECALL ?}`Y� ( �}4x�copy fr:�\*.* vir�t:\tmpba�ck�Q=>192�.168.4�P46:8144 �R��_�_�_�K}5�Ua��_�_�V�_goyo�o}�9�Ts:orde�rfil.dat�.l@oVo�o�o}0�Rmdb:+o�oRc �odv�a�_2o? U��
�o��So�d�v����
xyz�rate 61 �+�=�O������|����6788 �� ҏc�u����o�o56� ٟ���"��5�џ�b�t����6����e�mp:�6976 �W������.��*.d��Ʈϯ`�r�����1 +�=�O���� �)�Ҳ��ҿc�uχ� ����5�ͧ������� "���̨��b�t߆ߙ ����:�V�����������6 ��g�y�� �ϰ�9�T�����	�� ��@���c�u�����-� ?����������� N�_q����1��� ���&��J�[ m����7���� �"�F�i/{/ ����2/D/V/�/�/?��x284>��/a? s?�?��349�?�? �?"�?58�?bOtO��O���?��81392 WO�O�O�O��O�J �Oa_s_�_�/��<_N_ �_�_o?(?�S�_�_ couo�o�?�?5O�G�o �o�oO"O�o�H�ob t���/�/QcU� �
�/��T`�g� y����o�o9T��� 	���@ҏc�u�������$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1����?���% ֟��&�	��\�?� f���u��������ϯ ��"��F�)�;�|�_� ������ֿ��˿�� �B�%�f�I�[Ϝ�� ���ϵ�������,�� 6�b�E߆�i�{߼ߟ� ����������L�/� V��e������� �����6��+�l�O� v��������������� 2V9K�o ������� &R5vYk�� ���/��<// F/r/U/�/y/�/�/�/ �/?�/&?	??\??? f?�?u?�?�?�?�?�? �?"OOFO)O;O|O_O �O�O�O�O�O�O_�O _B_%_f_I_[_�__ �_�_�_�_�_�_,oo 6oboEo�oio{o�o�o �o�o�o�oL/ V�e����� ���6��+�l�O��v�������PARAoM �����_ �	��P�����OFT_�KB_CFG  �ヱ���PIN_�SIM  ����C�U�g�����RV�QSTP_DSB�,�򂣟����SR� �/�� & � ULTIROBOTTASK������TOP_O�N_ERR  ����PTN �/�@��A	�RING_P�RM� ��VD�T_GRP 1�<ˉ�  	���� ��������Я���� �*�Q�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߣߠ߲����� ������0�B�i�f� x������������ �/�,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZ�~���� ���/ /G/D/V/ h/z/�/�/�/�/�/�/ ?
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_�8___\_��VPRG�_COUNT�q�@���RENBU��UM�S��__UP�D 1�/�8  
s_�oo*oSo No`oro�o�o�o�o�o �o�o+&8Js n������� ��"�K�F�X�j��� ������ۏ֏���#� �0�B�k�f�x����� ����ҟ������C� >�P�b���������ӯ�ί�����UYS�DEBUG�P�P��)�d�YH�SP_PwASS�UB?Z��LOG ��U��S)�#�0� � ��Q)�
MC�:\��6���_MPAC���U���Qñ�8� �Q�SAV ������ǲ&��ηSV;�TEM�_TIME 1���[ (m�7&��4:�}YT1SVGgUNS�P�U'�U����ASK_OPTION�P�U�Q�Q���BCCFG 3��[u� n�A�a�`a�gZo��� �ߕ��߹������� :�%�^�p�[���� ������ �����6�!� Z�E�~�i���������&�������&8�� nY�}�?�� ԫ ��(L :p^����� ��/ /6/$/F/l/ Z/�/~/�/�/�/�/�/ �/�/2?8 F?X?v? �?�??�?�?�?�?�? O*O<O
O`ONO�OrO �O�O�O�O�O_�O&_ _J_8_n_\_~_�_�_ �_�_�_�_o�_ o"o 4ojoXo�oD?�o�o�o �o�oxo.TB x��j���� ����,�b�P��� t�����Ώ��ޏ�� (��L�:�p�^����� ��ʟ��o��6� H�Z�؟~�l������� د���ʯ ��D�2� h�V�x�z���¿��� Կ
���.��>�d�R� ��vϬϚ��Ͼ����� ��*��N��f�xߖ� �ߺ�8��������� 8�J�\�*��n��� ���������"��F� 4�j�X���|������� ������0@B T�x�d���� �>,Ntb ������/� (//8/:/L/�/p/�/ �/�/�/�/�/�/$?? H?6?l?Z?�?~?�?�? �?�?�?O�&O8OVO hOzO�?�O�O�O�O�O �O
__�O@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<o^o�oro �o�o�o�o�o�o  J8n$O��� ��X���4�"��X�B�v��$TBC�SG_GRP 2��B�� � �v� 
 ?�  ������׏ �������1��U�g��z���ƈ�d,� ���?v�	 H�C��d�>�����e�CL  B�p��Пܘ������\)��Y  A��ܟ$�B�g�B�Bl�i�X�ɼ���X��  D	J���r�����C����үܬ	���D�@v�=�W�j� }�H�Z���ſ���������v�	�V3.00��	�m61c�	*`X�P�u�g�p�>���2v�(:�� ��p���  O�����p�����z�JCFG� �B��� �����������=��=�c�q� K�qߗ߂߻ߦ����� ���'��$�]�H�� l������������ #��G�2�k�V���z� ������������ �p*<N���l� ������#5 GY}h��� �v�b��>�// / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?d? R?t?v?�?�?�?�?�? O�?*OO:O`ONO�O rO�O�O��O�O�O_ &__J_8_n_\_�_�_ �_�_�_�_�_�_�_o Fo4ojo|o�o�oZo�o �o�o�o�o�oB0 fT�x���� ���,��P�>�`� b�t�����Ώ����� ��&�L��Od�v��� 2�����ȟʟܟ� � 6�$�Z�l�~���N��� ��دƯ�� �2�� B�h�V���z�����Կ ¿����.��R�@� v�dϚψϪ��Ͼ��� ����<�*�L�N�`� �߄ߺߨ����ߚ�� �����\�J��n�� ���������"��� 2�X�F�|�j������� ��������.T Bxf����� ��>,bP �t�����/ �(//8/:/L/�/�� �/�/�/h/�/�/�/$? ?H?6?l?Z?�?�?�? �?�?�?�?O�?ODO VOhO"O4O�O�O�O�O �O�O
_�O_@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<oro`o �o�o�o�o�o�o�o &�/>P�/�� �������4� F�X��(���|����� ֏����Ə0��@� B�T���x�����ҟ�� ����,��P�>�t� b������������� ��:�(�^�L�n��� ����2d�����̿ �$�Z�H�~�lϢϐ� �������Ϻ� ��0� 2�D�zߌߞ߰�j��� �������
�,�.�@� v�d��������� ����<�*�`�N��� r������������� &J\�t�� B������ F4j|��^����/�  2 6# 6&J/6"��$TBJOP_�GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� ƞ6$ @2 �"	� �C�� �&b�  Cق'�!�!>ǌ��
559>��0+1�33=��CL� fff?>+0?�ffB� J1��%Y?d7�.��/>;��2\)?0��5���;��h{CY� �  @� ~�!B�  A�P?��?�3EC�  D��!�,�0*BO���?�3JB��
:�/��Bl�0��0�$��1�?O6!Aə�3AДC�1D�G6Ǌ=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__<�O�O>B�\JU�O�HH�1ts�A@g33@?1� C�� ��@�_�_&_8_>��D�UV_0�LP�Q30O<{�zR� @�0 �V�P!o3o�_<oRifo Po^o�o�o�oRo�o�o �o�oM(�ol��p~��p4�6&��q5	V3.0}0�#m61c�$�*(��$1!6�A�� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�IR�CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;S@;Q�U�|8�`rz@/&�8�6&<��1��w�^$ESTPAR�S  *({ _#H�R��ABLE 1%�p+Z�6#|�Q�Q � 1�|�|�|��5'=!|�	|�
|��|�˕6!|�|�:|���RDI��z!ʟܟ� ��$���O������¯ԯ�����S��x# V���˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���U-����ĜP�9� K�]�o��-�?�Q�c��u���6�NUM  ��z!� �>  Ȑ����_CF�G �����!@�b IMEBF_T�T����x#��a�VE�R��b�w�a�R {1�p+
 (3�6"1 ��  6!�� �������� �9�$�:� H�Z�l�~���������@������^$��_���@x�
b MI_�CHANm� x� >kDBGLV;0o��x�a!n ETHE�RAD ?�
� �y�$"�\&�n ROUT��!�p*!*�SN�MASK�x#�255.h�fx�^$OOLOFS_�DI��[ՠ	OR�QCTRL � p+;/���/+/=/ O/a/s/�/�/�/�/�/���/�/�/!?��PE?_DETAI���PON_SVOF�F�33P_MON� �H�v�2-9S�TRTCHK ����42VTCOMPATa8�24�:0FPROG �%�%MULTIROBOTTOx!O06�PLAY���L:_INST_M�P GL7YDUS8���?�2LCK�LPKQUICKMEt ��O�2SCRE�@}�
tps�@�2�A�@�I��@_Y����9�	SR_GR�P 1�� ���\�l_zZg_@�_�_�_�_�_�^�^� oj�Q'ODo/ohoSe ��oo�o�o�o�o�o �o!WE{i�������	1234567�h�!���X�E1�V[�
 �}ipn�l/a�gen.htmno��������ȏ�~�Panel� setup̌}��?��0�B�T�f� ��񏞟��ԟ� ��o����@�R�d�v� �����#�Я���� �*���ϯůr����� ����̿C��g��&� 8�J�\�n�����϶� ��������uϣϙ�F� X�j�|ߎߠ����;� ������0�B��*N�UALRMb@G ?�� [��� ���������� ��%� C�I�z�m�������v�SEV  �����t�ECFG CՁ=]/BaA$�   B�/D
 ��/C�Wi{� ������4 PRց; �To�\o�I�6?K0(%����0���� �//;/&/L/q/\/`�/�/�/l�D ��Q�/I_�@HIS�T 1ׁ9  �(  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1 Ec0p?�?�?�?/C�� >?P=962 n?�?
OO.O�?�?�136c?|O�O�O�OAO SO�?�O__0_�O�O _Lu_�_�_�_:_�/�_ �_oo)o;o�__oqo �o�o�o�oHo�o�o%7I~��a81�o u������o� ��)�;�M��q��� ������ˏZ�l��� %�7�I�[������� ��ǟٟh����!�3� E�W����������ï կ�v���/�A�S� e�Pb������ѿ� �����+�=�O�a�s� ϗϩϻ�������� ��'�9�K�]�o߁�� �߷��������ߎ�#� 5�G�Y�k�}���� �����������1�C� U�g�y���v������� ����	�?Qc u��(���� )�M_q� ��6���// %/�I/[/m//�/�/ �/D/�/�/�/?!?3? �/W?i?{?�?�?�?�� ���?�?OO/OAOD? eOwO�O�O�O�ONO`O �O__+_=_O_�Os_ �_�_�_�_�_\_�_o o'o9oKo�_�_�o�o �o�o�o�ojo�o# 5GY�o}�������?��$UI�_PANEDAT�A 1������  	�}�0�B�T�f�x��� )����mt� ۏ����#�5���Y� @�}���v�����ן�� �����1��U�g�N�\����� �1�� Ïȯگ����"�u� F���X�|�������Ŀ ֿ=������0�T� ;�x�_ϜϮϕ��Ϲ� �����,ߟ�M�� j�o߁ߓߥ߷���� ��`��#�5�G�Y�k� �ߏ���������� ����C�*�g�y�`� ��������F�X�	 -?Qc����߫ ����~; "_F��|�� ���/�7/I/0/ m/�����/�/�/�/�/ �/P/!?3?�W?i?{? �?�?�??�?�?�?O �?/OOSOeOLO�OpO �O�O�O�O�O_z/�/ J?O_a_s_�_�_�_�O �_@?�_oo'o9oKo �_oo�oho�o�o�o�o �o�o�o#
GY@ }d��&_8_�� ��1�C��g��_�� ������ӏ���^�� �?�&�c�u�\����� ��ϟ���ڟ�)�� M�����������˯ ݯ0�����7�I�[� m����������ٿ� ҿ���3�E�,�i�P� �ϟφ��Ϫ���Z�l�}���1�C�U�g�y���)߰�#�������  ��$�6��Z�A�~� e�w��������� ��2��V�h�O������v�p��$UI_P�ANELINK �1�v� � �  ���}1234567890����	 -?G ���o�� ���a��#5G�	����p&���  R��� ��Z��$/6/H/ Z/l/~//�/�/�/�/ �/�/�/
?2?D?V?h? z??$?�?�?�?�?�? 
O�?.O@OROdOvO�O  O�O�O�O�O�O_�O �O<_N_`_r_�_�_�0,���_�X�_�_�_  o2ooVohoKo�ooo �o�o�o�o�o�o� �,>r}����� �������/� A�S�e�w�������� я���tv�z��� �=�O�a�s������� 0S��ӟ���	��-� ��Q�c�u�������:� ϯ����)���M� _�q���������H�ݿ ���%�7�ƿ[�m� ϑϣϵ�D������� �!�3�Eߴ_i�{�
 �߂����߸������ /��S�e�H���~� ��R~'�'�a��:� L�^�p����������� ���� ��6HZ l~���#�5�� � 2D��hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?�/�?�?�?�? �?�?m?OO&O8OJO \O�?�O�O�O�O�O�O �O[�_��4_F_)_j_ |___�_�_�_�_�_�_ o�_0ooTofo��o ��o��o�o�o ,>1bt��� �K����(�:� ���{O������ʏ ܏�uO�$�6�H�Z� l���������Ɵ؟� ���� �2�D�V�h�z� 	�����¯ԯ����� �.�@�R�d�v���� ����п���ϕ�*� <�N�`�rτ��O�Ϻ� Io���������8�J� -�n߀�cߤ߇����� �����o1�oX��o |����������� ��0�B�T�f���� ����������S�e�w� ,>Pbt��' �����: L^p��#�� �� //$/�H/Z/ l/~/�/�/1/�/�/�/ �/? ?�/D?V?h?z? �?�?�???�?�?�?
O O.O��ROdO�߈OkO �O�O�O�O�O�O_�O <_N_1_r_�_g_�_7O�M�m�$UI�_QUICKME�N  ���_AobRESTORE 1��  ��|��Rto�o�im �o�o�o�o�o: L^p�%��� ���o����Z� l�~�����E�Ə؏� ��� �ÏD�V�h�z� ��7�������/���
� �.�@��d�v����� ��O�Я�����ß ͯ7�I���m������� ̿޿����&�8�J� �nπϒϤ϶�a��� ����Y�"�4�F�X�j� ߎߠ߲������ߋ����0�B�T�gSC�RE`?#m�u1sco`uU2��3��4��5��6��7��8��bUGSERq�v��Tp঑�ks����4��5*��6��7��8��`�NDO_CFG ��#k  n` �`PDATE ����Non�ebSEUFRA_ME  �TA��n�RTOL_AB�RTy�l��ENB�����GRP 1��ci/aCz  A�����Q�� $�6HRd��`U������MSK  ������Nv�%��U�%���bVI�SCAND_MA�X�I��FAIL_IMG� ��PݗP#��IM�REGNUM�
�,[SIZ�n`��A�,VONT�MOU��@����2��a���a����F�R:\ � �MC:\�\wLOG�B@F� !�'/!+/O/�U�z MCV��8#UD1r&E�X{+�S�PPO�64_��0'f�n6PO��LI�b�*�#V���,�f@�'�/� =	��(SZV�.�����'WAI�/ST�AT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_�JMPERR 1��#k
  �23�45678901 dF�ψO{O�O�O�O�O �O_�O*__N_A_S_x�_
� MLOWc>8
 �_TI�=��'MPHASOE  ��F��P�SHIFT�15 9�]@<�\� Do�U#oIo�oYoko�o �o�o�o�o�o�o6 lCU�y�� ��� ��	�V�-��e2����	VSwFT1�2	V�M�� �5�1G� ����%A�  BU8̀̀�@ pك�Ӂ˂�у��z�ME�@�?�{��!c>&+%�aM1��k�0��{ �$`0TDI�NEND��\�O � �z����S��w���P���ϜRELE�Q��Y���\�?_ACTIV��<:�R�A ��e���e�:�RD� ���YBOX �9��د�6��02����190.0m.�83���254��QF�	� �X�j��1�robot����   px�૿�5pc�� ̿�����7�����-�^f�ZABC�����,]@U��2ʿ�eϢ� �ϛϭϿ����� �� �V�=�z�a�s߰�E�	Z��1�Ѧ