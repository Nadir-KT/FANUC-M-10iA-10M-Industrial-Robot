��   38�A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����UI_CON�FIG_T  �T ($NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$DU�MMY36CME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  u�7�ODE�
]8CFOCA ��9CPS)C��\g 
HAN� � �TIMEOU�P�IPESIZE �� MWIN�P�ANEMAP� � � NU_FA�VB ?� 
$H�LP> _DIQ?y� mELEMVF}UR� h� So��$HMI�R�O'XW ADO�NLY� �TOwUCH�PROoOMMO?$��ALAR< �FI�LVEW�ENAB=!%bC -"�USER6)FCT�N6)WI�� I�* _ED�h"R!_�TITL�  �&USTOM0� t $} RT�_SPID��$Cܨ$*PAG� ?~ZDEVICE�)oSCREqEF����'N�@$FL�AG�@ �"US�RVI 1  < \� +2�n,1PRI�m� yA� K0TRIP�"�m�$$CLAS�S  ����l1��R��Ra0VI�RTO1j?|0'2 )��E�)�O`�R	 /�,��;����2�0�3�3�1��� , � � �?��
 ��s1,O>OPObOtO�O�O (O�O�O�O�O_ _�O;_M___q_�_�_ $_�_�_�_�_oo%o �_Io[omoo�o�o2o �o�o�o�o!�oE Wi{���@� ����/��S�e� w�������<�я������+�=� /TPTX��͈`��r�  sH����$/softpa�rt/genli�nk?help=�/md/tpmenu.dg?�ٟ� ���ȏ3�E�W�i�{� �����ïկ���� ���A�S�e�w����� *���ѿ�������+9���F�6�3C�($��p���^ϗ��ϻ���s1�1���?�K������̛3�" �1�5�2 \��6 RE�C VED��U�g��wholemod�.htm{�sin�gl��doub~��trip��brows�� ��h�
��.���R�d� v�����R�<�v߈�_dev.s��l�4��(�1�	t?��� (����������|��������G�  �0_q����� ��0\1C gy��I�B< ����//*/</ N/`/r/�/�/�/�/�/ �/�/?��??B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �OT�O�O�O�O	__ -_?_Q_c_^�_�_h_ z_�_�_���O)o$o 6oHoqolo~o�o�o�o �o�o�o ID V$?vp���� ��
��.�@�R�d� v���������Џ⏰O �/�A�S�e�w����� �����_���ğ֟+� =��_o쏅������� ͯȯگ���"�4� ]�X�j�|�������� ҿ̿����0�B�T� f�xϊϜϮ������� ����,�>��yߋ� �߯���������	�� �?�Q� �2���P� b�H������� �)�$� 6�H�q�l�~������� ������ܿ.( Vhz����� ��
.@Rd v��h����/ ///A/S/e/w/r�/��/|/�/�/�/:�$�UI_USERV�IEW 1���R 
�A��6?H?�mg? �?�?�?�?�?{?�?O  O2ODO�?hOzO�O�O �O[?�O�O�OSO_._ @_R_d__�_�_�_�_ �_�_�_oo*o<oNo �O[omoo�_�o�o�o �o�o&8J\n ������o� ��}/�X�j�|��� ��C�ď֏������ 0�B�T�f�x�#����� ��������,�ϟ P�b�t�������M�ί ������#�5�G� ����������ʿm��  ��$�6�ٿZ�l�~� �Ϣ�M�W�����E���  �2�D�V�h�ߌߞ� ������w���
��.� @���M�_�q��߬�� ��������*�<�N� `�r������������ ��������J\n ��5����� �"4FXj �����// 0/�T/f/x/�/�/?/ �/�/�/�/?�(