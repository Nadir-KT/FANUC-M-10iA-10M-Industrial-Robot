��   �A��*SYST�EM*��V7.5�0130 3/�19/2015 �A ���$$�CLASS  O���(��D���D VIRTUA�L%7MNUFR�AME AF�D� �� 	 88�?���}��y�� ����1= gQs�������	/�/?/��WN_UM  ��>l� ontWTOO=La4 
wY/ �/5/�/�/�/?5?? A?k?U?w?�?�?�?�? �?�?O�?	OCO-O?O aOcOuO�O�Om&�!{&����&�a