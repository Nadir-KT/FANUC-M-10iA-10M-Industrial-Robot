��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5M�AUTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{� �BL� OU&R ,A�0�!z� B� LM_O�z
eR�"CAM_;�1 xr$�ATTR4�@� A�NNN@5IMG_�HEIGH�AXcWoIDTH4VT� ��UU0F_ASP�EC�A$M�0E�XP�.@AX�f��CF�D X '$GR� � S�!.@=B�PNFLI�`�d� UIRE 3T!GOITCH+C�`N� MS�d_LZ`AC�"��`EDp�dL� J�4S�0� <za�!p�;G0 � 
?$WARNM�0f�!�@� -s�pNST�� CORN�"a1F�LTR{uTRAT�� T}p  $ACCa1�p��|{��rORI�P�C�kR�T0_S~B\qHG�,I1 [ Th�`�"3I�pTYD(�@*2 3`#@� X�!�B*HDDcJ* TCd�2_�3_�4_�U5_�6_�7_�8_��94FCO�$ <� �o�o�hK3 1#`�O_Mc@AC t� � E#6NGPvABA� �c1�Q 8��`,��@nr1��� d�P�0e���axnpUP&Pb26��4�p�"J�p_R�rPB�C��J�rĘߜJV �@U� B��s}�g1�"vYtP_*0OFS&Rw @� RO_K8�T��aIT�3T�NOM_�0�1p�34 >��D �� Ќ@�2�hPV��mEX�p� Ĝ0g0ۤ�p�r
$�TF�2C$MD3&i�TO�3�0U� F�/ ��Hw2tC%1(�Ez�g0#E{"F�"F�>�@�a�2 �@$�PPU8�3N)ύR&ևAX�!DU��;AI�3BUF�F=�@1 |pp���pkPIT� PP�EM�M�y��F�SIMQSI�"ܢ8VAڤT�)?�w' T�`(zM��P��B�qFACTb�@EW�P1�BTu�A?�MC� �$*1JB`p�*1DEC��F��ŏ��� �H0CHN�S_EMP1�$G��8��@_4�3�p2|@P��3�TCc�(r /�0-sx��ܐ� MB0i��!����JR� i�_SEGFR��Iv *�aR�TpN�C���PVF��?�bx &��f{uJc!� Ja��� !28�ץ�AJ���SIZ�3S�c�B��TM���g��JaRSINFȑb���q�� ��н����L�3��B���CRC�e�3CCp����c��mc� �b�1J�cѿ�.����D$ICb�Cq�5r��`���@v�'���EV����zF��_��F,pN��ܫ�?�4�0A�! �r���h�� ���p�2�͕a�� ��د\qR�Dx Ϗ��o"27��!ARV�O`C�$L	G�pV�B�1�P��@��t�aA�0'�|�+0Ro�� MEp`"1 �CRA 3 AZ�V�g6p�O �FCCb�`�`F�`K������ADI��a�A �bA'�.p��p�`�c¢`S4PƑ�a�AMP$��-`Y�3P�M�r��UR��QUA1  $.@TITO1/S@S��!����"0�DBP�XWO��B0!5��$SK���2�DBdq�!"�"�PR��? 
C�D=���΁!# S q1$�2�$z���L�)$$�/Xr��� %�/�$�C�!&?�$ENE��q.'*?�#� R�E�p2(H z��O�0#$L|3$$�#�B[�;���F�O_D��RO�Sr�#������3R�IGGER�6PA�pS����ETURN��2�cMR_8�TUrw��0EWM�ҍM�GN�P���BL�AH�<E���P��'&$P� �'P@�Q"3�CkD{��DQ���4�11��FGO_A7WAY�BMO�ѱQ�#!�DCS_޾)  �PIS � I gb {s�C��A��[ �B$�S��A�bP�@�EW-�TNT	Vճ�BV�Q.�C�(c`�UWr�P�J��P�$0���SAFE���V_�SV�bEXCLUt��nONL2�b�SY�*a&�OT�a'�HI_V�4��B<���_ *P0� r9�_z��p �"v�@SG�� +nr r�@6Acc*b��G�#@�E�V.iHb?fANNcUN$0.$fdID�	U�2�SC@�`�i�ax��j�f����z���@I$2,O�$F�ibW$}�OT9@�1� $DUMMY T��da��dn�� � ��E- ` ͑HE4(sg�*b�SAB���SUFFIW�V�@CA=�c5�gu6r� MSW�E�. 8Q�KEYI5���TM�10s�qA&�vIN����D���/ D��HOST_P!�rT��ta��t0n��tsp�pEMӰV���� SBLc UL>I�0  8	=�ȳ���DTk0�!1� � $S��ESAMPL��j�۰f爒�f���I�0��[ $SUB�k�#0�Cp��T�r#a�SAVʅ ��c���C��P�f�P$n0E�w YN�_B#2 0Q�D�I{dlpO(��9#�$�R_I�� �ENC2_S� 3  5�C߰�f�- �SpU����!!4�"g�޲�1T���5X�j`ȷg��0��0K�4�AaŔAV�ER�qĕ9g�DSP�v��PC��r"�(���ƓVALU�ߗHE�ԕM+�I�Pճ��OPP ���TH��֤��P�SH� �۰F��df��J� �ѸC1+6� H�bLL_DU s�~a3@{��3:����OTX"���sȣR_NOAUTO�!7�p$)�$�*��c�4�(�C� 8�C�, �"�!&�L�� �8H *8�L H <6����c"�`,  `Ĭ�kª�q��q��Psq��~q��7��8���9��0����1��1�̺1ٺ1�1�1� �1�1�2(�2T����2̺2ٺ2�U2�2 �2�2ʕ3(�3��3��̺3�ٺ3�3�3 �3��3�4(��(q���?��!9 <�9�&�z��I��1��׌M��QFE@'@� :� ,6��Q? ��@P?9��5�9�E�@A�!�A� �;p$TP�$VARI:�Z���7UP2�P< ���TDe���K`Q��r����Ќ�BAC�"G= T�p��e$)_,p�bn�kp+ IFIG� kp�H  ��P�Ȣ�F@`�!>t �;E��sC�ST �D� D���c�<�� 	C��{��_����l���R  ���FO�RCEUP?b��FWLUS�`H�N>�xF ���RD_CM�@E������ ��@vMP.��REMr F�Q��@1k@���7Q
K4	9NJ�5EFFۓ:f�@IN2Q��OVO�OVA�	TRO�V���DTՀ�DTMX� ��@�
�ے_PH"p��CL��_TpE�@�pK	_(�Y_T��v(���@A;QD� �������!0tܑ0R�Q���_�a����M̝7�CL�dρRIqV'�{��EARۑIOHPC�@����B�B��CM9@���R{ �GCLF��e!DYk(M�ap#5TuDG��� �%���SSD �s? PP�a�!�1���P_�!��(�!1��E�3�!3z�+5�&�GRA��J7�@��;�PW���ONn��EBUG�_SD2HP�{�_E� A`�=��/TERM`5Bi5K@O�ORI#e0Ci5�{�SM_�PԌ�e0Di5Ң0TAڧ9E�9UP\�Fg� -�A{�AdP|w3S@B$SEG�:v� EL{UUSE�@NFIJ�B$�;1x젎4�4C$UFlP=�$,�|QR@��_G90Tk�D�~SwNST�PAT��<��APTHJ3Q�E�p%B`�'EC����AR$P�I�aS�HFTy�A�A�H_�SHORР꣦6 ��0$�7PE��E�O#VR=��aPI�@��U�b �QAYLOW���IE"�r�A��?���ERV��XQ� Y��mG>@�BN��U�\��R2!P.uAScYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC���EaP;�uP;�6WOR>@�M`�!�GRSMT6�G3�GR��13�a�PAL@��P��q�uH� � ���T�OCA�`P	P�`$OP����p�ѡ��`0O��RE�`R4C�AO�p낎Be�`R�Eu�h�A���e$PWR�IMu�RR_�cN��q.=B I&2H���p�_ADDR��H_LENG�B�q�q�q�$�R��S�JڢSS��SKN��u\��u̳�uٳSE�A�jrmS��MN�!K������b����OL�X��p����`ACRO3pJ�@��X�+�p�Q��6�OUP3��b_�IX��a�a1 ��}򚃳���(��H ��D��ٰ��氋�+IO2S�D���x��	�7�L $l�<�`Y!_OFFr�oPRM_�����_HTTP_+�H:�wM (|pOBJ]"l�p��$��LE~C�d���N � \��֑AB_�Tq�b��S�`H�LVh��KR"uHITC�OU��BG�LO�q���h�����`���`SS� ���HQW�#A:�Oڠ<`�INCPU2VISIOW�͑��n��t�o��to�ٲ �IO�LN��P 8��R���p$SLob� PUT_n�$�p��P& ¢��Y F�_AS�"Q��$AL������Q  U�0�	P4A��^���ZPH�Y��-��p�UOI �#R `�K���@�$�u�"pP�pk���$�����q1UeJ5�S-���NE6W�JOGKG̲DISĖ��Kp���#T �(�uAVF�+`�CTyR�C
�FLAG2v�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w� m� _�{0a�^��cg���4� ����Ǝ���{0��� �SCH_���a7�NT�d�VW���E�"����4��UM�Aљ`�LJ�@�DAUf�E�AU�p��d|�r�GH��b/���BOO��W�L ?�6 ITp��y0�REC��GSCR ܓ�D
�<\���MARGm�!���զ ��d%�����S�����W���U� �J{GM[�MNCHJ���FNKEY\�Kn��PRG��UF���7P��FWD��HL.��STP��V��=@X��А�RS��HO`����C9T��b ��7�[�UL���6�(RD�� ����Gt��@POЛ�������MD�FO{CU��RGEX���TUI��I��4� @�L�����P@����`��P��NE���CANA��Bj�V7AILI�CL !�U?DCS_HII4�D�s�O�(!�S�$��S��� ���BUFF�!X�?PTH$m���vP`�ěԬ�AtrY��?P��j�3��`OS1Z2Z3Z�@�|�� Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�C���K�&&8���![ LQ��+00� 	P���`#qdt
�U�dw�<���_ \ ��`4Г�\��Ѩ#��MC4�] ��C�LDPL��UTRQ�LI��dڰ�)�$F�LG&�� 1�#�D���'B�LD�%�$�%ORGڰ5�2�PV� �VY8�s�T�r �#}d^ ���$6��$�%�S�`T� �B0�4>�6RCLMC�4]?0o?�9�9MI�p}dg_ d=њRQ�=�DSTB�p�c ;F�HHAX�R� JHdLEXCE�SryBM!p�a`���/B�T�F��`a�p=F_A7Ji��K�bOtH�0K�db \�Q���v$MBC�L�I|�)SREQUI�R�R�a.\o�AXDE�BUZ� �ML
t M��c�b�{P��4��2ANDRѧ``d;�2�ȺSDC��N�INl�K�x`찄�X� N&��aZ���UPST� enzrLOC�RIrp�EX<fA�p�9A�AODAQ��f �XY�OND�rMF ,Łf�s"��}%�e�/� �8FX3@IG}G�� g ��@t"��ܓs#N�s$R�a%��iL��hL�v<�@�DATA#?pAE�%����Y�N�h t $MD
`qI}�)nv� ytq�ytHP`�Pxu��(�zsANSW)�yt@��
yuD+�)\b���0o��i �@CUw�V��p 0XeRR2��j� Du�{Q��7Bd$OCALIA@��G�:�2��RIN��"�=<9INTE��C�k�r^�آXb]���_N�qlk���9�D����Bm��DIVFD�H�@���qnI$�V,��S�$���$Z�X�o�*�����oH �$�BELT�u!ACCEL�.�~�=��IRC�� ���D�T<�8�$PS�@�"L�@�r��#^�S�xEы T�PATH3����I���3x�p�A_@W��ڐ���2nC���4�_MG�$D�D��T���$FW��Rp9��I�4��D}E7�PPABN��ROTSPEE�[g�� J��[�C@�4��@$USE_d+�VPi��SYY����1 �aYN!@A��ǦOFF�qǡM�OU��NG���O9L����INC�tMa�6��HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]�ౌB��VE��#�y�2�3_UP񕋳LOWL���p� B���Du�9B#P`�x ����BCv�r�MOSI���BMOU��@�7P�ERCH  ȳOV��â
ǝ���� D�ScF�@MP����B� Vݡ�@y�j�LU0k��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A���x�����N`�F�RT1I�A$��MOUІЀHB�BS0�p7D5����ë�Z�DUM2�ԓS_BCKLSH_Cx�k���� ϣ���=���ޡ ��1CLAL"q��1М�@��CHK� �S�RTY��^�%�E1Qq_�޴_UM��@�C#��SCL�0�r�LMT_J1_L��9@H�qU�EO�p�b�_�e�k�e�SPC��u���N�PC�N�Hz \P�2�C�0~"XT��CN_:�N9��I�SF!�?�V���U� /���x�T���CB!�SH�:��E�E1TрT����y���T��P�A ��_P��_ � =������!�����J6 L�@��OG|�G�TORQU��ONֹ��E�R��H�LE�g_W2���_郠����I�IJ�I��Ff`xJ�1X�~1�VC3�0BD:B�1�@SB�JRKF9�0D�BL_SM��2M��P_DL2GR�V����fH�_��d���COS���LNH� �������!*,��aZ���fMY��_(�TH��)T�HET0��NK2a3���"��CB�&CB�CAA�B�"�0�!��!�&SB� 2N�%GTS�Ar�CI Ma�����,4#97#$DU���H\1�  �:Bk62�:AQ(rSf'$NE�D�`I��HB+5��$̀�!A�%��5�7���LPH�E�2���2SC% C%�2-&FC0JM&̀EV�8V�8߀LVJUV!KV/KV=KVKKVYKVgIH�8FRPM��#X!KH/KH=KUHKKHYKHgIO�<�O�8O�YNOJO�!KO/KO=KOKKO
YKOM&F�2�!+i%�0d�7SPBALA�NCE_o![cLE60H_�%SPc� &��b&�b&PFUL�C�h�b�g�b%p�1=k%�UTO_���T1T2�i/�2N ��"�{�t#�Ѱ`�0(�*�.�T��OÀ<�>v INSEG"�ͱ�REV4vͰl�DI�F�ŕ�1lzw��1m��OBpq�я?��MI{���nLCHgWARY�_�AB��~!�$MECH�!�o ��q�AX��P�����7Ђ�`n 
p�d(�U�ROB���CRr�H����(��MSK_f`�p� P �`_��R /�k�z�����1S�~��|�z�{���z��qIN�Uq�MTCOM�_C� �q  ����pO�$NO�REn����pЂ7r 8p GRe�u�SD�0AB�$?XYZ_DA�1a���DEBUUq�������s z`$��COD�� L���p��$BUFIwNDX|�  <��MORm�t $فUA��֐����r�<��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p} =�C�}pt�@b�D��FRIrӚ�T��RO@ \�E�}�����OPWO�Yq�v0Y�SY�SBU/@v�$SO!Pġd���ϪUΫ}p�PRUN����PA�D���rɡL�_O�Uo顢q�$^)�IMAG��w���0P_qIM��L�I�Nv�K�RGOVCRDt��X�(�P*�J�|��0L_�`]�L�0�RB1�0��M��ED}��p J��N�PMֲ��c��w�SL�`q�w x $OVSL4vwSDI��DEX�@���#���-�V} *�N4�\#�B�2�G�4B�_�M�y�q|�E� x Hw���p��ATUSW����C�0o�s���BT�M�ǌ�I�k�4p��x�԰q�y Dw�!E&���@E�r��p7��жЗ�EXE���ἱ�����f q�z3 @w���UP'��3$�pQ�XN����������� �PG�΅{ h $S#UB����0_���!��MPWAIv�PL7ã�LOR�٠F\p�˕$RCVFA�IL_C��٠BW�D΁�v�DEFS}P!p | Lw����Я�\���UN!I+�����H�R�+�}_L\pP��x�t���p�}H�> �*�j��(�s`~�N�`KET�B�%�J�PE Ѓ~z��J0SIZE�����X�'���S�OR~��FORMAT�``��c ��WrEM�t��%�UX��G�G��LI��p�  �$ˀP_SWIp�p{��J_PL��?AL_ ����ХA��B��� C��Dn�$E��.��C_�U�� �� � ���*�J�3K0����TIA4��5��6��MOM���������ˀB��AD����������PU� NR�������u��m��� A$PI�6q��	 �����K4�)6��U��w`��SPEEDgPG������ ��Ի�4T�� �p @��SAMr`���\�]��MOV _�_$�npt5��5���1���2���������'�S�Hp�IN�'�@�+�����4($4+T+GAM�MWf�1'�$GE�T`�p���Da���
�
pLIBR>�II.2�$HI=�_g�t�$�2�&E;��(A�.� �&LW�-6<�)56��&]��v�p��V��$PDCK��D�q��_?����� q�&���7��4���9�+� �$IM_SR�pD�s�rF�L�r�rLE���Om0H]��0���pq���PJqUR_S�CRN�FA���S_?SAVE_D��dE@�NOa�CAA�b� d@�$q�Z�Iǡs	�I � �J�K� ����H� L��>�"hq��� ���ɢ�� bW^U�S�A���M4� ��a��)q`��3�WW� I@v�_�q���MUAo��� � $PY�+�$W�P�vNG�{��P:��RA��RH��RO�PL�����qP� ��s'�X;�OI��&�Zxe ���m�� p��ˀ�3s�O�O��O�O�O�aa�_т� |��q�d@��.v��.v��d@��[wFv��E����%s�t;B�w�t|�tP���PMA��QUa ��Q�8��1٠QTH�H{OLW�QHYS��3ES��qUE�pZB���Oτ�  ـP�ܐ(�A����v�!�t�O`�q��u�"���8FA��IROG�����Q2���o�"��p�^�INFOҁ�׃hV����R�H�OI���� (�0SLEQ ������Y�3����Á��P0Ow0��5�!E0NU���AUT�A�COPAY�=�/�'��@Mg��N��=�}1������ ���RG��Á���X_�P�$;ख�`
��W��P��@��������EXT_CY�C bHᝡRpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�H�SdB����2�$��F�p���GPLeAdA
�TAR �Б@���P�2��裔d� ,�0FL�`�o@YN��K�Mz��Ck��PWR+��9ᘐ��DELA�}�dY�pAD�a�u�QSKIP4�� �A�$�OB`NT2�} ��P_$�M� ƷF@\bIpݷ�ݷ� ݷd����빸��Š��Ҡ�ߠ�9���J2R� ��� 46V�EX� TQQ�� ��TQ������ ��`��H�RDC�V� �`��X)�R�p������r��m$RGEA�R_� IOBT�2FcLG��fipER��DTC���Ԍ���2T�H2NS}� 1����G T\0 ����u�M\Ѫ`I��dG�REF�1�Á� l�h��ENsAB��cTPE�0 4�]����Y�]��ъQ n#��*��"�������2�Қ�߼���������3�қ'�9�K�P]�o���4�Ҝ��@�����������5���!�3�E�W�i�{��6�Ҟ�������������7�ҟ-?PQcu�8�Ҡ��������SM+SKÁ�l��a���EkA0��MOT-E6�����@��݂TQ�IO}5�I8STP��POW@��� �pJ����p�����E�"$DS?B_SIGN�1UQ��x�C\��S23�2���R�iDEVICEUS�XRSR�PARIT��4!O�PBIT�QI�O?WCONTR+�TQX��?SRCU� MpS�UXTASK�3Nx�p�0p$TATU�P#E#�0�����p�_XPC)�$FREEFROMS	p�na�GET�0��U�PD�A�2��RS�P� :��� !>$USAN�na8&����ERI�0�&RpRYq5*"_j@�qPm1�!�6WRK9�KD���6��QFR�IEND�Q�RUFxg�҃�0TOOL�6�MY�t$LEN�GTH_VT\�FCIR�pC�@ˀE> �+IUFIN-RM�ΕRGI�1ÐAITI�$GXñ3IvFG2v7G1���p3��B�GPR�p�1F�Oa_n 0��!RE��0p�53҅U�TC��3A�A�F �G(��":���e1n!��J�8 �%���%]��%�� 74��X O0�L
��T�3H&��8���%�b453GE�W�0�WsR�TD����T��M�����Q�T]�$V �2����1�а91T�8�02�;2k3�;3�:ifa�9-i�aQ0��NS��ZR$V��2B�VwEV�	V�B;�����&�S�`��F�"��k�@�2a�PS�E���$r1C��_3$Aܠ6wPR��7vMU�cS�t '�/89�G� 0G�aV`��p�d`���50�@��-��
25S�� �"�aRW����B�&�MN�AX�!�A:@�LAh��rTHIC¤1I���X�d1TF�Ej��q�uIF_C	H�3�qI܇7�Q�pG1RxV���]��:��u�_JF~�PR|ԀƱ�RVAT��� ��`���0R�榀DOfE��COU�Ա��AXI���O�FFSE׆TRIGNS���c����h������H�Y��IG#MA0PA�pJ�E��ORG_UNEV��J� �S������d �$CА��J�GROU����TqOށ�!��DSP���JOGӐ�#��_Pӱ�"O�q����@�&7KEP�IR��ܔ2�@M}R��AP�Q^��Eh0��K�SYS��q"K�PG2�BRAK�B��߄�pY�0=�d����`AD_������BSOC���N���DUMMY14�p@SV�PDE_�OP�#SFSPD�_OVR-���C���ˢΓOR٧3N�]0ڦF�ڦ��OV���SF��p���F�+�r!���CC��1q"L�CHDL��REC�OVʤc0��Wq@M������RO�#��Ȑ9_+��� @0�e@�VER�$OF�Se@CV/ �2WD��}��Z2���T�R�!���E_F�DO�MB_CM4���B��BL�bܒ#��adtVQR�$0pd���G$�7�AM5�`�� eŤ��_M;��"'����8$CA�'�E�8�8$HB�K(1���IO<�8����QPPA�������
��Ŋ����DVC_DBhC;��#"<Ѝ�r!S�1[ڤ�S�y3[֪�ATIOq 1q� ʡU�3���CABŐ�2�CvP���9P^�B���_� �S�UBCPU�ƐS �P �M�)0NS�c�M�"r�$HW_AC��U��S@��SA�A~�pl$UNITm�l_�AT���e�Ɛ�CYCLq�NEC�A���FLTR_2_FIO�7(��)&�B�LPқ/�.�_S[CT�CF_`�Fb�l���|�FS(!E�e�CHA�1��4�D°"3�RSD��$"}�����_Tb�PROX����� EMi_��ra�8!�a !�̹a��DIR0�RAOILACI�)RMr�CLO��C���Qq���#q�դ�PR=�S��AC/�c 	���FUNCq�0rRINP�Q�0��2�!3RAC �B ��[8���[WARn���#BL�Aq�A�����DAk�\���LD0���Q��q2eq�TI"r8��K�hPRIA�!r"AF��Pz!=�;���?,`�RK���MǀI�!�DF_@B�%1�n�LM�FAq@H�RDY�4_�P@R�S�A�0� �MUL�SE@���a ���ưt��m�m$�1$�1$1�o����� x*�EG� ����!cAR���Ӧ�09�2�,%� 7�AXE��RKOB��WpA��_l-���SY[�W!‎&S&�'WRU�/-1��@��STR������Eb� 	�%��J��A�B� ���&9�����O�To0 	$��A�RY�s#2��Ԓ�	�ёFI@��$LGINK|�qC1�aI_�#���%kqj2XYZ��t;rq�3�RC1j2^8'0B���'�4����+ �3FI���7�q����'���_Jˑ���O3�QO�P_�$;5���AT�BA�QBC��&�D�Uβ�&6��TURN߁"r�E11:�p��9GFL�`_���* �@�5�*7��Ʊ 1��� KŐM��&8����"r��ORQ ��a�(@#p=�j��g�#qXU�����mTOVEtQ:�M��i�� �U��U��VW�Z�A �Wb��T{�, ��@;� uQ���P\�i��UuQ�W`e�e�SERʑ
e	��E� O���UdAas��4S�/7����AX��B�'q ��E1�e��i��irp �jJ@�j�@�j�@�jP �j@ �j�!�f��i� �i��i��i��i� y�y�'y�7yTq�HyDEBU8�$ 32���qͲf2G �+ AB����رnSVS�7� 
#�d�� L�#�L��1W��1W�JA W��AW��AW�QW�@!�E@?D2�3LAB��29U4�Aӏ��C 7 o�ERf�5�� � $�@_ A6��!�PO��à��0#�
�_MRA�t�� d � T��ٔERR����;STY&���I��V�0��cz�TOQ�d�PL [ �d�"�� ?�w�!_ � pp`T)0���_V1Vr�aӔ����2ٛ2�E�����@�H�E���$W������V!��$�P��o�cI��aΣ�	 HELL_C�FG!� 5���B_BASq�SqR3��� a#QSb���1�%��U2��3��4��5���6��7��8���RaO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CO,. U�OUG�P~ ��`��m�������TPհ�_KAR�l�_�R�E*��P���7Q�UE���uP����C�STOPI_AL 7�l�k0��h��]�l0GSEM�4�(�M4�66�TYN�SO���DIZ�~�A�����m�_TM�MANR�Q��k0E����$�KEYSWITCaH���m���HE��OBEAT��E- �LE~�����U��F�!Ĳ���B�O_HOuM=OGREFUP�PR&��y!� [�Cr��O��-ECOC�|�Ԯ0_IOCMWD<
�a��(k���� � Dh1���U�X���M�βgPgCFgORC��� ���m�OM.  � Q@�5(�U�#P, Q1��, 3��45~��NPX_ASt�w� 0��ADD�о�$SIZ���$VAR���TI�P/�.��A�ҹ�M�ǐ��/�1�+ U"S��U!Cz���FRI	F��J�S���5Ԓ��NF�� �� � mxp`SI��TE�C\���CSGL��TQ2��@&����� ��S'TMT��,�P �&�BWuP��SHOW�4���SV�$��� �Q�A00 �@Ma}���� ��ਅ�&���5��6��7*��8��9��A��O ����Ѕ�Ӂ���0��F ��� G��0G���0 G���@G��PG��U1	1	1	1+	U18	1E	2��2��U2��2��2��2��U2��2��2��2��U2	2	2	2+	U28	2E	3��3��U3��3��3��3��U3��3��3��3��U3	3	3	3+	U38	3E	4�4��U4��4��4��4��U4��4��4��4��U4	4	4	4+	U48	4E	5�5��U5��5��5��5��U5��5��5��5��U5	5	5	5+	U58	5E	6�6��U6��6��6��6��U6��6��6��6��U6	6	6	6+	U68	6E	7�7��U7��7��7��7��U7��7��7��7��U7	7	7	7+	e78	7E��VP���UPDs�  ��`NЦ�5�YSL}Ot�� � L�`��d���A�aTA�80d��|�ALU:ed��~�CUѰjgF!aIgD_L�ÑeHI�j�I��$FILE_X���d��$2�Ue;SA>�� hO��`?E_BLCK��b|$��hD_CPUy�M�yA��c�o�d��Y�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA�i�J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP��_(�g����pr��� `�`GROU�w`��B��NFL�IC��f�REQUwIRE3�EBU�0�qB���w�2����p����q5�p�� \^��APPR��C}��Y�
ްEN٨CL9O7��S_M��H����u�
�qu�� ���MC�����9�'_MG��C�Co��`pM�в�N�BRKL�GNOL|�N�[�R���_LINђ�|�=�J����Pܔ�������� ���������6ɵ�̲8k�{���q��ď� ��
��qx)��7�PATH3ǀL�B�L��H�wࡠ�6J�CN�CA�Ғ�lڢB�IN�rUCV��4a��C!�UM��Y,���aE�p�����ʴ���PAYLO�A��J2L`R_AN�q�Lpp����$�M�R_F2LgSHR��N�LO���Rׯ�`ׯ�ACRL_G�ŒЛ� ��9Hj`߂$HM��үFLEXܣ�qJ>�u� :�� �����������1�F1�V�j�@�R� d�v�������E���� ȏڏ����"�4�q� ��6�M���~��U�g�Hy�ယT��o�X�� H������藕?��� ��ǟِݕ�ԕ�����%�7��JJ�� � V�h�z���`cAT�採@�EL��S S��J|�Ŝ�;JEy�CTR��~��TN��FQ��HA_ND_VB-����v`�� $��F20M����ebSW�rD��'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aDM)F�AW�Z`i�Aw�AA��X X�'pi�Dw��D��Pf�G�p�)S�Tk��!x��!N��DY�pנM�9$`%Ц� H��H�c�׎���0� ��Pѵڵ���������D�J��� ���1��R�6��QOASYMvř����v��J���cі�_SH>��ǺĤ�ED����������J�İ%�p�C�IDِ�_VI��!X�2PV_UN!IX�FThP�J��_R �5_Rc�cTz�pT�V�݀@���İ�߷��U $����D���Hqpˢ3��aEN�3�SDI����O4dD��`J�� x g"IJAAȱz�aabp�coc��`a�pdq�a� �^�OMME��� h�b�RqT(`PT�@ � S��a7�;�Ƞ�@ȷh�a�iT�@<� �$DUMMY9�Q�$PS_��R�FC��$v �����Pa� XXƠ���STE����SBRY�M21_�VF�8$SV_E�RF�O��LsdsCLRJtA��Odb`�O�p � D ?$GLOBj�_LO���u�q�cAp�rܛ@aSYS�qADqR``�`TCH  � ,��ɩb�oW_NA����7���TSR���l ���
* ?�&Q�0"?�;'?�I) ?�Y)��X���h���x� �����)��Ռ�Ӷ�;� �Ív�?��O�O�O�D>D�XSCRE栘p5����ST��s#}y`���Ea/u_HA�q� TơgpTYP�b���PG�aG���Od0�IS_䓀eАUEMd� ����ppyS�qaRSM_�q�*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCO�U��S�Ԕ 1�!�UE&��Ubwr���PROGM�FL�@$CUgpPOX�Q��5�I_�`H�� � 8�� �_�HE�PS�#��`RY ?�qp�b�t�dp�OUS��� � @6p�v_$BUTTp�Rp>R�COLUMq�e���SERV5�P�ANEH�q� �; �@GEU����Fy��)$HELyPõ)BETERv�)ෆ���A � � ��0��0��0ҰSIN簪c�@N���IH�1��_� �֪�LN�rؓ �qpձ_ò=�s$H��TEXl�����FLA@��RELV��D`����j����M��?,�Š��m����"�U�SRVIEW�q�S <6p�`U�`��NFI@;�FOC�U��;�PRI@�m�`�QY�TRIP>�qm�UN<`Md�� #@p�*eWA�RN)e6�SRTO�L%��g��ᴰO�NCORN��RAU䘠��T���w�VI�N�Le� $�גPATH9�גCwACH��LOG�!�LIMKR����v����HOST��!�b�R��OB�OT�d�IM>� �� ���Zq��Zq;�VCPU_A�VAIL�!�EX
	�!AN���q��10r��1r��1 �ѡ�.�p�  #`C����@$TOOL��$��_JMP� ����e$SS�����VSHIF��Nc�P�`ג��E�ȐR����OSU�R��Wk`RADILѮ��_�a��:�9a���`a�r��LULQ�$OUTPUT_3BM����IM�ABp �@�rTIL'SCO��C7� ������&��3 ��A���q���m�I�2G��pq�y@Md��}��yDJU��N_�WAIT֖�}Ҵ�{�%! NE�u��YBO�� ��� $`�t�S�B@TPE��NE�Cp�J^FY�nB_T��R�І�a$�H[YĭcB��dM� ��F� �p�$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"�`�"��[���P?� EaZABC~%��  $�"�R��
E`�$$C�LAS�������!pE`� � VI�RT]��/ 0ABS�����1 5�� < �!F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZi{0�-�AXL�p2��!�n63  �{tIN��qztPRE�����v��p�uLARMRECOV 9l�rwtNG�� .;	 A   �|.�0PPLIC���?5�p��Handlin�gTool o� �
V7.50P�/23-�  �P�B��
��_S�Wt� UP�!�� x�F0��t���A�ϐv� 86-4�� �it�y�� N�" �7DA5�� j�� QB@<��o�Noneisͅ�˰ ��T��]�!LAAx>�_l�V�uT��s9�UTO�"�Њt��y��HGAPON�
0g�1��Uh�D [1581�����̟ޟry����Q 1���p�,� 蘦���;�@��q_���"�" �c�.�H���D�HTTHKYX� �"�-�?�Q���ɯۯ 5����#�A�G�Y�k� }�������ſ׿1��� ��=�C�U�g�yϋ� �ϯ�����-���	�� 9�?�Q�c�u߇ߙ߫� ����)�����5�;� M�_�q������� %�����1�7�I�[� m����������!�� ��-3EWi{ ������ )/ASew�� ��/��/%/+/ =/O/a/s/�/�/�/�/ ?�/�/?!?'?9?K? ]?o?�?�?�?�?O�?��?�?O#O]���TO��E�W�DO_CL�EAN�����CNMw  � ��__/_A_S_�DS�PDRYR�O��H	Ic��M@�O�_�_�_ �_oo+o=oOoaoso��o�o���pB��v �u���aX�t������>9�PLUGG���G\��U�PRCvPB�@E��_�orOr�_��SEGF}�K [mwxq�O�O���p��?rqLAP�_ �~q�[�m�������� Ǐُ����!�3�x�TOTAL�f yx�_USENU�p��� �H���B��RG_�STRING 1�u�
�M�n�S5�
ȑ_I�TEM1Җ  n 5�� ��$�6�H�Z� l�~�������Ưد����� �2�D�I�/O SIGNA�L̕Tryout Modeӕ�Inp��Sim�ulatedב�Out��OV�ERR�P = 1�00֒In c�ycl��בProg Abor���ב��Statu�sՓ	Heart�beatїMH� Faul��Aler'�W�E�W�iπ{ύϟϱ������� �CΛ�A����8� J�\�n߀ߒߤ߶��� �������"�4�F�X�8j�|���WOR{pΛ ��(ߎ����� ��$� 6�H�Z�l�~���������������� 2PƠ�X ��A{ ������� /ASew��p���SDEV[ �o�#/5/G/Y/k/ }/�/�/�/�/�/�/�/�??1?C?U?g?y?PALTݠ1��z? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�Op�O�O_�?GRI�` ΛDQ�?_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o2_l�R��a\_�o" 4FXj|��� ������0�B�<T��oPREG�>��  f���Ə؏����  �2�D�V�h�z��������ԟ���Z��$�ARG_��D ?�	���;���  	�$Z�	[O�]�O��Z�p�.�SBN�_CONFIG S;��������CII_SAVE  Z�����.��TCELLSET�UP ;�%HOME_IOZ�~Z�%MOV_��
�REP�lU�(�UTOBACKܠ���FRwA:\z� \�,z�Ǡ'`�z���\ǡi�INI�0z����n�MESS�AG���ǡC���ODE_D������%��O�4�n�PAUS�X!�;� ((O>��ϞˈϾϬ� ���������*�`߀N߄�rߨ߶�g�l TSK  wͥ�_��q�UPDT+��d�!�A�WSM_C5F��;���'�>-�GRP 2:�?�+ N�BŰA��%��XSCRD1�1
N7� �ĥĢ�� ��������*����� ��r�����������7� ��[�&8J\n���*�t�GROU�N�UϩUP_N5A�:�	t���_ED�17�
� �%-BCKEDT-�2�'K&�`���-t��z�q�q�z����2t1������q�k�(/��ED3/��/�.a/�/;/M/ED4�/t/)?��/.?p?�/�/ED5`??�?<?.�?O�?�?ED6O�?qO��?.MO�O'O9OED7�O`O_�O.�O\_�O�OED8L_,�_�^-�_ oo_�_�ED9�_�_]o�_	`-9o�oo%oCR _ 9]�oF�o�k�� � NO_DEL���GE_UNU�SE��LAL_?OUT �����WD_ABOR�ﰨ~��pITR_�RTN��|NO�NSk���˥C�AM_PARAM� 1;�!�
 8�
SONY X�C-56 234�567890 �ਡ@���?}��( А\��
���{����^�H�R5q�̹��ŏR5y7ڏ�Aff���KOWA SC�310M
�x��>��d @<�
� ��e�^��П\�� ��*�<��`�r�g��CE_RIA_I��!�=�F���}�z� ��_LeIU�]������<��FB�GP 1.��Ǯ�M�x_�q�0�C*  ��V��C1��9��@��iG���CR�C]��Ud��l��s��R��T���[Դm��v���������� C����(�����=�{HE�`ONFIǰ��B�G_PRI 1�{V���ߖπ�Ϻ����������C�HKPAUS�� ;1K� ,!uD� V�@�z�dߞ߈ߚ��� �������.��R�<�hb���O���������_MOR��� �6��� 	 �����*��N�<��������?��q?$;�;����K��9��P���çaÃ-:���	�

 ��M���pU�ð��<���,~��DB����튒)
mc:c?pmidbg�f��:�  3���¥�p�/���������0� �s>ܑ۰��W�?�*�pY�pZUg�/V� ԋ��Uf��M/w�O/�
DEF 3l��s)�< buf.txts/��t/��ާ�)�	�`�����=L�Ͷ�*MC��1�����?43��1���t�īCz  BH�H�B�^B�$��B5�5@@��C���>'��Y
K�D\nD���C�|@8���.D�� @���=F�&��E�CeE�d��<�X�F��B��IY	���'w�K1���s���U.�p������BD�w�M@x8�K�C�2�����g@D�p@�0�EYK�EX��EQ�EJP �F�E�F� �G��>^F �E�� FB� �H,- Ge���H3Y��:�  �>�33 ����~  n8�~@F��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMO�FS�p�.8��)T}1��DE ��fF 
Q��;�(PG  B_<_��R�����	op6C4P�Y
s@ ]AQ�2s@�C�0B3�MaC{@@�*cw��UT�pFP?ROG %�z�o�oigI�q���v��ld�KEY_TBL � �&S�#� �	
��� !"�#$%&'()*+,-./01i��:;<=>?@A�BC� GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������vq���͓���������������������������������耇����������������������p`LCK�l4�p`��`STAT ��S_AUTO_DO����5�INDT_'ENB!���R�Q?��1�T2}�^�STO�Pb���TRLr`L�ETE��Ċ_S�CREEN ~�Zkcsc���U��MMENU �1 �Y  <�l�oR�Y1�[��� v�m���̟�����ٟ �8��!�G���W�i� �������ïկ��4� ��j�A�S���w��� ��迿�ѿ����T� +�=�cϜ�sυ��ϩ� ��������P�'�9� ��]�o߼ߓߥ���� ����:��#�p�G�Y� ����������$� ���3�l�C�U���y� ���������� ��	�VY)�_MANU�AL��t�DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�mg�(&/~&lMZ�IdPx�@P@#ONTIM6ه� d�`&��
�e�MOTNE�ND�o�RECO_RD 1(�[g2�/{�O��!�/k y"?4?F?X?�(`?�? �/�??�?�?�?�?�? )O�?MO�?qO�O�O�O BO�O:O�O^O_%_7_ I_�Om_�O�_ _�_�_ �_�_Z_o~_3o�_Wo io{o�o�_�o o�oDo �o/�oS�oL �o����@�� �+�yV,�c�u�� ������Ϗ>�P��� ��;�&���q���򏧟 ��P�ȟ�^������ I�[����� ���$��6��������"TO�LERENCwB����L�Ϳ C�S_CFG )��/'dMC:�\U�L%04d.'CSV�� c��/#[A ��CH��z� �//.ɿ��(S�R�C_OUT *���1/V�SGN� +��"��#��09-FEB-�20 18:44~027-JANp��21:48+ P;��ɞ�/.���f�pa�m�?�PJPѲ���VERSION �Y�V2.�0.�ƲEFLO�GIC 1,� 	:ޠ=�ޠ�L��PROG_E�NB��"p�ULS�k' ����_WRSTJNK ��"f�EMO_OPT_�SL ?	�#
� 	R575 /#=�����0�B��>��TO  �ݵ�l���V_F EX��d�%��PATHw AY�A\�����5+ICT�F�u-�j�#�egS�,�ST?BF_TTS�(�	�d���l#!w�� M�AU��z�^"MSWX�.�<�4,#�Y�/�
!J�6%�ZI~m��$SB�L_FAUL(�0��9'TDIA[�1�<�<� ����12345678#90
��P��H Zl~����� ��/ /2/D/V/h/��� P� ѩ �yƽ/��6�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�,/�gUMP���� ��ATR���1OC@P�MEl�OOY_TE{MP?�È�3F�8��G�|DUNI��.��YN_BRK �2_�/�EMGDI�_STA��]��EN�C2_SCR 3�K7(_:_L_^_ l&_�_�_�_�_)��C�A14_�/oo/o�AoԢ�B�T5�K�ϋo~ol�{_�o�o �o'9K]o �������� �#�5��/V�h�z��� �`~�����ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T���x������� ��ү�����,�>� P�b�t���������ο ����(�f�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ���������:�  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� �����*<N `r������ �&8J\n ���������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?��? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O��O�O__NoETM�ODE 16�5]�Q �d�X�
X_j_|Q�PRRO�R_PROG �%GZ%�@��_  ��UTABLE  G[�?oo)oRj�RRSEV_NU�M  �`WP��QQY`�Q_AU�TO_ENB  q�eOS�T_NOna� 7G[�QXb�  *��`��`��`��`d`+�`�o�o�o�dHISUc�QOP��k_ALM 18.G[ �A��l�P+�ok}������o_Nb�`  �G[�a�R
�:PTC�P_VER !�GZ!�_�$EXTLOG_REQvs�i\�SIZe�~W�TOL  �Q{Dzr�A W�_BWD�p��xf́�t�_DI�� 9�5�d�T�QsRֆSTEP��:P�_OP_DOv�f��PFACTORY�_TUNwdM�E�ATURE :��5̀rQH�andlingT�ool �� \s�fmEngl�ish Dict�ionary��r�oduAA �Vis�� Mas�ter����
E�N̐nalog �I/O����g.f�d̐uto So�ftware U�pdate  F� OR�mati�c Backup~��H596,��ground E�ditޒ  1 �H5Came�ra�F��OPL�GX�ell𜩐IwI) X�ommՐsshw���com��sco���\tp����pane��  �opl��tyle select��/al C��nJ�Ց�onitor��R�DE��tr��R�eliab𠧒6�U�Diagnosx(�푥�5528��u��heck S�afety UI�F��Enhanc�ed Rob S�erv%�q ) �"S�r�User �Fr[�����a��xt. DIO ��fiG� sŢ��e�ndx�Err�L&F� pȐĳr됮�� ����  !��F�CTN Menu�`�v-�ݡ���TPw Inېfac��  ER J�GC�pבk Ex�ct�g��H558���igh-Spe�x�Ski1�  2�
P��?���mm�unic'�ons��&�l�ur�ې���ST Ǡ��co�nn��2��TXP�L��ncr�st�ru����"FAT�KAREL �Cmd. LE�u�aG�545\��R�un-Ti��En=v��d
!����ؠ++�s)�S/W���[�LicegnseZ��� 4T��0�ogBook(�Syڐm)��H5�4O�MACROs�,\�/Offsen��Loa�MH��ܽ���r, k�Me�chStop P�rot���� li�c/�MiвShiqf����ɒMixx���)���xSPS�M�ode Swit�ch�� R5W�M�o�:�.�� 74� ���g��K�2~h�ulti-T=��M���LN (�Pos�Regi�ڑ������d�ݐt 'Fun�ǩ�.�����Num~����� �lne��ᝰ A�djup����� � - W��tat�uw᧒T�R�DMz�ot��scWove U�9����3Ѓ�uest' 492�*�o������62;�SNPX� b ���8 J7<`���Libr��J�#48���ӗ� �Ԅ��
�6O�� Par�ts in VCCMt�32���	��{Ѥ�J990��/�I� 2 P��T_MILIB��H�:��P�AccD�L�o
TE$TX��n��ap1S�Te����pkey��w����d��Une�xceptx�mo�tnZ��������є�� O����� 90J�єSP CSXC<�f���6�� Py�We}���gPRI�>vrЮt�men�� ��iPɰa������vGrid�pl�ay��v��0�)�H�1�M-10iA�(B201 �2�\� 0\k/�Ascii�l�Т�ɐ�/�Col��ԑGu�ar� 
�� /Pl-�ޠ"K��st{�Pat ��!S�C�yc�҂�ori�e��IF8�ata- quҐ�� ƶ���mH574��RL���am���Pb�H_MI De3�(b�����PCϺ�Pa�sswo+!��"P�E? Sp$�[���t�p��� ven��T�w�N�p�YELL�OW BOE	k$A;rc��vis��y3*�n0WeldW��cial�7�V#t&�Op����1y�� 2F�a�por1tN�(�p�T1�T�0 �� ��xy]�&kTX��tw�igjx�1� b� ct\��JPN ARCPSU PR��oݲ�OL� Sup�2f�il� &PAɰאc{ro�� "PM(�X���O$SS� eв7tex�� r���z=�t�ssagT��P��P@�Ȱ�����rtW��H'>�r�dpn��n1�
t�!� z ��a�scbin4ps�yn��+Aj�M �HEL�NCL �VIS PKGS� PLOA`�MB� �,�4VW�R�IPE GET_�VAR FIE �3\t��FL[�O�OL: ADD �R729.FD �\j8'�CsQ�QE���DVvQ�sQNO? WTWTE��}PD  �^��biR�FOR ��ECT�n�`��ALSE �ALAfPCPMO�-130  M"� #h�D: HANG FROMmP��AQfr��R70�9 DRAM A�VAILCHEC�KSO!��sQVPC�S SU�@LIM�CHK Q +P~dF_F POS��F�Q� R5938�-12 CHAR�Y�0�PROGRAy W�SAVEN`wAME�P.SV��7��$En*��p?F�U�{�TRC|� S�HADV0UPDA�T KCJўRST�ATI�`�P MU�CH y�1��IM�Q MOTN-0�03��}�ROBO�GUIDE DA�UGH�a���*�t�ou����I� Šh�d�ATH�PepMO�VET�ǔVMX�PACK MAY ASSERT�Dn��YCLfqTA�r�BE COR v�r*Q3rAN�pRC� OPTIONS�J1vr̐PSH-�171Z@x�tcǠSU1�1Hp^9R!�Q��`_T�P��'�j��d{tby ap?p wa 5I�~d��PHI���p�aTE�L�MXSPD �TB5bLu 1��UBl6@�qENJ`CE2��61��p��s	�m�ay n�0� R�6{�R� �Rtrasff)�� 40*��p��fr��sys�var scr �J7��cj`DJUD��bH V��Q/�PSET ERR`�J` 68��PND�ANT SCRE�EN UNREAh��'�J`D�pPA��z�pR`IO 1����PFI�pB�pGROUN�PD��G��R��P�QnRSVIP �!p�a�PDIGIT� VERS�r}BL�o�UEWϕ P0�6  �!��MAG`p�abZV�DI<�`� SSUE�ܰ��EPLAN J=OT` DEL�pݡ�#Z�@D͐CAL9LOb�Q ph��RޫQIPND��IM�G�R719��MwNT/�PES �puVL�c��Hol�08Cq���tPG:�`C��M�canΠ��p�g.v�S: 3D� mK�view ed�` �p��ea7�:��b� of �Py����ANNOT ACCESS M��tƁ*�t4s a���lok��Flexj/:�Rw!mo?�PA?�-�����`n�pa SNBPJ? AUTO-�06f�����TB��PIAB{LE1q 636���PLN: RG$�pul;pNWFMDB��VI���tWIT �9x�0@o��Qui�#0�ҺPN RRS�?pUSB�� t & remov�@� )�_��&AxEPF�T_=� 7<`�pP�:�OS-144 ��h s�g��@�OST� � CR�ASH DU 9^��$P�pW� �.$��LOGIN���8&�J��6b04�6 issue �6 Jg��: Solow �st��?c (Hos`�c����`IL`IMPR�WtSPOT:Wh�:0�T�STYW ./�VMGR�h�T0wCAT��hos���E�q��� �O:�S:+pRTU' k�e-S� ����E:���pv@�2�� t\h�ߐ��m ��alļ�0�  $�H� W�A͐��3 CNT�0 T�� Wro>U�alarm���0s�d � �0SE1���t�r R{�OMEBp����K� 55��R�EàSEst��g �    �KA7NJI�no����INISITALcIZ-p�dn1weρl<��dr�� lx`~�SCII L�fails w��y ��`�YSTEa�p��o��Pv� IIH����1W�Gro>Pmo ol\wpSh@��P��Ϡn cfl�xL@АWRI �OGF Lq��p?�F��up��de-re�la�d "AP�o SY�ch�Abe�twe:0IND 1t0$gbDO����r� `�GigE��#operabi-lf  PAbHi�H`���c�lead�\�etf�Ps�r�O�S 030�&: fi=g��GLA )P ���i��7Np tpkswx�B��If�Ag������5aE�a EXCE#dU�_��tPCLOS��"r[ob�NTdpFa�U�c�!���PNI�O V750�Q1p��Qa��DB ��b�P M�+P�QED��DET��-� \r�k��ONLINEhSBUGIQ ߔĠ,i`Z�IB�S ap�ABC JARK�YFq� ���0MI�L�`� R�pNД \�p0GAR��D*pqR��P�"! jK�0cT�P�Hl#n�a��ZE V�� TA;SK�$VP2(�4`�
�!�$�P�`WIB�PK05�!FȐB�/��BUSY R7UNN�� "��d���R-p�LO��N�DIVY�CUL���fsfoaBW�p���30	V���ˠIT`�a50�5.�@OF�UN#EX�P1b�af�@�}E��SVEMG� �NMLq� D0pC?C_SAFEX 0c��08"qD �PETr�`N@�#J87��B��RsP�A'�M��K�`K�H GU�NCHG۔MEC�H�pMc� T�  �y, g@�$ OR?Y LEAKA�;�ޢSPEm�Ja��V�tGRIܱ�@އCTLN�TRpk�FpepR�j50�EN-`IN�����p� �`�Ǒk!��T3�/dqo�STO�0A�#�L�p �0�@�Q��АY�&�;pb1T!O8pP�s���FB�@�Yp`�`DU��aO��supk�t4 � P�F�� Bnf�Q�PSV�GN-1��V�SRSR)J�UP�a2�Q�#D�q l O���QBRKCTR 5Ұ�|"-�r�<pc��j!INVP�D ZO� ��T`h#�Q�cH�set,|D��"D�UAL� w�2*BRVO117 A]��TNѫt�+bTa24�73��q.?��sAU�z�i�B�compl�ete��604.�� -�`han�c�U� F��eN8��  ��npJtPpd!q��`��� 5h'596p�!5d�� @"p�P�P�Q�0�P2�p �A� xP��R(}\xP�e� aʰI���E���1��p� j  �� xS?P�^P �A��AxP�q 5 sig:��a��"AC;a���
�bCexPb_p���.pc]l<bHbc?b_circ~h<n�`tl1�~`xP`o�d�xP�b]o2�� �cb��c�ixP�jupfr�m�dxP�o�`exe��a�oFdxPtped�}o��u`�cptli1bxzxP�lcr�xrxP\�blsazEdxP_fm�}gcxP�x�� �o|sp�o�mc(��o'b_jzop�u6��wf��t��wms�1�q��sld�)��jm!c�o\�n��nuhЕ�ƭ|st�e��>�pl�qp�iwck���u�vf0uߒ��lvi�sn�Cgacul�wQ
E F  !� Fc.fd�Qv��� qw���Data� Acquisi��nF�|1�RR63�1`��TR�QDMCkM �2�P75H�]1�P583xP1��[71��59`�5�P57<PxP�Q����a(���Q��o pxP^!daq\�oA���@�� ge/�et�dms�"DMER9"؟,�pgdD����.�m���-��qaq1.<᡾xPmo��h����f{�u�`13��M�ACROs, Sksaff�@z����0E3�SR�Q(��Q6��E1�Q9ӡ�R�ZSh���PxPJ643�@7bؠ6�P�@�PRS�@����e �Q�UС P�IK�Q52 PT�LC�W��xP3 (��p/O��!�Pn� �xP5��03\�sfmnmc "MNMCq�<��Q��5\$AcX�FM��� ci,Ҥ�X����cdpql+�
�sk�SK�<xP�SH560,P���,�y�refp �"REFp�d�A�jlxP	�of�OFc�l<gy�to�TO_�x���ٺ���+j�e�u��caxis�2�xPE�\�e�q"I�SDTc��]�pr7ax ��MN��<u�b�isde܃h��\�w�xP! isb�asic��B� yP]��QAxes��R6������.�(B9a�Q�ess�� xP���2�D�@�z�atis���(�{������~��m��FM�c�u�{�
ѩ�MNIS��ݝ����x�����ٺ��x� j75���Devic�� �Interfacx�RȔQJ754��� xP�Ne`�� xP�ϐ2�б����{dn� "DNE�����
tpdnui�5UI��ݝ	bd��bP�q_rso�fOb
dv_aro��u�����stchkc��zp	 �(}onl��G!ffL+H�J( ��"l"/�n�b��<�z�hamp��T�eC�!i�a"�59�0�S�q��0 (�+P�`o�u�!2��xpc_2�pcchm��CH�MP_�|8бpev�ws��2쳌pcs|F��#C SenxPacro�U·�-�R6�Pd�xPk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GEM�,\i(��Dgesnd�5���H{�}Ha�@csy���c�Isu�xD��Fmd��I��7�4����u���AccuCal�P�4� ��ɢ�7ޠB0��6+6f�6��99\aFF q��S(�U��2�
X�p0�!Bd��cb_�Sa{UL��  �� �?�ܖto��otp�lus\tsrnPغ�qb�Wp��t����1��Tool (?N. A.)�[K�7�Z�(P�m���țbfcls� k9�4�"K4p��qtp{ap� "PS9|H�stpswo��0�p�L7��t\�q�� ��D�yt5�4�q��w��q��� �M�uk��rkey����s��}|t�sfeatu6�CEA��� cf)t\Xq`�����d�h5����LRC0�md�!�5!87���aR�(�����2V��8c?u3l\�pa3}H�&r-�Xuļ��t,�� �q " �q�Ot��~,���{�/ ��1c�}����y�p� r��5���S�XAg�-�xy���Wj874�- iRVis���Queu�� �@��-�6�1���(����u���tӑ�����
�tpvtsn "VTSN�3C�+�:� v\pRDV����^*�prdq\�Q�&�vstk=P�������nm&_�դ�c�lrqν���ge�t�TX��Bd���apoQϿ�0qstr�D[� ��t�p'Z�����npv��@�enl IP0��D!x�'�|���csc ߸��tvo/@��2�q���vb� ���q���!���h]����(� Cont�rol�PRAX:�P5��556�A@�59�P56.@56r@5A�J69$@�982 J552 IDVR7�hqA���16�H���La��� ��Xe�frlparm.f�7FRL�am��C9�@(F�����w6�{���A��QJ64�3�� 50�0LS�E
_pVAR $SGSYSC���RS_UNITS� �P�2�4tA�TX�.$VNUM_OLD 5�1�xP{�ƈ50+�"�` Funct���5tA� P}��`#@�`3�a0�c�ڂ��9���@H5 נ� �P���(�A�� ��۶}����ֻ�}��bPRb�߶~pp=r4�TPSPI�3�}�r�10�#;A� �t�
`���1���96�����%C�� Aفz��J�bIncr�	 ����\���1o5�qni4�MNIN�p	xP�`���!��H�our  �� 2�21 ~�AAVM��̳�0 ��TU�P ��J54s5 ��6162��VCAM  �(�CLIO= ��R6�N2��MSC "P� �STYL��C�28~ 13\��NRE "FH�RM SCH^��DCSU%OR�SR {b�04 ~�EIOC�1{ j 542 � �os| � egiCst�����7��1�MASK6�934"7 ��OOCO ��"3��8��2���� 0� HB��� 4�"39N� Re�� ��LCHK
%OPL�G%��3"%MHCMR.%MC  ; 4? ���6 dPI�5�4�s� DSW%M�D� pQ�K!637��0�0p"�1�Р"4� �6<27 CT�N K � 5 ����"7��<25�%/�T��%FRDM� �Sxg!��930 FB�( NBA�P� ( HLB  Men��SM$@jB( PVC� ��20v��2H�TC�CTM�IL��\@PAC c16U�hAJ`SAI N\@ELN��<29s�UECK �b��@FRM �b�O�R���IPL��R>k0CSXC ����VVFnaTg@HT�TP �!26 ���G�@obI�GUI"%IPGS|�r� H863 qbp�!�07r�!34 �r>�84 \so`!� Qx`CC3 Fb�21��!96 rb!531 ���!53R% E1!s3!��~�.p"�9js VATFUJG775"��pLR6^R�P�WSMjUCT�O�@xT58 F!890���1XY ta3!�770 ��88M5�UOL  GTSox
�{` LCM �r�| TSS�EfP6 |W�\@CPE `���0VR� l�QNL�"��@001 imrb�c3 =�b�0���0�`6 w�b-P�- R-�b8n@5EW�b9 �Ґa� ���b�`ׁ�b2 2'000��`3��`	4*5�`5!�c�#$��`7.%�`8 h6�05? U0�@B6iE"aRp7� !Pr�8 t�a@�tr2O iB/�1vp3�&vp5 Ȃtr9Σ�a�4@-p�r3 F��r5&�re`u��r�7 ��r8�U�p9? \h738�a�_R2D7"�1f���2&�7� �3 S7iC��4>w5Ip��Or60 C�L�1lbEN�4 I�pyL�`uP��@N�-PJ8�2N�8NeN�9 H�r`�E�b7]�|���q8�Вࠂ9 2���a`0�qЂ5�%U�097 0��@18�0���1 (�q�3 5R���0����mpU��0�0�7�*�H@(q�\P"R;B6�q124�b;�0�@���@06� x�3 pB/x�u ��~x�6 H606�a�1� ��7 6 ����p�b155� ����7jUU1632 �3 g���4*�65 2e 1"_��P�4U1`��ҢB1���`0'�17�4 �q��P�E18�6 R ��P�7 t��P�8&�3 (��90 B/�s1981����@202���6 3���A�RU�2� d��2 b2$h`��4�᪂2�4�&��19v Q�2��u�2d�Tpt2� ��H"�a2hP�$�5���!#U2�p�p
�2�p��B�@5�0-@��8 @�9��TX@�� �e�5�`rb26Af�2 ^R�a�2Kp��1y�bQ5Hp�`
�5�0@�0gqGA���a52ѐ��Z��6�60ہ5� Jׁ2��8�E��9�ESU5@ٰ\�q5hQT`S�2ޖ5�p\w�@۲�pJ �-P��5�p�1\t�H�4��PC2H�7j��phiw�@���P�x��559 ldu� P�D���Q�@������� �`.��Pt>��8�581�"6�q58�!AM۲T��A iC�a589`��@�x����5 �a��12׀0.�1����,�2����,�!P\hI8��Lp ��,�7���6�0840\��A?NRS 0C}A��0p��{��ran��FRA��Д�е� ��A%���ѹ�Ҍ� ����(����Ќ��� �З���������ь����$�G��1��ը����������� xS�`q�  X�����`64��M���iC/50T-H�������*��)p46���� C��N����mw75s֐� Sp��b46��v�����^�M-71?�7�������42������dC��-�а�70�r$�E��/h�����O$��rD���c7c7C�q��Ѕ���L��/��2\imm7c7�g������`���(�� e�����"������`�a r��c�T,����"��,�� ��x�<Ex�m77t����k���5�����)�;iC��-HS- � B
_�>���+����7U�]���Mh7�s��7�������-9?�/260L_������Qҡ������]�9pAA/@���q�S�������h6251��c��92���p����.�)92c0� g$�@�����)$��85$���pylH"O"�
�21���t?�350����p��`$�
�� �350!����0��9�U/0�\m9��M9A3���4%� s��3�M$��X%u���"him98J3����� i Ad�"m4~�103p�x� ����h794̂�&R���H�0����\� ���g�5AU��՜��0 ���*2��00��#06�АՃ�է!07{r ������� ��kЙ@����EP�#������?��8#!�;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?���CD25L�����0�"l�2BL 
#��B��\20�2_� r�re���X��1�� N����A@��z��`�C�pU��`��0�4��DyA�\�`f Q��sU���\�5�  ��� �p�^P��<$85����+P=�ab1l���1LT��lA8��!uDnE(�20T⧰J�1 e�bH85����b�Ռ�5[�16�Bs��������d2p��x��m6t! `Q����bˀ���b#�(�6iB;S�p�!� �3� ��b�s��-`�_�W8�_�����6I	$�X5�1�U815��R�p6S��� �/�/+q�!�q��`��6o��5m[o)�m6�sW��Q�?��se�t06p ��3%H�5��10p$����g/��JrH��  s��A�856�Ȝ��F�� ���p/2���h�܅�✐)�5���̑v��(��m	6��Y�H�ѝ̑m�Q6�Ҝ��a6�DM��F��-S�+��H2� ����Ҽ�� �r̑���✐��l���p�1���F���2�\t;6h T6H��� �Ҝ�'Vl���ᜐ��V7ᜐ/����;3A7��p~S��������4�`圐�V���*!3��2�PM[���%ܖO�chn��v�el5����Vq���_arp#��̑�.���?2l_hemq$�.�'�6415���5� ��?����F�����A5g�L�ј[���1��Ȝ�𙋹1����M7NU�М��eʾ�����uq$D;��-�4��3&H�f�c�Ĝ�h� ������u��� 㜐��ZS�!ܑ4���M-����S�$̑��� �� 0��<�����\07shJ�H�v �À�sF��S*󜐳� ��̑���vl�3�A�T�#��QȚ�Te��q�cpr����T@75j�5�dd�̑1�(UL�&� (�,���0�\�?���̑��a�� xSPA���a�e�w�2��d(�	�2�C��A/����\�+p�����21s (ܱ�CL S�� ��B̺��7F���4?�<�lơ1L����c� ���u9�0����Ce/q��O���9�K��r9 (��,�Rs��ז�5�G�m2�0c��i��w�2 ��:�0`�$��2�2lҀ0�k�X�S� ,�ι2���O���1!41�w���2T@� _std��G�y� �ң�H� jdgm����w0 \� �1L���	�P�@~�W*�b��t 5��(����3�,���AE{������L��&�5\L��3�L�@|#~���~!���4�#@��O����h�L6A�������2璥����44�����[6\j4s��·���# ��ol�E"w�8Pk� ����?0xj�H1�1Rr��>��]�2a�2�Aw�P ��2��|41 �8��ˡ��{� �%�A<��� +�?�l��0�&0�"��|�`Am1�2� �ػ��3�HqB�� ��K�R��ˑb�W��� Fs���)�ѐ�!����a�1����5��16�16C��C����0\imBQ��d�P���b��\B5�-���DiL���O�_�<ѠPEtL�E�RH�Z�p�Pgω�am1l�� u���̑�b�<����<�$�T�̑�F���@�Ȋ�Dpb��X"��hr��p� ����^P��9�0\� j�971\kckrcfJ�F�s�����c���e "CTME��r���ɛ��a�`ma�in.[��g�`r#un}�_vc�#0 �w�1Oܕ_u����bctme��Ӧ�`ܑޅj735�- �KAREL UsKe {�U���J�P�1���p� Ȗ �9�B@��L�9��7�j[�atk208� "K��Kя��\��9��a��̹���N�cKRC�a�o ��kc�qJ�&s����� Grſ�fsD��:y��s��ˑ1X\j|хrd�tB�, ��`.v�q�� �sǑIf�Wf�j52�TKQut_o Set��J�w H5K536(��932���91�58�(�9�BA�1(�74�O,A$�(TCP �Ak���/�)Y� ��\tpqtoo�l.v��v���!? conre;a#��Control �Re�ble��CNRE(�T�<�4�2����D�)���S�5524��q(g�� (򭂯�4X�cOux�\sfwuts�UTS`�i�栜���t�棂Č�? 6�T�!�SA OO+D6����@�����,!��6cp+� igt�t6i��!I0�TW8 ���la��vo58�o�bF� �򬡯i�Xh��!X�k�0Y!8\m6e��!6EC���v��6����������<16�A���A�6s�����U�g�T|ώ���r1"�qR��˔Z4�T��@���,#�eZp)g� ���<ONO0���uJ���tCR;��F�a� x�SP�f��prds�uchk �1��2H&&?���t��*D%$ �r(�✑�娟:r���'�s�qO��<sc�rc�C�\At�trldJ"o�\�V�����Paylo�n�firm�l�!�87��7��A�3ad�! �?ވI�?p4lQ��3��3"�q��x pl�`���d7��l�calC�uDup���;��mov��<���initX�:s�8O��a�r4 ��r�67A4|�e Ge?neratiڲ����7g2q$��g R� (Sh��c �,|�bE��$Ԓ\��:�"��4��4X�4�. sg��5�ЌF$d6"e;Qp "SHAP�TQ ongcr pGC��a(�&"� ��"GD�A¶��r6�"axW�/�$dataX<:s�"tpad��[q�%tput;a__O7@;a�o8�1�yl+s�Ar�?�:�#�?�5x�?�:c O�:y O�:�$IO�s`O%g�qǒ��?�@0\��"o�j9�2;!�Ppl.Co�llis�QSkip#��@5��@J��D���@\ވ�C@X�7ҥ�7�|s2��pt7cls�LS�DU��k?�\_ ets�`�< \�Q��@����`dcKqQ�FC�;��J,�n��` (���4eN����T �{���'j(�c������/IӸaȁ��̠H������зa�e�\mcclmt �"CLM�/��� moate\��lmp�ALM�?>p7qm!c?����2vm�q��8%�3s��_sv90�_x_msu�2L^va_� K�o�{in�8�(3r<�c_logpr��rtrcW񊬯 �v_3�~yc0��d�<�te���der$cCe� Fiρ�R��Q��?�l�enter ߄|��(Sd��1ثTX�+fK�r�a9�9sQ9+�5�r\�tq\� "FND�R���ST�Dn$LANG.�Pgui��D⠓0�S������sp�!ğ֙uf�ҝ�s����$�����e+�=���� �����������w�H�r\fn_�ϣ��$`�x�tcpma��-� TCP�����R638 R�Ҡ�V�38��M7p,�� �Ӡ�$Ӡ�8p0Р�VSl,�>�tk��99�a ��B3���PզԠ��D�2�����UI��t��� hqB���8��������p����re�ȿ��exe@4φ�B���e388�ԡG�rmpWX���var@�φ�3 N�����vx�!ҡ��~q�RBT $c�OPTN a�sk E0��1�R� MAS0�H59}3/�96 H50�Vi�480�5�H0Ԉ�m�Q�K��7�0�g�Pl�h0ԧ�2�OR�DP��@"��t/\mas��0�a�� "�ԧ�����k�գR����ӹ`m��b��&7�.f��u�d��}r��splayD��E���1w�UPDT� Ub��887 (&��Di{���v�Ӛ� �Ԛ⧔��#�B��㟳>��o  ����a�䣣��60q��B��|���qscan���B���ad@�������q`�䗣�#�p�К�`2�� vlv ��Ù�$�>�b����! S��Easy</К�Util���>��511 J���r��R7 ��Nor֠>��inc),<6Q
�� �`c��"4�[����986FVRx bSo����q�nd6� ���P��4�a\ (��
   �������d��K�rbdZ���men7����- Me`tyFњ�Fb�0�TUaN�577?i3R��\�5�u?��!� n���f������l\mh�Ц�ű8E|hmn�	��B<\O���e�1"�� l!��y���
��\|p����B���Ћmh�@��:. aG!���/�t�5�5�6�!X�l�.us���Y/k)ensubL���eK�h�� �B \1;5g?y?�?�?D���?*rm�p�?Ktbox O2K|?�G��C?A%ds���?1��#� �TR��/��P �4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ăd�Q3t.�P׀al��P+OP517F��IN0a��Q(}g���PESTf3ua@�PB�l�ig�h�6�a�q��P � x9S��`  n�0m�bumpP�Q969g�69�Qq��P0��baAp�@Q� B�OX��,>vche8�s�>vetu㒣^=wffse�3�Ā�]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q8<twaǂ tp�Q҄�Taror Re'cov�b�O�P�642����a�q���a⁠QErǃ�Qr!y�з`�P'�T�`�a�ar������	{'�paok971��71��`m���>�pjot���PXc��C�1�adb �-�ail��nagx���b�QR629�a�Q��b�P  ��
  �P���$$CL[q �����������$�PS_DIGsIT���"�!�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*���1:PRODU�CT�Q0\PGS�TK�bV,n��99�\����$FEAT_IN�DEX��~��� 搠IL�ECOMP ;���)��"��S�ETUP2 <����  �N !�_AP2�BCK 1=�  �)}6/E+%,/i/��W/�/ ~+/�/O/�/s/�/? �/>?�/b?t??�?'? �?�?]?�?�?O(O�? LO�?pO�?}O�O5O�O YO�O _�O$_�OH_Z_ �O~__�_�_C_�_g_ �_�_	o2o�_Vo�_zo �oo�o?o�o�ouo
 �o.@�od�o� ��M�q��� <��`�r����%��� ̏[�������!�J� ُn�������3�ȟW� �����"���F�X�� |����/���֯e��� ���0���T��x��� ���=�ҿ�s�ϗ�@,ϻ�9�b�� P/� 2) *.V1Riϳ�!�*����`������PC�|7�!�FR6:"�"c��χ��T��� ��Lը��ܮx��ﶏ*.F��>� �	�N�,�k��ߏ��STM �����Qа����!�iPen�dant Panel���H��F����4������GIF �������u����JPG&P��<�����	PANE�L1.DT��@������2��Y�G��
3 w�����//�
4�a/�O///�/��
TPEINSO.XML�/����\�/�/�!Cust�om Toolb�ar?�PAS�SWORD/��FRS:\R?? �%Passwo�rd Config�?��?k?�?OH� 6O�?ZOlO�?�OO�O �OUO�OyO_�O�OD_ �Oh_�Oa_�_-_�_Q_ �_�_�_o�_@oRo�_ voo�o)o;o�o_o�o �o�o*�oN�or� �7��m�� &���\�����y� ��E�ڏi������4� ÏX�j��������A� S��w�����B�џ f�������+���O�� �������>�ͯ߯t� ���'���ο]�򿁿 �(Ϸ�L�ۿpς�� ��5���Y�k� ߏ�$� ���Z���~�ߢߴ� C���g�����2��� V����ߌ���?�� ��u�
���.�@���d� �����)���M���q� ����<��5r �%��[� &�J�n�� 3�W���"/� F/X/�|//�/�/A/ �/e/�/�/�/0?�/T? �/M?�??�?=?�?�? s?O�?,O>O�?bO�? �OO'O�OKO�OoO�O _�O:_�O^_p_�O�_ #_�_�_Y_�_}_o�_��_Ho)f�$FIL�E_DGBCK �1=��5`��� ( ��)
SUMMA�RY.DGRo�\�MD:�o�o
`�Diag Sum�mary�o�Z
C?ONSLOG�o�o�a
J�aCon�sole log�K�[�`MEMCHECK@'�o��^qMemory� Data��W��)�qHAD�OW���P��s�Shadow C?hangesS�-c�-��)	FTAP=��9����w`q�mment TB�D׏�W0<�)�ETHERNET�̏�^�q�Z��aE�thernet �bpfigurat�ion[��P��DCSVRFˏ��Ïܟ��q%�� ve�rify all�ߟ-c1PY���DIFFԟ��̟a��p�%��diffc���q��1X�?�Q��� ����X=��CHGD��¯ԯi��px��� ����2`�G�Y�� ��� �GD��ʿܿ�q��p���Ϥ�FY�3h�O�a��� ��(�GD�������y��p�ϡ�0�UPDATES.������[FRS:\������aUpda�tes List����kPSRBWLOD.CM.��\���B��_pPS_ROBOWEL���_�� ��o��,o!�3���W� ��{�
�t���@���d� ����/��Se�� ���N�r � =�a�r� &�J���/� 9/K/�o/��/"/�/ �/X/�/|/�/#?�/G? �/k?}??�?0?�?�? f?�?�?O�?OUO�? yOO�O�O>O�ObO�O 	_�O-_�OQ_c_�O�_ _�_:_�_�_p_o�_ o;o�__o�_�o�o$o �oHo�o�o~o�o7 �o0m�o� �� V�z�!��E�� i�{�
���.�ÏR��� �������.�S��w� �����<�џ`���� ��+���O�ޟH�������8���߯n�����$FILE_��P�R���������� �M�DONLY 1=�4�� 
 � ��w�į��诨�ѿ�� �����+Ϻ�O�޿s� ��ϩ�8�����n�� ��'߶�4�]��ρ�� �߷�F���j����� 5���Y�k��ߏ��� B�����x����1�C� ��g������,���P� ��������?��L�u�VISBCK�R�<�a�*.VD�|�4 FR:\���4 Vis�ion VD file� :Lb pZ�#��Y� }/$/�H/�l/� /�/1/�/�/�/�/�/  ?�/1?V?�/z?	?�? �???�?c?�?�?�?.O �?ROdOO�OO�O;O �O�OqO_�O*_<_�O�`_�O�__%_�_�M�R_GRP 1>�4�L�UC4 w B�P	 ]��ol`�*u����RHB ���2 ��� ��� ���He �Y�Q`orkbIh�oJd�o�Sc�o�oO\�d�Nc�Ly���F�5U�aTǪ؋�o�o �A�B�-\�A�.�Q6��ߞ;o%F}?R?��?��Zlq�Q�?�5�xq}E�?� F@ �r�d��a}J��NJk��H9�Hu���F!��IP��sX~�`�.9��<9�8�96C'6<?,6\b�1��,.�g�R���6x�PA�����|�ݏx��� %��I�4�F��j��� ��ǟ���֟��!���E�`r�UBH�P� �~�������W
�6�P;�uPI��a˯�o�e�Q cB��P5���@�33�@���4�m�,�@U�UU��U�~w�>u?.�?!x�^���ֿ���3��=[�z�=�̽=�V6<�=�=��=$q��~���@8�i7G���8�D�8?@9!�7ϥ��@Ϣ���cD�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p���������>p�� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__>���  DE_�Hly_�\@@m_B�=��vR/��I�O�SMT
�G�SUoo&o�RHOSTC�19H�I� ��zM�SM�l[�bo�	127.�0�`1�o  e �o�o�o#z�oF�Xj|�l60s	a�nonymous������� (ao�&�&��o� x��o������ҏ�3 ��,�>�a�O���� ������Ο�U%�7�I� �]����f�x����� ���ү����+�i� {�P�b�t�������� ����S�(�:�L� ^ϭ�oϔϦϸ���� ��=��$�6�H�Zߩ� ��Ϳs���������� � �2���V�h�z�� �߰���������
�� k�}ߏߡߣ���߬� ��������C�*< Nq�_����� �-�?�Q�c�eJ�� n������ �/"/E�X/j/|/ �/�/�%'/? [0?B?T?f?x?��? �?�?�?�??E/W/,O�>OPObO�KDaENT� 1I�K P!\�?�O  �P�O �O�O�O�O#_�OG_
_ S_._|_�_d_�_�_�_ �_o�_1o�_ogo*o �oNo�oro�o�o�o	 �o-�oQu8n �������� #��L�q�4���X��� |�ݏ���ď֏7����[���B�QUICC0��h�z�۟��A1ܟ��ʟ+���2,����{�!ROU�TER|�X�j�˯!?PCJOG̯���!192.168.0.10���}GNAME !��J!ROBOT��vNS_CFG �1H�I ��Auto-s�tarted�$FTP�/���/�? ޿#?��&�8�JϏ? nπϒϤ�ǿ��[���`���"�4�G�#��� ��������������� �����&�8�J�\�n� ������������� �/�/�/F���j��ߎ� ������������ 0S�T��x��� ��!�3��G,{� Pbt��C�� ��/�:/L/^/ p/�/���	/�/ =?$?6?H?Z?)/~? �?�?�?�/�?k?�?O  O2ODO�/�/�/�/�? �O�/�O�O�O
__�? @_R_d_v_�_�O-_�_ �_�_�_oUOgOyO�O �_ro�O�o�o�o�o�o �_&8Jmo�o �����o)o;o MoO!��oX�j�|��� ��oď֏����/����B�T�f�x���^�S�T_ERR J�;�����PDUSI�Z  ��^P�����>ٕWRD �?z���  �guest ���+�=�O�a�s�*��SCDMNGRPw 2Kz�Ð���۠\��K��� 	P01.�14 8�q  � y��B    ;�����{ �����������������������~ �ǟI�4�m�X��|��  i�  �  
����� ����+��������
����l�.x��
��"�l�ڲ۰s��d�������_G�ROU��L�� e��	��۠07K�QUPD  ����PČ�TYg������TTP_A�UTH 1M��� <!iPen'dan���<�_��!KAREL�:*�����KC�%�5�G��VISION SETZ���|��Ҽߪ��� ������
�W�.�@����d�v���CTRL� N�������
��FFF9E�3���FRS:DEFAULT��FANUC �Web Server�
������q�������������W�R_CONFIGw O�� ����IDL_CPU�_PC"��B���= �BH#MI�N.�BGNR_�IO��� ���% N�PT_SIM_D�Os}TPMO_DNTOLs �_PRTY�=!OLNK 1P���'9K]|o�MASTEr ������O_CFG���UO����C�YCLE���_?ASG 1Q���
 q2/D/V/h/ z/�/�/�/�/�/�/�/p
??y"NUM����Q�IPCH���£RTRY_�CN"�u���SC�RN������ ���R����?���$J23_D_SP_EN������0OBPROC��3��JOGV�1�S_�@��8��?�';ZO'??0CP�OSREO�KANJI_�Ϡu�A$#��3T ���E�O�ECL_LM B2e?��@EYLOGGI�N�������L�ANGUAGE Y_�=� }Q���LG�2U������ �x�����PZC � �'0������MC:\RSCH\00\˝�LN_DISP V�������T�OC�4Dz\A��SOGBOOK W+��o���o�o���Xi�o�o�o�o��o~}	x(y��	�ne�i�ekElG�_BUFF 1X���}2���� Ӣ������'� T�K�]����������� ɏۏ���#�P���~�qDCS Zxm =���%|d1h�`���ʟܟ�g�IOw 1[+ �?'����'�7�I�[�o� �������ǯٯ��� �!�3�G�W�i�{��������ÿ׿�El TM  ��d��#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U��g�yߋߝ߈t�SE�V�0m�TYP�� ��$�}�A�RS"�(_�s�2FLg 1\��0��� �����������5�STP<P���DmNGNAM�4�U�nf�UPS`GI�5��A�5s�_LOA�D@G %j%=@_MOV�u�����MAXUALRMB7�P8��y���3��0]&q��Ca]�s�3�~�� 8@=@^�+ طv	��V0+�P�A5d�cr���U� �����E( iTy����� ��/ /A/,/Q/w/ b/�/~/�/�/�/�/�/ ??)?O?:?s?V?�? �?�?�?�?�?�?O'O OKO.OoOZOlO�O�O �O�O�O�O�O#__G_ 2_D_}_`_�_�_�_�_ �_�_�_o
ooUo8o yodo�o�o�o�o�o�o��o�o-��D_LDXDISA^�� �MEMO_APX��E ?��
 �0y�����������ISC ;1_�� �O� ���W�i�����Ə �����}��ߏD�/� h�z�a��������� �����@���O�a� 5������������u� �ׯ<�'�`�r�Y��� ���y�޿�ۿ��� 8Ϲ�G�Y�-ϒ�}϶� ������m�����4���X�j�#�_MSTR� `��}�SCD 1as}�R���N� �������8�#�5�n� Y��}��������� ���4��X�C�|�g� �������������� 	B-Rxc�� �����> )bM�q��� ��/�(//L/7/ p/[/m/�/�/�/�/�/ �/?�/"?H?3?l?W?��?{?�?�?�?n�MK�CFG b����?��LTARM_��2cRuB� �3WpTNBpME�TPUOp�2�����NDSP_CM�NTnE@F�E�� d���N�2A�O|�D�EPOSCF�G��NPSTOL �1e-�4@�<#�
;Q�1;UK_YW7_ Y_[_m_�_�_�_�_�_ �_o�_oQo3oEo�o�io{o�o�a�ASIN�G_CHK  ��MAqODAQ2Cf�O�7J�eDEV �	Rz	MC:>'|HSIZEn@�����eTASK �%<z%$1234?56789 ��u��gTRIG 1g.�� l<u%����3���>svvYP�aq��kEM_IN�F 1h9G� `)AT?&FV0E0(����)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏ P��t�������]�ί �����(�۟�^� �#�5�����k�ܿ�  ϻ�ů6��Z�A�~� ��C���g�y������ ��2�i�C�h�ό�G� ���ߩ��ߙϫ���� ����d�v�)ߚ��߾� y��������<�N� �r�%�7�I�[���� ��9�&��J[��g��>ONIT�OR�@G ?;{ �  	EXESC1�3�2�3�E4�5��p�7�8�9�3�n�R �R�RRR R(R4R@RTLR2Y2e2qU2}2�2�2�U2�2�2�3Y�3e3��aR_G�RP_SV 1i�t��q(�5�
���5��۵MO�~q_DCd~�1PL�_NAME !�<u� �!De�fault Pe�rsonalit�y (from �FD) �4RR2�k! 1j)TEX�)TH��!�AX d�?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�Ox2-?�O�O�O__0_ B_T_f_x_�b<�O�_ �_�_�_�_�_o o2o�DoVoho&xRj" 1�o�)&0\�b, Ӗ9��b�a @oD�  �a?��c�a?�`�a�aA'��6�ew;�	l��b	 �xoJp��`��`	p �<; �(p� �.r� �K�K ���K=*�J���J���JV��k0q`q�P�x�|�� @j�@T;f�r�f�q�ac^rs�I�� ��p����p�r�ph}�3��´  ���>��ph�`z���꜖"�Jm�q� H�N��a`c��$�dw��  ��  P� Q�� �� |  ��m�Əi}	'� �� �I� �  �����:�È�È=G���(��#�a	����I  �n @H�i~�ab�Ӌ�b!�$w���"N0���  'Ж�q�p@2��@����r��q5�C�pC0C��@ C�����`
�A1]w@�B�V~X�
nwBD0h�A��p�ӊ�p@����aDz���֏࿯�Я	�pv�(� �� -���I��-�=��A�a��we_q�`�p �??�ff ��m�|�� �����Ƽ�!@ݿ�>1�  P�apv(�`ţ�� �=�qst��?˙��`x`�� <
�6b<߈;����<�ê<�? <�&P�ς��AO��c1��ƍ�?offf?O�?&���qt@�.�J<?�`��wi4� ���dly�e߾g;ߪ� t��p�[ߔ�߸ߣ� ���� ����6�wh�F0%�r�!�����1ى����E��� E�O�G+� F�!���/���?�e�`P���t���lyBL�cB��Enw4������� +��R��s���������h�yÔ�>���I�mXj���A�y�weC��������#/*/c/�N/wi�����v/C�`� CHs/`
=$��p�<!�!��ܼ�'��3A�A�AR�1AO�^?��$�?������
=ç>�����3�W
=�s#�]�;e��?������{�����<�>(��B�u���=B0�������	R��zH�F��G���G���H�U`E����C�+��}I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*O ONO9OrO]O�O�O�O �O�O�O�O_�O8_#_ \_G_�_�_}_�_�_�_ �_�_�_"oooXoCo |ogo�o�o�o�o�o�o �o	B-fQ� u������� ,��P�b�M���q��� ��Ώ���ݏ�(�� L�7�p�[������ʟ ���ٟ���6�!�Z��E�W���#1( �ٙ9�K���ĥ ������Ư!3��8���!4Mgqs��,�IB+8��J��a���{�d�d�����ȿ��쿔ڼ%P8�P�= :GϚ�S�6�h�z���R�Ϯ����������  %�� ��h� Vߌ�z߰�&�g�/9�$�������7�����A�S�e�w�   ������������̿2 F�$�&Gb��������!C���@���8������F� Dz�N�� F�P �D�������)#�B�'9K]o#?_���@@v
4$�8�8��8�.
 v��� !3EWi{�����:� ���ۨ�1��$M�SKCFMAP � ���� ���(.�ONREL  ��!9��EXC/FENBE'
#7%�^!FNCe/W$JO�GOVLIME'dtO S"d�KEYE'u�%�RUN�,��%�SFSP�DTY0g&P%9#S�IGNE/W$T1M�OT�/T!�_C�E_GRP 1p��#\x��?p� �?�?�?�?�?O�? OBO�?fOO[O�OSO �O�O�O�O�O_,_�O P__I_�_=_�_�_�_ �_�_oo�_:o��TCOM_CFG 1q	-�vo�o��o
Va_ARC_�b"�p)UAP_�CPL�ot$NOCHECK ?	+ �x�% 7I[m���������!�.+N�O_WAIT_L� 7%S2NT^ar�	+�s�_ERR�_12s	)9��  ,ȍޏ��x����&��dT_MO��t>��, *oq��9�PARAM��u	+��a�ß'g�{�� =?�345?678901�� ,��K�]�9�i�����`��ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDS�P�c#6p(OFFSET_CART�oη�DISƿ��PE?N_FILE尨!��ai��`OPTIO�N_IO�/��PW�ORK ve7s# ��V�ؤ�p�p�4�p�	 ����p��<���RG_DSBL  ���P#��ϸ�RIE�NTTOD ?�Cᴭ !l�UT__SIM_D$�"����V��LCT w}�h�iĜa[�1ԟ_PEXE�j�R�ATvШ&p%� ��2�^3j)TEX)T�H�)�X d 3�������%�7�I� [�m��������������!�3�E���2 ��u���������������c�<d�AS ew������`��Ǎ�^0OUa0�o(��(�����u2, ����O H @D��  [?�aG?��cc�D][�Z��;�	ls��xJ��������<� ��� ���2�H(��H3�k7HSM5G��22G���Gpc
͜�'f�/,-,2�CR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t3�!�/ �/�"�t32����/6 W ��P%�Q%��%�|T��S62�q?�'e	'� � ��2I� � � ��+==�̡ͳ?�;	�h	�0��I  �n �@�2�.��Ov;���ٟ?&gN�]O  �''�uD@!� C�C��@F#H!�/�O�O Nsb
���@�@E��@�e`0B��QA�0Yv: �13Uwz$oV_�/z_�e_�_�_	��( �� -�2@�1�1ta�Ua�c����:A-���.  �?�ff���[o"o�_!U�`oXÜQ8���o:�j>�1  Po�V(���eF0�f�Y����L�?����x�b�P<
6b<�߈;܍�<��ê<� <�#&�,/aA�;r��@Ov0P?fff?��0?&ip�T@�.�{r�J<?�`�u#	�Bdqt�Yc �a�Mw�Bo�� 7�"�[�F��j����� ��ُ����3�����,���(�E��� E��3G+� F��a��ҟ������,��P�;���B�pAZ�>��B��6�<O ίD���P��t�=����a�s�����6j�h�y�7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�<%?��?������(���#	Ę��P �N�||CH���Ŀx������@I�_��'�3A�A�A�R1AO�^??�$�?��� ��±
=ç>�����3�W
=�#� U��e����B��@��{�����<����(�B�u���=B0�������	�b�H��F�G���G���H�U`E����C�+��I�#�I��H�D�F��E��RC�j=[��
I��@H��!H�( E?<YD0߻� �������� �9�$� ]�H�Z���~������� ������#5 YD }h������ �
C.gR� ������	/� -//*/c/N/�/r/�/ �/�/�/�/?�/)?? M?8?q?\?�?�?�?�? �?�?�?O�?7O"O[O mOXO�O|O�O�O�O�O��O�O�O3_Q(���3���b��gUU���W_i_2�3ǭ8��_�_2�4M�gs�_�_�RIB+��_�_�a���{�miGo5okoYo(�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�u�,��  �p���o ��/��S��z
uү ܠ�������ڱ������������  /�M�w�e�������~�l2 F�$��'Gb��t��a�`�,p�S�C�y�@p�5��G�Y�۠F� D�z�� F�P D��]����پ��ʯܯ� ��~ÿ?���@@�J?�K�K���K���
 �|��� ����Ŀֿ������0�B�T�fϽ�V� ����{��1��$�PARAM_ME�NU ?3���  �DEFPULS�Er�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L��	�OPT���PTB4�.�C��R_DECSN ���e��ߑߣ����� ������!�3�\�W��i�{���USE_PROG %��q%�����CCR����e����_HOSoT !��!��:���T�`�V��/��X����_TIMqE��^��  ��?GDEBUG\�����GINP_FL'MSK����Tfp�����PGA  ��̹�)CH����TY+PE������� ����� - ?hcu���� ���//@/;/M/ _/�/�/�/�/�/�/�/��/??%?7?`?��W�ORD ?	=�	RSfu	P�NSUԜ2JO�K�DRTEy�]T�RACECTL �1x3��� }�` &�`��`�>�6DT Q�y3�%@�0D �� �c��a:@V�@BR�2ODOVOhO�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V�.Iv��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p��j�����  $6HZl~ �������/  /2/D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o��o 0BTfx��� ������,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l�~� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ����������*��$�PGTRACEL�EN  )�  ��(���>�_UP z/���m�u�Y��n�>�_CFG7 {m�W�(��~���PКӂ�DEFSPD |���'�P��>�IN~��TRL }���(�8����PE__CONFI��~m՟�mњ�\�ղ�LID�����=�GRP 1���W��)�A ����&ff(�A�+33D�� D�]� CÀ A)@1��Ѭ(�d�Ԭ����0�0�� 	 �1�ح֚��� �������B�9�����O�9�s�(�>�?T?�
5��������� =��=#�
����P ;t_�����<��  Dz (�
H�X~i ������/��/D///h/S/�/���
V7.10be�ta1��  �A�E�"ӻ�A (�� ?!G���!>���"�܇��!���!BQ��!A\� �!��T�!2p����Ț/ 8?J?\?n?};� ����/��/�?}/�?�? OO:O%O7OpO[O�O O�O�O�O�O�O_�O 6_!_Z_E_~_i_�_�_ �_�_�_�_'o2o�_ VoAoSo�owo�o�o�o �o�o�o.R=�v1�/�#F@  �y�}��{m��y=� �1�'�O�a��?�?�? ������ߏʏ��'� �K�6�H���l����� ɟ���؟�#��G� 2�k�V���z������� �o��ίC�.�g� R�d����������п 	���-�?�*�cώ� ��Ϯ������ B�;�f�x�������D� ���߶��������7� "�[�F�X��|��� ��������!�3��W� B�{�f��������� � ����/S>w bt������ =OzόϾψ ����ϼ� /.�'/ R�d�v߈߁/0�/�/ �/�/�/�/�/#??G? 2?k?V?h?�?�?�?�? �?�?O�?1OCO.OgO RO�OvO�O�O���O�O �O__?_*_c_N_�_ r_�_�_�_�_�_o�_ )oTfx�to�� �/�o/>/P/ b/t/mo�|�� �����3��W� B�{�f�x�����Տ�� �����A�S�>�w� b����O��џ����� �+��O�:�s�^��� ����ͯ���ܯ�@o Rodo�o`��o�o�o�� ƿ�o���*<N� Y��}�hϡό��ϰ� �������
�C�.�g� Rߋ�v߈��߬����� 	���-��Q�c�N�� �����l������� �;�&�_�J���n��� ��������,�>�P� :L��������� ���(�:�3��0 iT�x���� �/�///S/>/w/ b/�/�/�/�/�/�/�/ ??=?(?a?s?��? �?X?�?�?�?�?O'O OKO6OoOZO�O~O�O �O�O�O*\&_8_�r���_�_��$�PLID_KNO�W_M  ��� Q�TSoV ���P��?o"o 4o�OXoCoUo�o R��SM_GRP 1���Z'0{`�@R�`uf�e�`
�5 � �gpk' Pe]o�����������SMR��c��mT�EyQ}? yR����������� ����ӏ�G�!��-� ����������韫��� ϟ�C���)������������寧���QS�T�a1 1���)���P0� A 4��E2�D�V�h��� ����߿¿Կ���9� �.�o�R�d�vψ���P�Ͼ����2�0�N Q�<3��3�/�A�S��4l�~ߐ����5���������A6
��.�@��7Y�k�}���8���������MAD  �)��PAR�NUM  !��}o+��SCHE� �S�
��f���S��UPDf�x��_CMP_�`H�� ��'�UER_wCHK-���ZE*<RSr��_�QG_MOG���_�~X�_RES_G��!���D�>1 bU�y������/�	/��� �+/�k�H/g/l/� �Ї/�/�/�	��/�/ �/�X�?$?)?��� D?c?h?����?�?�?�V 1��U�ax�@c]�@t@(�@c\�@�@D�@c[�*@��T?HR_INRr�J���b�Ud2FMASS6?O ZSGMN>OqC�MON_QUEUE ��U�V P~P� X�N$ UhN8�FV�@END�A���IEXE�O�E��B�E�@�O�COPTI�O�G��@PROG�RAM %�J%��@�?���BTAS�K_IG�6^OCFG ��Oz��_�P�DATA�c��[@Ц2=�DoVoho zo�j2o�o�o�o�o�o�);M jIN+FO[��m��D �������� 1�C�U�g�y����������ӏ���	�dwpt��l )�QE DI�T ��_i��^W�ERFLX	C�RGADJ �tZA�����?נʕFA~��IORITY�G�W���MPDSP(NQ����U�GD��oOTOE@1�X� (!AF:@�E� c�Ч!t�cpn���!u�d����!icm����?<�XY_�Q�X���Q)� a*�1�5��P�� ]�@�L���p������� �ʿ��+�=�$�a��Hυϗ�*��POR�T)QH��P�E���_CARTRE�PPX��SKSTyA�H�
SSAV�@��tZ	2500H863���_x�
Ԫ'��X�@�s�wPtS�ߕߧ���UR�GE�@B��x	WFF��DO�F"[W\��������WRUP_�DELAY �|X���R_HOTqX�	B%�c���R_NORMALq^R��v�SEMI�����9�QSKIP'��vtUr�x 	7� 1�1��X�j�|�?�tU �������������� $J\n4�� ������4 FX|j��� ����/0/B//�R/x/f/�/�/�/tU�?$RCVTM$��D��� DCR'����Ў!?��L�B�'�CE��>�x�=���8.(gC�����e��ߠ��?����:�o?��� <
6b<�߈;܍�>�u.�?!<�&�?h?�?�?�@ >��?O O2ODOVOhO zO�O�O�O�O�O�?�O �O__@_+_=_v_Y_ �_�_�?�_�_�_oo *o<oNo`oro�o�o�o �_�o�o�o�o�o8 J-n��_��� ����"�4�F�X� j�U������ď��� ӏ���B�T��x� ��������ҟ���� �,�>�)�b�M����� �������ïկ�Y� :�L�^�p��������� ʿܿ� ����6�!� Z�E�~ϐ�{ϴϗ��� ��-�� �2�D�V�h� zߌߞ߰��������� 
���.��R�=�v�� k���������� *�<�N�`�r������� ���������& J\?����� ���"4FX�j|��!GN_A�TC 1�	; �AT&FV�0E0�AT�DP/6/9/2{/9�ATA��,AT%G�1%B960��+++�,�H�/,�!IO_TY�PE  �%�#�t�REFPOS�1 1�V+ x�u/�n�/j �/
=�/�/�/Q?<?u? ?�?4?�?X?�?�?�+/2 1�V+�/�?��?\O�?�O�?�!3 1�O*O<OvO�O�O|_�OS4 1��O��O�O_�_t_�_+_S5 1�B_T_f_�_�o	oBo�_S6 1��_�_�_5o�o�o�o>UoS7 1�lo~o��o�oH3l�oS8 1�%_����SMASKw 1�V/  
?��M��XNOS/�r�������!MOTE�  n��$��_CFG ����q���"PL_RANG������POWER ������SM�_DRYPRG �%o�%�P��T?ART ��^�UME_PRO-��?����$_EXEC_ENB  ���GSPD��Րݘ���TDB��
�R�M�
�MT_'�T�����OBOT�_NAME �o����OB_O�RD_NUM ?��b!H?863  �կ����PC_TIMEOUT��{ x�S232Ă�1�� L�TEACH PE�NDAN��w���-��Mai�ntenance Cons���s��"���KCL/!Cm��

���t�ҿ� No Us�e-��Ϝ�0�NPqO�򁋁���.�CH_L�������q	��s�MAVAIL������糅��SPACE�1 2��, �j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��ߤ� �ߚ� �2�D���h� ��|��`������ ���� �2�D��h� ��|���`���������y���2����0� B���f�����{���3); M_����� �/� /44F Xj|*/���/�/@�/?(??=?5Q/ c/u/�/�/G?�/�/�?�O�?$OEO,OZO6 n?�?�?�?�?dO�?�? _,_�OA_b_I_w_7�O�O�O�O�O�_�O _(oIoo^oofo�o8�_�_�_�_�_�o o6oEf){����G �o�� ���
M� ���*�<�N�`�r� ������w���o������d.��%�S� e�w�����������Ǐ َ���Θ8�+�=�k� }�������ůׯ͟�� ��%�'�X�K�]��� ������ӿ�����p�#�E�W� `� @�������x�����\�e������ �����R�d߂�8�j� �߾߈ߒߤ������ ����0�r���X�� ����������8�����
�ύ�_MO�DE  �{��S ��{|�2�0�A����3�	S�|)CWORK_{AD���K�+/R  �{�`� ��� _INTVA�L���d���R_O�PTION� ���H VAT_G�RP 2��up(N�k|��_�� ���/0/B/��h� u/T� }/�/�/�/�/ �/�/?!?�/E?W?i? {?�?�?5?�?�?�?�? �?O/OAOOeOwO�O �O�O�OUO�O�O__ �O=_O_a_s_5_�_�_ �_�_�_�_�_o'o9o �_Iooo�o�oUo�o�o �o�o�o�o5GY k-���u�� ���1�C��g�y� ��M�����ӏ叧�	� �-�?�Q�c������� ��������ǟ��;�M�_����$SC?AN_TIM��_%�}�R �(�#((�<04_d d 	
!D�ʣ���u�/������U��25���@�dD5�P�g��]	����������dd�x� � P���� ��  8� ҿ�<!���D��$�M� _�qσϕϧϹ���������ƿv���F�X��/� ;��ob��pm��t�_DiQ|̡  � l� |�̡ĥ�������!� 3�E�W�i�{���� ����������/�A� S�e�]�Ӈ������� ������);M _q������ �r���j�Tf x������� //,/>/P/b/t/�/��/�/�/�/�%�/  0��6��!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O*�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo�O�OJ�o�o�o �o�o�o�o 2D Vhz�����`��
�7?  ;� >�P�b�t��������� Ǐُ����!�3�E��W�i�{�������ß �ş3�ܟ��&� 8�J�\�n�������������ɯ�����,� �+�	�12345678^�� 	� =5���f�x�������������
��.�@� R�d�vψϚ�៾��� ������*�<�N�`� r߄߳Ϩߺ������� ��&�8�J�\�n�� ������������� "�4�F�u�j�|����� ����������0 _�Tfx���� ���I>P bt������ �!/(/:/L/^/p/��/�/�/�/�/�/� 2�/?�#/9?K?]?��iCz  Bp�˚   ��h2���*�$SCR_�GRP 1�(��U8(�\x�d�@ >� �'��	  �3�1�2�4(1*�&�I�3�F1OOXO}m��D�@�0ʛ)����HUK�LM-�10iA 890�?�90;��F;�M61C D�:�CP�*�1
\&V�1	��6F��CW�9)A7Y	�(R�_�_�_�_�_�\���0i^�oO UO>oPo#G�/���o�'o�o�o�o�oB�B0�rtAA�0*  @�Bu&Xw?��ju�bH0{Uz�AF@ F�` �r��o����� +��O�:�s��mBqrr`����������B�͏ b����7�"�[�F�X� ��|�����ٟğ���N����AO�0�B�CU
�L���E�jqBq=���Ҕ�$G@�@pϯ B���G�I
E��0EL_DEFA�ULT  �T�_�E���MIPOWERFL  
E*��7�oWFDO� *���1ERVENT �1���`(��� L!DUM_�EIP��>��j!AF_INE�<¿C�!FT�������!o:� ���a�!RPC�_MAINb�DȺ8Pϭ�t�VIS}�C�y�����!TP���PU�ϫ�d��E�!�
PMON_PR'OXYF߮�e4ߑ���_ߧ�f����!RDM_SRV��r��g��)�!R�dIﰴh�u�!
v��M�ߨ�id���!?RLSYNC��>��8���!ROS��4��4��Y�(� }���J�\��������� ����7��["4 F�j|�����!�Eio�ICE_KL ?%�� (%SVCPRG1n>���3D��3���4/D/�5./3/�6V/[/�7~/�/��D�/�9�/�+�@��/ ��#?��K?�� s?� /�?�H/�?� p/�?��/O��/;O ��/cO�?�O�9? �O�a?�O��?_� �?+_��?S_�O{_ �)O�_�QO�_�yO �_��Os���� >o�o}1�o�o�o�o�o �o�o;M8q \������� ��7�"�[�F��j� ������ُď���!� �E�0�W�{�f����� ß���ҟ���A� ,�e�P���t���������ί�y_DEV� ��M{C:�@`!�OUT��2��?REC 1�`e��j� �� 	 �����˿���ڿ��
 �`e��� 6�N�<�r�`ϖτϦ� �Ϯ�������&��J� 8�n߀�bߤߒ��߶� ������"��2�X�F� |�j���������� ����.�T�B�x�Z� l������������� ,P>`bt� �����( L:\�d��� �� /�$/6//Z/ H/~/l/�/�/�/�/.� �/?�/2? ?V?D?f? �?n?�?�?�?�?�?
O �?.O@O"OdORO�OvO �O�O�O�O�O�O__ <_*_`_N_�_�_x_�_ �_�_�_�_oo8oo ,ono\o�o�o�o�o�o �o�o�o "4j X������� ���B�$�f�T�v� �����������؏� �>�,�b�P�r���p�oV 1�}� P
��ܟ� ���TY�PE\��HELL_CFG �.�z�͟  	�<����RSR���� ��ӯ�������?� *�<�u�`��������������  �%�3�E��Q̊\���M�o�p�)�d��2��d]�KϾ:�HK 1�H� u�������A� <�N�`߉߄ߖߨ��� ��������&�8��~=�OMM �H����9�FTOV_E�NB&�1�OW_?REG_UI��8��IMWAIT��\a���OUT�������TIM������VAL����_U�NIT��K�1�MO�N_ALIAS �?ew� ( he�#������������ ��);M��q� ���d�� %�I[m�< ������!/3/ E/W//{/�/�/�/�/ n/�/�/??/?�/S? e?w?�?�?F?�?�?�? �?�?O+O=OOOaOO �O�O�O�O�OxO�O_ _'_9_�O]_o_�_�_ >_�_�_�_�_�_�_#o 5oGoYokoo�o�o�o �o�o�o�o1C �ogy��H�� ��	��-�?�Q�c� u� �������ϏᏌ� ��)�;��L�q��� ����R�˟ݟ��� ��7�I�[�m��*��� ��ǯٯ믖��!�3� E��i�{�������\� տ�����ȿA�S� e�wω�4ϭϿ����� �����+�=�O���s� �ߗߩ߻�f������ �'���K�]�o��� >����������#� 5�G�Y��}����������o��$SMON�_DEFPRO ������� *S�YSTEM*  �d=��RECA�LL ?}�� �( �}3cop�y frs:or�derfil.d�at virt:�\tmpback�\=>inspi�ron:2636`��r��o�}*.mdb:*.*C�U
Y���	.x.:\�8R�n(���/.a6H _^�//�-? Qb/t/�/�/�F/� �/�/??)�M�/ p?�?�?�8?J?��?� OO�%
xyzrate 61 �?@�?�?nO�O�O�%.G>R(4940 HOZO �O�O_"/4/�/�Ga_ s_�_�_�/E_�HY_�_ �_o!?3?FO�C�_no �o�o�?6oHo�@^o�o &O8O�o�omx��O�J8124�O Y���!3s����n�������I2488G�Y�����!_ 3_�_��a�s������_ E���Y�����!o3o Fݟn������o6� H�ŀ^����&�8� ��ܟm��������ȟ Z�����"�4�ǯX� i�{ύϠ���C�֯�� ����0�B�T�e�w� �ߜ���I�ҿ����� �,Ͽ�P�a�s��� ��;���`�����(�������o����������� 13164  I�[�����#�5������fx�����A 8028HZ��"�4.�@߸bt�� }+��I�Z ��/��4�G���o/�/�/&�0��?/�
 _/�/??'9�� n?�?�?��/�[?�?��?O!��$SNP�X_ASG 1�����9A�� P 0 �'%R[1]�@1.1O �?�$�%dO�OsO�O�O�O �O�O�O __D_'_9_ z_]_�_�_�_�_�_�_ 
o�_o@o#odoGoYo �o}o�o�o�o�o�o�o *4`C�gy �������	� J�-�T���c������� ڏ�����4��)� j�M�t�����ğ���� ��ݟ�0��T�7�I� ��m��������ǯٯ ���$�P�3�t�W�i� �������ÿ���� :��D�p�Sϔ�wω� �ϭ��� ���$��� Z�=�dߐ�sߴߗߩ� ������ ��D�'�9� z�]��������� 
����@�#�d�G�Y� ��}������������� *4`C�gy ������	 J-T�c��� ���/�4//)/ j/M/t/�/�/�/�/�/��/�/?0?4,DPA�RAM �9E}CA �	��:�P�4�0$HOF�T_KB_CFG�  q3?E�4PI�N_SIM  9K�6�?�?�?�0,@�RVQSTP_DSB�>�21On8J0�SR ��;� G& =O{Oq0�6�TOP_ON_E_RR  q4�9~�APTN �5��@A�BRING_PRM�O� J0VDT_G�RP 1�Y9�@  	�7n8_(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2Dkhz �������
� 1�.�@�R�d�v����� ����Џ�����*� <�N�`�r��������� ̟ޟ���&�8�J� \�����������ȯگ ����"�I�F�X�j� |�������Ŀֿ�� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�tߛߘߪ� ����������(�:� a�^�p������� ���� �'�$�6�H�Z� l�~���������������3VPRG_CO7UNT�6��A�5NENB�OM=��4J_UPD 1}��;8  
 q2������  )$6Hql~� ����/�/ / I/D/V/h/�/�/�/�/ �/�/�/�/!??.?@? i?d?v?�?�?�?�?�? �?�?OOAO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_��_�_YSDEBSUG" � �Pdk	��PSP_PASS�"B?�[LOG� ��mr�P�X�_  �g~�Q
MC:\d<�_b_MPCm�H�o�o�Qa�o �~vfSAV �m�:dUb�U\gS�V�\TEM_TI�ME 1�� �(�P[�TZ�o	T1SVGUNS} �#'k�spAS�K_OPTION�" �gospBC?CFG ��|c �b��z`� ���4��X�C�|�g� ����ď֏������ 	�B�-�f�Q�c����� �����ϟ��,�>�)�b��YR���S��� ƯA������ ��D� �nd��t9�l������� ��ڿȿ�����"� X�F�|�jϠώ��ϲ� ��������B�0�f� T�v�xߊ��ߦؑ��� ����(��L�:�\� ��p���������� � �6�$�F�H�Z��� ~������������� 2 VDzh�� �������4 Fdv���� ��//*/�N/</ r/`/�/�/�/�/�/�/ �/??8?&?\?J?l? �?�?�?�?�?�?�?�? OO"OXOFO|O2�O �O�O�O�OfO_�O_ B_0_f_x_�_X_�_�_ �_�_�_�_oooPo >otobo�o�o�o�o�o �o�o:(^L np�����O� �$�6�H��l�Z�|� ����Ə؏ꏸ���� 2� �V�D�f�h�z��� ��ԟ����
�,� R�@�v�d��������� ίЯ���<��T� f�������&�̿��ܿ ��&�8�J��n�\� �π϶Ϥ�������� ��4�"�X�F�|�jߌ� �ߠ����������� .�0�B�x�f��R��� ���������,��<� b�P�������x����� ����&(:p ^�������  6$ZH~l ��������/ &/D/V/h/��/z/�/��/�/�/�&0�$T�BCSG_GRP� 2��%��  �1 
? ?�  /?A? +?e?O?�?s?�?�?�?��?�;23�<d�, �$A?1	� HC���6>�@E�5CL  �B�'2^OjH4Jݸ�B\)LFY g A�jO�MB��?F�IBl�O�O�@�JG|_�@�  D	�15_ __$YC-P{_F_$`_j\��_�]@0�> �X�Uo�_�_6oSoo�0o~o�o�k�h�0	V3.00'2�	m61c�c	�*�`�d2�o�e>əJC0(�a�i �,p�m-  �0�����omvu1JC�FG ��%� 1 #0vz��r8Br�|�|��� �z� �%��I�4�m� X���|��������֏ ���3��W�B�g��� x�����՟������ ��S�>�w�b����� '2A ��ʯܯ����� �E�0�i�T���x��� ÿտ翢����/�� ?�e�1�/���/�Ϝ� ���������,��P� >�`߆�tߪߘ��߼� �������L�:�p� ^����������� � �6�H�>/`�r�� ��������������  0Vhz8�� ����
.� R@vd���� ���//</*/L/ r/`/�/�/�/�/�/�/ �/�/?8?&?\?J?�? n?�?�?�?�?���?O O�?FO4OVOXOjO�O �O�O�O�O�O__�O B_0_f_T_v_�_�_�_ z_�_�_�_oo>o,o boPoroto�o�o�o�o �o�o(8^L �p������ �$��H�6�l�~�(O ����f�d��؏��� 2� �B�D�V������� n����ԟ
���.�@� R�d����v������� �Я���*��N�<� ^�`�r�����̿��� ޿��$�J�8�n�\� �π϶Ϥ�������� ��(�:�L���|�jߌ� �ߠ����������0� B�T��x�f���� ���������,��P� >�t�b����������� ����:(JL ^������  �6$ZH~l ��^���dߚ / /D/2/h/V/x/�/�/ �/�/�/�/�/?
?@? .?d?v?�?�?T?�?�? �?�?�?OO<O*O`O NO�OrO�O�O�O�O�O _�O&__6_8_J_�_ n_�_�_�_�_�_�_�_ "ooFo��po�o,o Zo�o�o�o�o�o0 Tfx�H�� �����,�>�� b�P���t��������� Ώ��(��L�:�p� ^�������ʟ���ܟ � �"�$�6�l�Z��� ~�����دꯔo�� &�ЯV�D�z�h����� ��Կ¿��
��.���R�@�v�dϚτ�  9���� ��������$TBJOP_GRP 2ǌ���  �?������������x�JBЌ��9� �< �X�=��� @���	 �C�� t�b  C���я>��͘Րդ�>�̚йѳ33=�CLj�fff}?��?�ffBGР�ь�����t�ц�>w�(�\)�����E噙�;���hCYj��  @�h��B�  A�����f��C�  �Dhъ�1��O��4�N����
:_���Bl^��j��i�l�l����Aəg�A�"��D���֊=qH���н�p�h�Q�;��A�j�ٙ�@L��D	2�����x��$�6�>B�\���T���Q�tsx�@�33@���C����y�1����>�#�Dh�����������<{�h�@ i� ��t��	 ���K&�j �n|���p�@/�/:/k/�ԇ����!��	V3.�00J�m61cI�*� IԿ��/�'� Eo�E���E��E��F��F�!�F8��F�T�Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G�,I�!CH`��C�dTDU�?�D��D��D�E(!/E\��E��E�h��E�ME��s�F`F+'\�FD��F`=�F}'�F���F�[
F����F��M;��;Q��T,8�4` *(�ϴ?�2���3\��X/O��ESTPARS  ��	����HR@ABLE K1����0��
H��7 8��9
G
HP
H����
G	
H

HQ
HYE��
H
Hu
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_$�^:BS _� �JGo Yoko}o�o�o�o�o�o �o�o1CUg y����`#oRL�y �_�_�_�_�O�O�O�O��OX:B�rNUM [ ���P���� V@P:B_CFG ˭�Z�h��@��IMEBF_�TT%AU��2@�V�ERS�q��R� 1���
 ($�/����b� ���� J�\���j�|���ǟ�� ȟ֟�����0�B��T���x�������2�_ԧ��@�
��MI__CHAN�� �} ��DBGLV����������ETHERAD ?��O�������h������ROUT��!��!������SNMASKD��U�255.���#������OOLOFS�_DI%@�u.�O�RQCTRL �����}ϛ3rϧϹ� ��������%�7�I߀[�:���h�z߯�APE_DETAI"��G�PON_SVO�FF=���P_MOON �֍�2���STRTCHK ��^�����VT?COMPAT��O������FPROG �%^�%GET�DAT����9�P�LAY&H��_IN�ST_Mް �������US�q��L�CK���QUIC�KME�=���SC�REZ�G�tps� ���u�z�����_��@@n�.�S�R_GRP 1о^� �O� ���
��+O=sa�쀚�
m�� ����L/C 1gU�y��� ��	/�-//Q/?/�a/�/	1234�567�0�/�/@X�t�1���
 �}�ipnl/� g?en.htm�?� ?2?D?V?`P�anel setupZ<}P�?�?�?�?�?�? �??,O >OPObOtO�O�?�O!O �O�O�O__(_�O�O ^_p_�_�_�_�_/_]_ S_ oo$o6oHoZo�_ ~o�_�o�o�o�o�o�o so�o2DVhz� 1'���
�� .��R��v��������ЏG���UALR�M��G ?9� �1�#�5�f�Y��� }�������џן����,��P��SEV � ����E?CFG ������A��   BȽ�
 Q���^� ���	��-�?�Q�c�@u�������������C �����I��?���(%D�6� � $�]�Hρ�lϥϐ��� ��������#��G����� �߿U�I_�Y�HIST 1վ�  (��� ��,/SOF�TPART/GE�NLINK?cu�rrent=editpage,��,1����,�;��� ����menu��962�߆���0��K�]�o�36u�
� �.�@���W�i�{��� ������R����� /A��ew��� �N��+= O�s��������f��f//'/ 9/K/]/`�/�/�/�/ �/�/j/�/?#?5?G? Y?�/�/�?�?�?�?�? �?x?OO1OCOUOgO �?�O�O�O�O�O�OtO �O_-_?_Q_c_u__ �_�_�_�_�_�_�� )o;oMo_oqo�o�_�o �o�o�o�o�o%7 I[m� �� �����3�E�W� i�{������ÏՏ� ������A�S�e�w� ����*���џ���� �ooO�a�s����� ����ͯ߯���'� ��K�]�o��������� F�ۿ����#�5�Ŀ Y�k�}Ϗϡϳ�B��� ������1�C���g� yߋߝ߯���P����� 	��-�?�*�<�u�� ������������ )�;�M���������� ������l�%7 I[������ �hz!3EW i������� v////A/S/e/P����$UI_PA�NEDATA 1������!�  	�}�w/�/�/�/�/?? )?>?��/i?{?�? �?�?�?*?�?�?OO OAO(OeOLO�O�O�O��O�O�O�O�O_&Y� b�>RQ?V_h_ z_�_�_�__�_G?�_ 
oo.o@oRodo�_�o oo�o�o�o�o�o�o *<#`G��}�-\�v�#�_�� !�3�E�W��{��_�� ��ÏՏ���`��/� �S�:�w���p����� џ������+��O� a���������ͯ߯ �D����9�K�]�o� �������ɿ���Կ �#�
�G�.�k�}�d� �ψ����Ͼ���n��� 1�C�U�g�yߋ��ϯ� ��4�����	��-�?� ��c�J������ ���������;�M�4� q�X����������� %7��[�� �����@� �3WiP�t �����/�// A/����w/�/�/�/�/ �/$/�/h?+?=?O? a?s?�?�/�?�?�?�? �?O�?'OOKO]ODO �OhO�O�O�O�ON/`/ _#_5_G_Y_k_�O�_ �_?�_�_�_�_oo �_Co*ogoyo`o�o�o �o�o�o�o�o-`Q8u�O�O}��@������)� >��U-�j�|������� ď+��Ϗ���B� )�f�M���������������ݟ�&�S�K��$UI_PANELINK 1�U�  ��  ��}1�234567890s���������ͯդ �Rq����!�3�E�W� �{�������ÿտm��m�&����Qo�  �0�B�T�f�x�� v�&ϲ���������� ��0�B�T�f�xߊ�"� �����������߲� >�P�b�t���0�� ����������$�L� ^�p�����,�>�����`�� $�0,&� [gI�m��� ����>P3 t�i��Ϻ�  -n��'/9/K/]/o/ �/t�/�/�/�/�/�/ ?�/)?;?M?_?q?�? �UQ�=�2"��?�? �?OO%O7O��OOaO sO�O�O�O�OJO�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5oGo�_ko}o�o�o �o�oTo�o�o1 C�ogy���� �B�	��-��Q� c�F�����|������ �֏�)��M���= �?��?/ȟڟ��� �"�?F�X�j�|��� ��/�į֯����� 0��?�?�?x������� ��ҿY����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z���� -���������
��. RdG��}� ���c���<�� `r������� �//&/8/J/�n/ �/�/�/�/�/7�I�[� 	�"?4?F?X?j?|?� �?�?�?�?�?�?�?O 0OBOTOfOxO�OO�O �O�O�O�O_�O,_>_ P_b_t_�__�_�_�_ �_�_oo�_:oLo^o po�o�o#o�o�o�o�o  ��6H�l~ a������� �2��V�h�K����� ��1�U
��.� @�R�d�W/�������� П������*�<�N� `�r��/�/?��̯ޯ ���&���J�\�n� ������3�ȿڿ��� �"ϱ�F�X�j�|ώ� �ϲ�A��������� 0߿�T�f�xߊߜ߮� =���������,�>� ��b�t�����+ ������:�L�/� p���e�����������  ��6���ۏ���$UI_QU�ICKMEN  }���}���RESTOR�E 1٩�  �
�8m3\n ���G���� /�4/F/X/j/|/' �/�/�//�/�/?? 0?�/T?f?x?�?�?�? Q?�?�?�?OO�/'O 9OKO�?�O�O�O�O�O qO�O__(_:_�O^_ p_�_�_�_QO[_�_�_ I_�_$o6oHoZoloo �o�o�o�o�o{o�o  2D�_Qcu�o �������.� @�R�d�v��������xЏ⏜SCRE� �?�u1�sc� u2�3��4�5�6�7��8��USER�����T���ksT'���4��5��6���7��8��� NDO_CFG ڱ�  �  � PD�ATE h���None�S�EUFRAME � ϖ��RTOL_ABRT�����ENB(��G�RP 1��	�?Cz  A�~�|��%|�������į֦��X�� UH�X�7�?MSK  K�S��7�N�%uT�%������VISCA�ND_MAXI��I�3���FAILO_IMGI�z �% �#S���IMREG�NUMI�
���S�IZI�� �ϔ�,�ONTMOU4'�K�Ε�&�����a��a���s�FR:\��� � M�C:\(�\LOGnh�B@Ԕ !{��Ϡ�����z �MCV����7UD1 �EX	��z ��PO64_t�Q��n6��PO!�LI�Oڞ�re�V�N�f@`��I�� =	_�SZ�Vmޘ��`�WA�Imߠ�STAT �k�% @��4�F��T�$#�x �2D�WP  ��P� G��=��������_JMP�ERR 1ޱ
�  �p2345678901��� 	�:�-�?�]�c����� ������������$�MLOW�ޘ�����g_TI/�˘'���MPHASE  �k�ԓ� ��SH�IFT%�1 Ǚ��<z��_� ���F/| Se������ �0///?/x/O/a/��/�/�/�/�/�����k�	VSFT1�\�	V��M+3 S�5�Ք p���ſA�  B8[0�[0�Πpg3a1Y2�_3Y�7ME��K�͗q	6e���&%���M���b��	���$��TDINEND3�4��4OH�+�G�1�OS2OIV I�{��]LRELEv�I��4.�@��1_AC�TIV�IT��B��A �m��/_��B�RDBГOZ�YBO�X �ǝf_\���b�2�TI�190.0.�P8�3p\�V254tp^�Ԓ	 �S��_�[b��r�obot84q_   p�9o\�pc�PZoMh�]�Hm�_Jk@1�o�ZA+BCd��k�,���P \�Xo}�o0); M�q����� ���>��aZ�b��_V