��   ��A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���D�RYRUN_T   � $'�ENB  $�NUM_PORT�A ESU@$STATE P _TCOL_��PM�PMCmGRP_�MASKZE� O�TIONNLOG�_INFONiA�VcFLTR_E�MPTYd $P�ROD__ L � P�C&J_  �4 $TYPE�NFST_IDX؞�_ICI � �MIX_BG�-�� G_NA�Mc %$MOD�c_USdCIFoY_TI< #�MKR-  �$LINc  { x_SIZa�#� .  �$USE_FL�GA�l�i�S�IMA�Q�QB��SCANRAX��IN�I��_C7OUNrRO�_�!_TMR_VA�gyh>� i�p'` ���H��!^%�$$CLA�SS  �����!��5��5� VIRTUR �/� '|/ �%5���U����8� ��!2�%I1�+ �M?_?q?�?�?�?�? �?�?�?OO%O7OIO`[OmO��+6W?�%{�! ��X�O�O�O  10�� ' 1�+G 4%zO*_��1 1_]_<_�_�_r_�_ �_�_�_�_�_#ooo Yo8oJo�ono1�C���-54�� �b1�d,1�!�a�o .@Rdv�� �����?~c�a 1&�8�J�\�n����� ����ȏڏ�����!��C�1�) U�g�y����� ����ӟ���	��-� �G�`�r��������� ̯ޯ���&�8�C� \�n���������ȿڿ ����"�4�F�Q�j� |ώϠϲ��������� ��0�B�M�_�xߊ� �߮����������� ,�>�P�[�t���� ����������(�:� L�^�i���������� ���� $6HZ e�w������� � 2DVh�F