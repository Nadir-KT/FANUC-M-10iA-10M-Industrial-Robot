��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 � �1�FP�CUREQ1 �� $SOFT�; T_ID�TO�TAL_EQ� �$� � NO�PS�_SPI_IND�E��$�X�S�CREEN_NA�ME �SIGN��� �PK_FIL	�$THKYMPA�NE�  	$_DUMMY � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"%�ASB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za4 q;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6�_�7_�8_�94:\qO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"YtP_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0�1p�3`?��D� �� Ќ@��hPV��mEX�p� �0g0�ۤ�p�r
$TF��2C$MD3i�T�O�3�0U� F� K��Hw2tC1(�	Ez�g0#E{"F�"F�40CP@�a2 m�@$�PPU�3N)ύRև�AX�!DU��AI�3BUF�F=�@�1 |pp���pP�IT� PP�M��M�y��F�SIMQSI�"ܢVA�ڤT��=�w T��`(zM��P�B�qF�ACTb�@EW��P1�BTv?�MC�� �$*1JqB`p�*1DEC���F���=�� ��H0CHNS_E;MP1�$G��8�B�@_4�3�p|@P��3�TCc�(r/�0-s x��ܐ� MBi��!����JR� i�SEGKFR��Iv �aR��TpN�C��PVF��?�bx & ��f{uJc!�Ja��� �!28�ץ�AJ���SI!Z�3S�c�B�TM����g��JaRSINF ȑb���q�۽�н脄���L�3�B���C3RC�e�3CCp�� ���c��mcҞb�1J��cѿ�.����D$ICb�Cq�5r�ե��@v�L'���EV���zF��_��F,pN��ܫ��?�4�0A�! �r���h�Ϩ��p �2�͕a�� �د��}R�Dx Ϗ ��o"27�!ARV�O`�C�$LG�pV�B@�1�P��@�t�aA�0�'�|�+0Ro�� M�Ep`"1 CRA 3 AZV�g6p��O �FCCb�`�`F��`K������ADI ��a�A�bA'�.p ��p�`�c�`S4PƑL�a�AMP��-`Y�3�P�M�]pUR��QU�A1  $@TITO1/S@S�!����"0�DBPXWO��zB0!5�$SK��L�2�DBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z���LB�)$�/���� %�/��$C�!&?�$ENE�q.'*?�Ú �RE�p2(H ���O�0#$L|3$$�#�B[�;�К�FO_D��ROSr�#������3�RIGGER�6P�ApS����ETUR�N�2�cMR_8�T�Uw��0EWM��M�GN�P���B#LAH�<E���P��O&$P� �'P@D�Q3�CkD{��DQฑ�4�11��FGO_oAWAY�BMO��t�Q#!� CS_�o)  �PIS�  I gb {s�C��A��[ �B$�S��AbP�@�EW-�TNTVճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_S}V�bEXCLU�:�nONL2��S1Y�*a&�OT�a'�HI_V�4��B���_ *P0� 9�y_z��p n�T;SG�� +nrr� @6Acc*b��G�#@E��V.iHb?fANNU�N$0.$fdID�U�2�SC@�`�i�a���j�fp�z��@I$2,�O�$FibW$}�O�T9@�1 $DUMMYk��da��d�n�� � �E- ` ͑HE4(sg��*b�SAB��SUFFmIW��@CA=��c5�g6r�!M�SW�E. 8Q�KgEYI5���TM�100s�qA�vIN���Ѹ�!��/ D��H7OST_P!�rk���ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  �8	=ȳ�r�DT�k0�!1 � $|S��ESAMPL��@j�۰f璱f���I�0|��[ $SUB��k�#0�C��T�r#a�SAVʅ��c���CX��P�fP$n0E��w YN_B#2 M0Q�DI{dlpO(���9#$�R_I��� �ENC2s_S� 3  5�C߰�f�- �SpU����!4�"g�޲�19T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9�g�DSP�v��PC���r"��(���ƓV7ALUߗHE�ԕ�M+�IPճ��OP5P ��TH��֤D��P�S� �۰F��df�J� ���C1�+6 H�bLL_DUs�~a3@{��3:���OTX"����s�r�0NOAUT5O�!7�p$)�$�*��c4�(�C�pR8�C, �""�L�� 8H *8�LH <6����c"�` , `Ĭ�kª�q��q���sq��~q��7��8J��9��0����1��U1̺1ٺ1�1�U1 �1�1�2(ʩ2����2̺2ٺ2��2�2 �2�2*�3(�3��3��̺U3ٺ3�3�3 ��3�3�4(%����?��!9 < �9�&�z��I��1���M��QFE@'@� �: ,6��Q? �@P?9��5�9�E�@A��a�A�z� ;p$TP�?$VARI:�Z�n��UP2�P< ���TDe���K`Q�p����q��BAC�"G= T�p��e$)_,p�bn�kp+ IFIG� kp�H  ��P����@`�!>t ;hE��sC�ST� D� D���c�<� 	C��{��_���l����R  ���FOR�CEUP?b��FL+US�`H�N>�F ����RD_CM�@E ������ ��@vMP��REMr F�Q��1������7Q
K4	NJ�5EFFۓ:�@3IN2Q��OVO��OVA�	TROV̷��DTՀ�DTMX� ��@�
ے�_PH"p��CL���_TpE�@�pK	_�(�Y_T��v(�J�@A;QD� �������!0tܑ0RQD���_�a����M��7�CL�dρRIV�'�{��EARۑI�OHPC�@����B��B��CM9@���R =�GCLF�e!�DYk(M�ap#5TuDG��� �%���FSSD �s? PP�a�!�1���P_�!��(�!1��E�3�!3z�+5�&�GRA��J7�@��;�PW���ONn��EBUG�_SD2H�P{�_E� A L��� �TERM`5B>i7 �ORI#e0�Ci5$Z �SM�_�P��e0D�9TA��9Ei6�PUP\�F�� -�A{�A�dPw3S@B$SEG��:� EL{UUSE.�@NFIJ�B$��;1젎4�4C$UFlP=�$,�|QR@"��_G90Tk�D��~SNST�PATx����APTHJ��E�p%B`�'EC���AR$P�I�aSHFTy�A�A�H_SHORР꣦6% �0$�7PE��E�GOVR=��aPI�@��U�b �QAYLOW���IE"�r�A8��?���ERV��XQ �Y��mG>@�BN��U���R2!P.uA�SYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC����EP;�uP;�6WOR�>@M`�0SM5T6�G3�GR��13�aPAL@���`�q�u_H � ���'TOCA�`P	P�`$OP����pѡ�`0O��R%E�`R4C�AO�p��Be�`R�Eu�h|�A��e$PWR�3IMu�RR_�cN�\�q=B I&2H���p_ADDR��H_LENG�B�q�qT�q$�R��S�JڢSS��SKN��u��0�u̳�uٳSE�A��jrS��MN�!K������b����O�LX��p����`ACRO3pJ�@��X��+��Q��6�OUP3�b_�IX��a�a1��}򚃳���(�� H��D��ٰ��氋�VIO2S�D������	�7�L $xd��`Y!_OFFr��PRM_��j^�aTTP_+�H:�wM (|pOBJ]"l�p��$��LE~C�d���N � \��֑AB_�Tq�b��S�`H�LVh��KR"uHITC�OU��BG�LO�q���h�����`���`SS� ���HQW�#A:�Oڠ<`�INCPU2VISIOW�͑��n��t�o��to�ٲ �IO�LN��P 8��R���p$SLob� PUT_n�$�p��P& ¢��Y F�_AS�"Q��$AL������Q  U�0�	P4A��^���ZPH�Y��-��x��UOI �#R `�K���@�$�u�"pP�pk���$�����&���UJ5�S-���NE�6WJOGKG̲DI�S���Kp���#T� (�uAVF�+`�C�TR�C
�FLAG�2�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w�  m�_�{0a�^��cg��� 4�����Ǝ���{0��� SCH_���a7��N�d�VW���E �"����4��UM�A�r�`LJ�@�DAUfՃEAU�p��d|�r�GqH�ba���BOO��WL ?�6 I�T��y0�REC���SCR ܓ�Dx
�\���MARGm� !��զ ��d%�����	S����W���U� ��JGM[�MNCH|J���FNKEY\��K��PRG��UF���7P��FWD��H]L��STP��V��=@��А�RS��HO`����C9T��b ��7�[�UL���6�(R�D� ����Gt��@P�O��������MD�F�OCU��RGEX.��TUI��I��4�@�L�����P����`��P��NE��CANA��Bj�oVAILI�CL !~�UDCS_HII4���s�O�(!�SH���S��ܜ�__BUFF�!X�5?PTH$m����v`�ěԃ�AtrY��?P��j�3��`O+S1Z2Z3Z�|�� Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�AC���K�&&z�� [ LQ��+0 0�	P���`#qdt
�U��dw<���_ \ ?�4Г�\��Ѩ#\0�C4�] ��CL�DPL��UTRQL�I��dڰ�)�$FLAG&�� 1�#�D����'B�LD�%�$�%ORGڰ5�2�PVŇV�Y8�s�T�r�$}d^ A���$6��$�%S�`�T� �B0�4�6RCLMC�4]?o?�9>���MI�p}dg_ d=њRQ�=�DSTB�p�c ;F�HHAX�R� JHdLEXCE�SrD�BM!p�a`���/B�Ta�B��`a�p=F_A7Ji��K�bOtH� K�db \�Q���v$MBC�L�I|�)SREQUI�R�R�a.\o�AXDESBUZ��ALt M���c�b�{P����2F�ANDRѧ`�`d;Ҙ2�ȺSDC��N�I�Nl�K�x`��X� N�&��aZ���UPS�T� ezrLO�C�RIrp�EX�<fA�p�9A�AOD�AQ��f XY�OND�rMF,Łf��s"��}%�e/� � w�FX3@IGG�� g ��t"���ܓs#N�s$R�a% ��iL��hL�v�@�ODATA#?pE��%�tR��Y�Nh �t $MD`qI�}�)nv� ytq�ytH�P`�Pxu��(�zsAN�SW)�yt@��yuD+�)AI^`���0o��i �@CUw�V��p 0XeRR2��j� Du�{Q��7Bd$OCALIA@��G�:�2��RIN��"��<E�NTE��Ck��r^�آXb]���_N�qlk���9�*����B�m��DIV��DH�@���qnI$V�,��S�$��$AZ�X�o�*�����oH �$B�ELT�u!ACC�EL�.�~�=�ICRC�� ���D�T��8�$PS�@�"L�@�r��#^�S�E�<� T�PATH3���DI���3x�p�A_W ��ڐ���2nC��4��_MG�$DDx��T���$FW��Rp9��I�4��DE�7�PPABN��R?OTSPEE�[g�� J��[�C@4�~�@$USE_+�2VPi��SYY��Z�1 qYN!@A��ǦOFF�qǡMO�U��NG���OL����INC�tMa6���HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]��BƉ�VE��#�y�23�_UP񕋳LOWL���p� B���Du�9B#P`�x ���ByCv�r�MOSI���BMOU��@�7PE�RCH  ȳOV ��â
ǝ����D �ScF�@MP����� !Vݡ�@y�j�LUk��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A��x������N`�F�RTI�A$��MOUЖ�HB@�BS0�p7D5����x��Z�DUM2ԓ�S_BCKLSH_Cx�k����ϣ����=���ޡ �	ACLAL"q��1м@N��CHK� �S�RTY��^�%E1rQq_�޴_UM�@r�C#��SCL0��r�LMT_J1_�L��9@H�qU�E�O�p�b�_�e�k�e�S�PC��u���N�P	C�N�Hz \P��C�0~"XT��C�N_:�N9��I�S	F!�?�V���U�/����x�T���CB!�SH�:��E�E1T�T�����y���T��PAL ��_P��_� �=������!����Jb6 L�@��OG��G�TORQU��ONֹ��E�R��H�E�&g_W2���_郅P���I�I�%I��Ff`xJ�1�,~1�VC3�0BD�B��1�@SBJ�RKF9�0DBOL_SM��2M�P�_DL2GRV�����fH_p��d���COS���LNH�� ������!*,�baZ���fMY��_(�TH��)TH�ET0��NK23����"��CB�&CB�CAA�B�"��!��!�&SB� 2�%'GTS�Ar�CIMa������,4#97#$DU���H\1� ���Bk62��AQ(rSf$NE�D�`I��B$+5��$̀�!A�%�5p�7���LPH�E�2���2SC%C�%�2-&FC0JM&̀V��8V�8߀LVJV�!KV/KV=KVKKV
YKVgIH�8FRM���#X!KH/KH=KH�KKHYKHgIO�<OR�8O�YNOJO!KUO/KO=KOKKOYKOM&F�2�!+i%0d��7SPBALANgCE_o![cLE0H_�%SPc� &�b�&�b&PFULC��h�b�g�b%p�1k�%�UTO_��Tg1T2�i/�2N�� "�{�t#�Ѱ`�0�*�.�T��OÀ<�v �INSEG"�ͱR�EV4vͰl�DIF��ŕ�1lzw��1m���OBpq�я?�M�I{���nLCHW3ARY�_�AB��!�?$MECH�!o X��q�AX��P��p��7Ђ�`n 
��d(�U�ROB��C�Rr�H���%��MSK_f`�p WP �`_��R/�k�z�����1S�~�|�`z�{���z��qINUq��MTCOM_�C� �q  ����pO�$NOR�En����pЂr� 8p GRe�uS�DZ�AB�$XYZ_DA�1a���DEBUUq�������s z`$��COD��� L���p��$BUFIN�DX|�  <�M{ORm�t $فUA��֐���r��<��rG��u � $SIMUL  �S�*�Y�̑a�OBJ�E�`̖ADJUS<�ݐAY_IS��D�3����_FI�=��Tu 7�~� 6�'��p} =�C�}p�@:b�D��FRIr��MT��RO@ \�E}z��y�OPWOY�q�v0Y�SYS�BU/@v�$SOP�ġd���ϪUΫ}pPgRUN����PA���D���rɡL�_OUbo顢q�$)�/IMAG��w��0�P_qIM��L�IN�v�K�RGOVR!Dt��X�(�P*�J�|��0L_�`]��0�RB1�����ML��ED}��p ��%N�PMֲ��oc�w��SL�`q�w x �$OVSL4vS;DI��DEX�� ��#���-�V} *�N4�\#�B�2�G�B�_�M�cy�q�>E� x Hw��p^��ATUSW����C�0o�s���BTMT�ǌ�I�k�4��x�԰q�y Dw�E&���@E�r��7�8�жЗ�EXE�����������f q�z �@w���UP'��$�pQ�XN�����x����� �PG΅�{ h $SUB����0_���!�_MPWAIv�P7�&��LOR���F\p˕�$RCVFAI�L_C���BWD�΁�v�DEFSP>!p | Lw����Я�\���UNI+�����H�R�+�}_L\pP��x�t���p�}H�> �*�j�(�ts`~�N�`KETB�J%�J�PE Ѓ~��=J0SIZE����hX�'���S�OR��?FORMAT�`�Ӱc ��WrEM�t���%�UX��G��P�LI��p�  �$ˀP_SWI��pq�J_PL��A�L_ �����AR��B��� C��D��$E��.�C�_�U�� � �� ���*�J3xK0����TIA4��u5��6��MOM��@������ˀB�ЃAD����������PU� NR�������m��� A$PI�6q��	� ����K4�)6��U��w`��SPEEDgPG������� �Ի�4T�� � 8@��SAMr`��p\�]��MOV_� _$�npt5��5���	1���2��������Ȣ'�S�Hp�IN �'�@�+�����4($4+T+GAMM�Wf�1'�$GETH`�p���Da���

pOLIBR>�II2�$HI=�_g�t��2�&E;��(A�.� �&LW�-6<�)56�&�]��v�p��V��?$PDCK���q"��_?�����q� &���7��4���9+�� �$IM_SR�pD�s�rF��r&�rLE���Om0H�]��0�-�pq���PJqUR_SC�RN�FA���S_SAVE_D��dE@�NOa�CAA�b�d@ �$q�Z�Iǡs	�I�  �J�K� ����H�L� �>�"hq����� �ɢ�� bW^UST�A��-M4��� a��)q`��3�WW�I@�v�_�=���MUAo�� � $PY+�θ�$W�P�vNG �{��P:��RA��RH��RO�PL�����q� (��s'�X;�OI�&��Zxe ���m�� p��ˀ�3s�O�O�O��O�O�aa�_т� |��q�d@��.v��.v@��d@��[wFv��E��P�%E�s;B�w�|�tP���PMA�Q]Ua ��Q8�ܾ1�QTH�HO�LG�QHYS��ES��qUE�pZB��]Oτ�  ��Pܐ@(�A����v�!�t�	O`�q��u�"���FA��IROG�����Q2���o�"��p��/INFOҁ�׃V�����R���OI���{ (�0SLEQ� �����Y�3����Á���P0Ow0����!E0NU��A�UT�A�COPY��=�/�'��@Mg�N@��=�}1������ ���RG��Á���X_�P�$;ख�`��W��P��@��������EXT_CYCB bHᝡRpÁ�r�n�_NAe!А����ROv`	��� � ���PO�R_�1�E2�SRV� �)_�I�DI��T_�k�}�'���dЇ�T����5��6��7��I8i�H�SdB���2�K$��F�p��GPqLeAdA
�TAR��@�@���P����裔d� ,�0FL�`�o@YN��K�Mz��Ck��PWR+��9ᘐ��DELA�}�dY�pAD�a}�#�QSKIP4�� �A�$�OB`NeT�} ��P_$� M�ƷF@\bIpݷ�ݷ �ݷd����빸��@Š�Ҡ�ߠ�9���J2R� ��� m4V�EX� TQQ� ����TQ������ ���`���RDC�V� )�`��X)�R�p������r��m$RGE7AR_� IOBT�2�FLG��fipER��DTC���Ԍ���2�TH2NS}� S1���G T\0' ���u�M\Ѫ`qI�d��REF��1Á� l�h��E�NAB��cTPE �04�]����Y�]��� �Qn#��*��"�����
��2�Қ�߼�����(����3�қ'�9�0K�]�o�� ����4�Ҝ������������5�ҝ!�3�E�PW�i�{��6�Ҟ��@�����������7���-?Qcu�8�Ҡ��������SMSKÁ��l��a��EkAޚ�MOTE6������@�݂TQ�IIO}5�IS�tR�9W@��� �pJ� ���p����E�"�$DSB_SIG!N�1UQ�x�C\��/S232���R�i�DEVICEUS��XRSRPARIT|��4!OPBIT�Q�I�OWCONT�R+�TQ��?SRCU�� MpSUXTAS�K�3N�p�0p$TATU�PE#�0������p_XPC)��$FREEFRO�MS	pna�GET\�0��UPD�A�2�aF"P� :���� !$USA�N�na&����ERI��0�RpRYq5*"_�j@�Pm1�!�6WR	K9KD���6��Q?FRIEND�Q�R�UFg�҃�0TOO�L�6MY�t$L�ENGTH_VT\�FIR�pC�@ˀyE> +IUFIN-R:M��RGI�1ÐOAITI�$GXñl3IvFG2v7G1�0��p3�B�GPR�p�1�F�O_n 0��!R�E��p�53҅U�TCp��3A�A�F �G(��":���e1n!� �J�8�%���%]��%�|� 74�X O0*�L��T�3H&��8P���%b453GE�W�0�WsR�TD����T���M����Q�T]�$V 2����1��R�91�8�02�;2k3�;3�:ifa�9-i��aQ��NS��ZR$V��2BVwEV�	V�B
;�����&�S�`���F�"�k�@�2a�PS�E��$r1C���_$Aܠ6wPR��7vMU�cS�t '�/89�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx������BSOC����N��DUMMY�14�p�0SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW_C�� �S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}����_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�S�A�pC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EG� �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G + AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC � o�ER|f�5� � $�@�_ A��!�PO���à�0#�
�_M�RAt�� d r� T��p�ERR��L=�;TY&���I��qV�0�cz�TOQ�d�PL[ �d�"�� ?�|w�! � pp`qT)0���_V1VrP�aӔ����2ٛ2薈E����@�H�E����$W�����V!��$�P��o�cI���aΣ	 HELL�_CFG!�� 5��B_BAS�q�SR3��� Ea#Sb���1�U%��2��3��4��U5��6��7��8����RO����I0�0NL�\CAB+�����ACK4�����,��p2@�&�?�_PUﳳCO. W�OUG�P�~ ����m�������T=Pհ_KAR�[@&_�RE*��P���|�QUE���uP�����CSTOPI_AL7�l�k0��h��]�l0SEM�4�(��M4�6�TYN�SO���DIZ�~�A������m_TM�MA'NRQ��k0E�����$KEYSWI�TCH���m���H=E��BEAT��|�E- LE~�����U±�F!Ĳ���B�O_�HOM=OGREFUPPR&��y!� �[�C��O��-EC�OC��Ԯ0_IOC1MWD
�a���m��� � Dh1���	UX���M�βgPgC�FORC��� �]��OM.  �� @�5(�U�#P�, 1��, 3��4�5���NPX_A�St�� 0��AD�D���$SIZ>��$VAR����TIP/�.��A�ҹM�ǐ��/�1�+ �U"S�U!Cz���F'RIF��J�S���5Ԓ�NF�� �� �� xp`SI��TqE�C���CSGL��	TQ2�@&����� ���STMT��,�P� �&BWuP��SHsOW4���SV��$�� �Q�A00�@Ma}���� ������&���5��6���7��8��9��A ��O ���Ѕ�Ӂ��� ��F��� G��0G ���0G���@G��PTG��1	1	1	U1+	18	1E	2��U2��2��2��2��U2��2��2��2��U2��2	2	2	U2+	28	2E	3��U3��3��3��3��U3��3��3��3��U3��3	3	3	U3+	38	3E	4�U4��4��4��4��U4��4��4��4��U4��4	4	4	U4+	48	4E	5�U5��5��5��5��U5��5��5��5��U5��5	5	5	U5+	58	5E	6�U6��6��6��6��U6��6��6��6��U6��6	6	6	U6+	68	6E	7�U7��7��7��7��U7��7��7��7��U7��7	7	7	�7+	78	7E��V�P��UPDs� � �`NЦ�
��SYSLOt�� � L��d���A�aTA�0d��|��ALU:ed�~�CU�ѰjgF!aID_L��ÑeHI�jI��$FILE_���d��c$2�
�cSA>�� hO��`E_B�LCK��b$��hD_CPUyM�yA���c�o�d�b����R ;�Đ
PW��!�[ oqLA��S=�8ts�q~tRUN�q st�q~t���qst�q�~t �T��ACC�s��X -$�qLEN;��tH��p�h�_�I��ǀLOWo_AXI�F1�q
�d2*�MZ���ă���W�Im�ւ�aR�TOR��pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v�������TCV��؁��T��ي�����t�V�H���V�Jj�R�MA�"��J��m�u�b����q2S�#�U�{�t�6K�JK��VK;���4H���3��J0�����JJ��JJ��AAAL��ڐ��ڐԖ4Օ5���N1���ʋ�ƀW�LP�_(�g�x,��pr�� `�`�GROUw`��B>��NFLIC��f�REQUIRE3�EBU��qB���w�2����p���q5�p��� \��APP�R��C}�Y�
ްE�N٨CLO7��SC_M��H���u�
�q�u�� �`�MCp�����9�_MG��C�Co��`M�в�N�wBRKL�NOL|�tN�[�R��_LIN�H��|�=�J����Pܔ ������������������6ɵ�̲8k�|D����� ���
��q)��7�PATH3�L�B�L��Hôwࡠ�J�CN�CaA�Ғ�ڢB�IN�r�UCV�4a��C!�U�M��Y,���aE��p����ʴ���PA�YLOA��J2L�`R_AN�q�L�pp���$�M�R_?F2LSHR��N�LOԡ�Rׯ�`ׯ�ACRL_G�Œ�ț� ��Hj`߂$yHM���FLEXܣ��qJ�u� :���������0����1�F1�V� j�@�R�d�v�������E����ȏڏ���� "�4�q���6�M���~�@��U�g�y�ယT��o�X��H������藕 ?�����ǟِݕ��ԕ����%�7�%|��J�� � V�0h�z���`AT�採6@�EL�� S���J|�Ŝ�JEy�C�TR��~�TN��F�Q��HAND_V�B-���v`�� $��F2M����eb�SW�b�'���O $$MF�:�Rg��(x�,4�%��0&A@�`�=��aM)F�AW�Z`i�Aw�A��X X�T'pi�Dw�D��Pf�G�p�)STk��!x��!N��DY�pנM� 9$`%Ц�H��H�c�@׎���0� ��Pѵ�ڵ��������9 ���� ����1��R�6��QASYIMvř���v��J�8��cі�_SH>��� �Ĥ�ED����������J�İ%��C�ID�.��_VI�!X�>2PV_UNIX�FThP�J��_R�5_Rc� cTz�pT�V��@���İ��߷��U ����Xd���Hqpˢ��faEN�3�DI�����O4d��`J�S� x g"IJAA�a z�aabp�coc�`a�p�dq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a�i�T�@<� $D�UMMY9Q�$7PS_��RFC��;$v �p���Pa� XƠ����STE���SBR�Y�M21_VF�8�$SV_ERF�O���LsdsCLRJtA���Odb`O�p �� D $GgLOBj�_LO����u�q�cAp�r�@aS;YS�qADR``�`TCH  �� ,��ɩb�W_N�A���7����TSR���l ���
*?�&Q� 0"?�;'?�I)?�Y)�� X���h���x������) ��Ռ�Ӷ�;��Ív��?��O�O�O�D�XS�CRE栘p��f��ST��s}y`L���Y�/_H�A�q� TơgpTYP�b���G�a�G���Od0ISb_䓀dEaUEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI@m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1 �ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���>EaVSHIF��Nc�P�`ג�E�ȐyR����OSUR��=Wk`RADILѮ��_�a��:�9a��`a��r��LULQ$O�UTPUT_BM����IM�AB �@��rTILSC	O��C7��� ����&��3��A����q���m�I�2"G�o�y@Md�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM�,�F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? ��ZABC%��  $�"R���
ϐ�$$CLA}S������!�p� � � VIRT8]��/ 0ABS�����1 5�� <  �!F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o �$6HZi{0-�A�XL�p��"�63  �{tIN��qztGPRE�����v�p��uLARMRECOV 9�rwt�NG�� .;	 A   �.�0�PPLIC��?�5�p�H�andlingT�ool o� 
�V7.50P/2�3-�  �Pfv��
��_SWt�w UP�!� x�#F0��t���A� v� 864��� �it�y� r�2 7wDA5�� �� ?Qf@��o��Noneisͅ�˰ ��T��~�!LAex>�E_l�V�uT��s9�UTO�"�Њt�y��?HGAPON
0g��1��Uh�D 1581����̟�ޟry����Q 1���p�,�蘦����;�@��q_��"{�" �c��.�H���D�HTTHK� Z��*� H�N���Ưد����  �2���V�h�z����� ��¿Կ���
��.� ��R�d�vϔϚϬϾ� ��������*߄�N� `�rߐߖߨߺ����� ����&��J�\�n� ������������� �"�|�F�X�j����� ������������ xBTf���� ����t> Pb������ ��//p/:/L/^/ |/�/�/�/�/�/�/�/  ??l?6?H?Z?x?~? �?�?�?�?�?�?�?OhO2O��TO�E�W��DO_CLEAN���7��CNM  � �__/_�A_S_�DSPDR3YR�O��HIc��M@�O�_�_�_�_oo +o=oOoaoso�o�o���pB��v �u���a�X�t������9�PL�UGG���G��U�P�RCvPB�@���_�orOr_7�SEGF}�K[mwxq �O�O�����?rqLAP�_�~q�[� m��������Ǐُ�����!�3�x�TOT�AL�f yx�USE+NU�p�� �H����B��RG_STR�ING 1u�
_�Mn�S5��
ȑ_ITEM1Җ  n5�� � �$�6�H�Z�l�~��� ����Ưد���� ��2�D�I/O �SIGNAL̕�Tryout �ModeӕIn�p��Simula�tedבOut���OVERR~�P = 100֒�In cycl���בProg OAbor��ב���StatusՓ	�Heartbea�tїMH Fa�ul��Aler '�W�E�W�i�{ύϟ�p�������� �C Λ�A����8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|���WOR{pΛ��(ߎ� ���� ��$�6�H�Z� l�~�������������p�� 2PƠ �X ��A{��� ����/A Sew�����SDEV[�o� #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1?�C?U?g?y?PALTݠ1��z?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_�?GRI�`ΛDQ�? _l_~_�_�_�_�_�_ �_�_o o2oDoVoho@zo�o�o�o2_l�R� �a\_�o"4FX j|����������0�B�T��oPREG�>�� f��� Ə؏���� �2�D� V�h�z�������ԟ����Z��$ARG�_��D ?	����;��  	$Z�W	[O�]O��Z��p�.�SBN_CONFIG ;�ꎱ����CII�_SAVE  �Z�����.�TCE�LLSETUP �;�%HOM�E_IOZ�Z�%�MOV_��
�R�EP�lU�(�UTOoBACKܠ���FRA:\�z� \�z�Ǡ'�`�z���ǡi�I�NI�0z���~n�MESSAG����ǡC���ODE_!D������%�O�4��n�PAUSX!�~;� ((O>� �ϞˈϾϬ������ ����*�`�N߄�r��߶�g�l TSK � wͥ�_�q�UP3DT+��d!�AſWSM_CF���;���'�-�GRgP 2:�?� N��BŰA��%�XSC�RD1�1
7� 	�ĥĢ�������� ��*�������r��� ��������7���[� &8J\n��*�>t�GROUN�UϾ�UP_NA��:�	t��_ED��17�
 �%�-BCKEDT�-�2�'K�`�ܵu�z�q�,q�z���2t1�����q�k�(/��ED3/��/��.a/�/;/M/ED4�/t/)?�/.?p?�/�/ED5`??�?�<?.�?O�?�?ED6O�?qO�?.MO�O'O9OED7�O`O_��O.�O\_�O�OEDa8L_,�_�^-p�_ oo_�_ED9�_�_]o�_	-9o�oo%oCR_ 9]��oF�o�k� � NO�_DEL��GE?_UNUSE���LAL_OUT �����WD_ABORﰨ~��pITR_RTN�=��|NONSk����˥CAM_PARAM 1;��!�
 8
SO�NY XC-56� 2345678�90 ਡ@����?��( �А\�
���{��:��^�HR5q�̹���ŏR57ڏ�A�ff��KOW�A SC310M�
�x�̆�d @<�
���e�^ ��П\����*�<���`�r�g�CE_R�IA_I�!��=�F��}�z� ]��_LIU�]�V����<��FB��GP 1���Ǯ�M�_�q�0�Cg*  ����C1���9��@��G���CVR�C]��d��l��Es��R�����[ԴUm��v�������_�� C����(������=�HE�`O�NFIǰ�B�G_�PRI 1�{ V���ߖϨϺ�����������CHKPA�US�� 1K� ,!uD�V�@�z�d� �߈ߚ��߾������.��R�<�b���OƯ�������_MkOR�� �^<:��� 	 ��� ��*��N�<����䡑��?��q?;�;�����K��9�P��|�ça�-:���	�

��M��@�pU�ð��<��,~���DB���튒)�
mc:cpmi�dbg�f�:�/  ��¥��p�/�  U���ȋ��� ��s>�  �ٕ�U�?U�苐�Ug�T/�W��XUf��M/w�O/�
DEF 3l��s)�< buf.txts/��t/��ާ�)�	�`�����=L�Ͷ�*MC��1�����?43��1���t�īCz  BH�H�CPUeB�$��BPI�7����C���C���Y
K�D�nyD���Cx�9�;�
D�� D���^�=Fr���E�CeE�� �=7Y�F��F�;�p4��*w�1����s���.��p����BDw�M@)x8��1Ҩ����g@5DPD�0EYK��EX�EQ��EJP F�E��F� G���>^F E�� �FB� H,- �Ge��H3Y���:�  >�33� ���~  in8�~@��5Y�E�>�ðA��Y<#�
"Q ���+_�'�RSMOFS�pؒ.8��)T1��DEg ��F 
Qv��;�(P  B_<_��R����	op6�C4P�Y
P]A(Q�2PC�0B3�Ma�C{@@*cw��UT��pFPROG !%�z�o�oigI�q����v��ldKEY_TOBL  �&S�#�� �	
��� !"#$%&'�()*+,-./�01i�:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�����������������������p`LCK�l4�p`�`STAT� ��S_AUTO_�DO���5�IN?DT_ENB!���1R�Q?�1�T2}�^��STOPb���TR�Lr`LETE���Ċ_SCREEN� �Zkc�sc��U��MME�NU 1 �Y  <�l�oR�Y 1�[���v�m���̟�� ���ٟ�8��!�G� ��W�i��������ï կ��4���j�A�S� ��w�����迿�ѿ� ���T�+�=�cϜ�s� ���ϩϻ������� P�'�9߆�]�o߼ߓ� ���������:��#� p�G�Y������� ����$����3�l�C� U���y������������ ��	VY)�_M�ANUA�0���$�DBCO[�RIG|ڇ
�DBNUM� Ҟ�B1 e
�PXWORK 1!�[�_U/4FX��_AWAY�^i�GCP  b=�Pj_AL� #�j��Y��܅ `�_�  �1"�[ , 
�od�&/~&l%MZ�IdPx@P@#�ONTIMه�& d�`&�
�e�MOTNEND�o��RECORD �1(�[g2�/{�O��!�/ky"?4? F?X?�(`?�?�/�?? �?�?�?�?�?)O�?MO �?qO�O�O�OBO�O:O �O^O_%_7_I_�Om_ �O�_ _�_�_�_�_Z_ o~_3o�_Woio{o�o �_�o o�oDo�o /�oS�oL�o�� ��@���+�y V,�c�u�������� Ϗ>�P�����;�&� ��q���򏧟��P�ȟ �^������I�[�� ��� ���$�6��������jTOLER7ENCwB����L�͖ CS_C�FG )�/'d�MC:\U�L�%04d.CSVd�� c��/#A ��+CH��z� //.�ɿ��(S�RC_O_UT *��~�SGN +���"��#�29-�JAN-20 2o3:09015l��10:51+ P/Vt�ɞ�/.���f�pa�m�?�PJPѲ���VERSION �Y�V2.�0.84,EFLO�GIC 1,� 	:ޠ=�ޠ�L��PROG_E�NB��"p�ULS�k' ����_WRSTJNK ��"f�EMO_OPT_�SL ?	�#
� 	R575 /#=�����0�B��>��TO  �ݵ�l���V_F EX��d�%��PATHw AY�A\�����5+ICT�F�u-�j�#�egS�,�ST?BF_TTS�(�	�d���l#!w�� M�AU��z�^"MSWX�.��4,#�Y�/�
!J�6%�ZI~m��$SB�L_FAUL(�0��9'TDIA[�1�<�� ����12345678#90
��P��H Zl~����� ��/ /2/D/V/h/��� P� ѩ �yƽ/��6�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�,/�gUMP���� ��ATR���1OC@P�MEl�OOY_TE{MP?�È�3F�8��G�|DUNI��.��YN_BRK �2_�/�EMGDI�_STA��]��EN�C2_SCR 3�K7(_:_L_^_ l&_�_�_�_�_)��C�A14_�/oo/o�AoԢ�B�T5�K�ϋo~ol�{_�o�o �o'9K]o �������� �#�5��/V�h�z��� �`~�����ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T���x������� ��ү�����,�>� P�b�t���������ο ����(�f�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ���������:�  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� �����*<N `r������ �&8J\n ���������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?��? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O��O�O__NoETM�ODE 16�5]�Q �d�X�
X_j_|Q�PRRO�R_PROG �%GZ%�@��_  ��UTABLE  G[�?oo)oRj�RRSEV_NU�M  �`WP��QQY`�Q_AU�TO_ENB  q�eOS�T_NOna� 7G[�QXb�  *��`��`��`��`d`+�`�o�o�o�dHISUc�QOP��k_ALM 18.G[ �A��l�P+�ok}������o_Nb�`  �G[�a�R
�:PTC�P_VER !�GZ!�_�$EXTLOG_REQvs�i\�SIZe�~W�TOL  �Q{Dzr�A W�_BWD�p��xf́�t�_DI�� 9�5�d�T�QsRֆSTEP��:P�_OP_DOv�f��PFACTORY�_TUNwdM�E�ATURE :��5̀rQH�andlingT�ool �� \s�fmEngl�ish Dict�ionary��r�oduAA �Vis�� Mas�ter����
E�N̐nalog �I/O����g.f�d̐uto So�ftware U�pdate  F� OR�mati�c Backup~��H596,��ground E�ditޒ  1 �H5Came�ra�F��OPL�GX�ell𜩐IwI) X�ommՐsshw���com��sco���\tp����pane��  �opl��tyle select��/al C��nJ�Ց�onitor��R�DE��tr��R�eliab𠧒6�U�Diagnosx(�푥�5528��u��heck S�afety UI�F��Enhanc�ed Rob S�erv%�q ) �"S�r�User �Fr[�����a��xt. DIO ��fiG� sŢ��e�ndx�Err�L&F� pȐĳr됮�� ����  !��F�CTN Menu�`�v-�ݡ���TPw Inېfac��  ER J�GC�pבk Ex�ct�g��H558���igh-Spe�x�Ski1�  2�
P��?���mm�unic'�ons��&�l�ur�ې���ST Ǡ��co�nn��2��TXP�L��ncr�st�ru����"FAT�KAREL �Cmd. LE�u�aG�545\��R�un-Ti��En=v��d
!����ؠ++�s)�S/W���[�LicegnseZ��� 4T��0�ogBook(�Syڐm)��H5�4O�MACROs�,\�/Offsen��Loa�MH��ܽ���r, k�Me�chStop P�rot���� li�c/�MiвShiqf����ɒMixx���)���xStS�M�ode Swit�ch�� R5W�M�o�:�.�� 74� ���g��K�2~h�ulti-T=��M���LN (�Pos�Regi�ڑ������d�ݐt 'Fun�ǩ�.�����Num~����� �lne��ᝰ A�djup����� � - W��tat�uw᧒T�R�DMz�ot��scWove U�9����3Ѓ�uest' 492�*�o������62;�SNPX� b ���8 J7<`���Libr��J�#48���ӗ� �Ԅ��
�6O�� Par�ts in VCCMt�32���	��{Ѥ�J990��/�I� 2 P��T_MILIB��H�:��P�AccD�L�o
TE$TX��n��ap1S�Te����pkey��w����d��Une�xceptx�mo�tnZ��������є�� O����� 90J�єSP CSXC<�f���6�� Py�We}���gPRI�>vrЮt�men�� ��iPɰa������vGrid�pl�ay��v��0�)�H�1�M-10iA�(B201 �2�\� 0\k/�Ascii�l�Т�ɐ�/�Col��ԑGu�ar� 
�� /Pl-�ޠ"K��st{�Pat ��!S�C�yc�҂�ori�e��IF8�ata- quҐ�� ƶ���mH574��RL���am���Pb�H_MI De3�(b�����PCϺ�Pa�sswo+!��"P�E? Sp$�[���t�p��� ven��T�w�N�p�YELL�OW BOE	k$A;rc��vis��y3*�n0WeldW��cial�7�V#t&�Op����1y�� 2F�a�por1tN�(�p�T1�T�0 �� ��xy]�&kTX��tw�igjx�1� b� ct\��JPN ARCPSU PR��oݲ�OL� Sup�2f�il� &PAɰאc{ro�� "PM(�X���O$SS� eв7tex�� r���z=�t�ssagT��P��P@�Ȱ�����rtW��H'>�r�dpn��n1�
t�!� z ��a�scbin4ps�yn��+Aj�M �HEL�NCL �VIS PKGS� PLOA`�MB� �,�4VW�R�IPE GET_�VAR FIE �3\t��FL[�O�OL: ADD �R729.FD �\j8'�CsQ�QE���DVvQ�sQNO? WTWTE��}PD  �^��biR�FOR ��ECT�n�`��ALSE �ALAfPCPMO�-130  M"� #h�D: HANG FROMmP��AQfr��R70�9 DRAM A�VAILCHEC�KSO!��sQVPC�S SU�@LIM�CHK Q +P~dF_F POS��F�Q� R5938�-12 CHAR�Y�0�PROGRAy W�SAVEN`wAME�P.SV��7��$En*��p?F�U�{�TRC|� S�HADV0UPDA�T KCJўRST�ATI�`�P MU�CH y�1��IM�Q MOTN-0�03��}�ROBO�GUIDE DA�UGH�a���*�t�ou����I� Šh�d�ATH�PepMO�VET�ǔVMX�PACK MAY ASSERT�Dn��YCLfqTA�r�BE COR v�r*Q3rAN�pRC� OPTIONS�J1vr̐PSH-�171Z@x�tcǠSU1�1Hp^9R!�Q��`_T�P��'�j��d{tby ap?p wa 5I�~d��PHI���p�aTE�L�MXSPD �TB5bLu 1��UBl6@�qENJ`CE2��61��p��s	�m�ay n�0� R�6{�R� �Rtrasff)�� 40*��p��fr��sys�var scr �J7��cj`DJUD��bH V��Q/�PSET ERR`�J` 68��PND�ANT SCRE�EN UNREAh��'�J`D�pPA��z�pR`IO 1����PFI�pB�pGROUN�PD��G��R��P�QnRSVIP �!p�a�PDIGIT� VERS�r}BL�o�UEWϕ P0�6  �!��MAG`p�abZV�DI<�`� SSUE�ܰ��EPLAN J=OT` DEL�pݡ�#Z�@D͐CAL9LOb�Q ph��RޫQIPND��IM�G�R719��MwNT/�PES �puVL�c��Hol�08Cq���tPG:�`C��M�canΠ��p�g.v�S: 3D� mK�view ed�` �p��ea7�:��b� of �Py����ANNOT ACCESS M��tƁ*�t4s a���lok��Flexj/:�Rw!mo?�PA?�-�����`n�pa SNBPJ? AUTO-�06f�����TB��PIAB{LE1q 636���PLN: RG$�pul;pNWFMDB��VI���tWIT �9x�0@o��Qui�#0�ҺPN RRS�?pUSB�� t & remov�@� )�_��&AxEPF�T_=� 7<`�pP�:�OS-144 ��h s�g��@�OST� � CR�ASH DU 9^��$P�pW� �.$��LOGIN���8&�J��6b04�6 issue �6 Jg��: Solow �st��?c (Hos`�c����`IL`IMPR�WtSPOT:Wh�:0�T�STYW ./�VMGR�h�T0wCAT��hos���E�q��� �O:�S:+pRTU' k�e-S� ����E:���pv@�2�� t\h�ߐ��m ��alļ�0�  $�H� W�A͐��3 CNT�0 T�� Wro>U�alarm���0s�d � �0SE1���t�r R{�OMEBp����K� 55��R�EàSEst��g �    �KA7NJI�no����INISITALcIZ-p�dn1weρl<��dr�� lx`~�SCII L�fails w��y ��`�YSTEa�p��o��Pv� IIH����1W�Gro>Pmo ol\wpSh@��P��Ϡn cfl�xL@АWRI �OGF Lq��p?�F��up��de-re�la�d "AP�o SY�ch�Abe�twe:0IND 1t0$gbDO����r� `�GigE��#operabi-lf  PAbHi�H`���c�lead�\�etf�Ps�r�O�S 030�&: fi=g��GLA )P ���i��7Np tpkswx�B��If�Ag������5aE�a EXCE#dU�_��tPCLOS��"r[ob�NTdpFa�U�c�!���PNI�O V750�Q1p��Qa��DB ��b�P M�+P�QED��DET��-� \r�k��ONLINEhSBUGIQ ߔĠ,i`Z�IB�S ap�ABC JARK�YFq� ���0MI�L�`� R�pNД \�p0GAR��D*pqR��P�"! jK�0cT�P�Hl#n�a��ZE V�� TA;SK�$VP2(�4`�
�!�$�P�`WIB�PK05�!FȐB�/��BUSY R7UNN�� "��d���R-p�LO��N�DIVY�CUL���fsfoaBW�p���30	V���ˠIT`�a50�5.�@OF�UN#EX�P1b�af�@�}E��SVEMG� �NMLq� D0pC?C_SAFEX 0c��08"qD �PETr�`N@�#J87��B��RsP�A'�M��K�`K�H GU�NCHG۔MEC�H�pMc� T�  �y, g@�$ OR?Y LEAKA�;�ޢSPEm�Ja��V�tGRIܱ�@އCTLN�TRpk�FpepR�j50�EN-`IN�����p� �`�Ǒk!��T3�/dqo�STO�0A�#�L�p �0�@�Q��АY�&�;pb1T!O8pP�s���FB�@�Yp`�`DU��aO��supk�t4 � P�F�� Bnf�Q�PSV�GN-1��V�SRSR)J�UP�a2�Q�#D�q l O���QBRKCTR 5Ұ�|"-�r�<pc��j!INVP�D ZO� ��T`h#�Q�cH�set,|D��"D�UAL� w�2*BRVO117 A]��TNѫt�+bTa24�73��q.?��sAU�z�i�B�compl�ete��604.�� -�`han�c�U� F��eN8��  ��npJtPpd!q��`��� 5h'596p�!5d�� @"p�P�P�Q�0�P2�p �A� xP��R(}\xP�e� aʰI���E���1��p� j  �� xS?t�^t �A��AxP�q 5 sig:��a��"AC;a���
�bCexPb_p���.pc]l<bHbc?b_circ~h<n�`tl1�~`xP`o�d�xP�b]o2�� �cb��c�ixP�jupfr�m�dxP�o�`exe��a�oFdxPtped�}o��u`�cptli1bxzxP�lcr�xrxP\�blsazEdxP_fm�}gcxP�x�� �o|sp�o�mc(��o'b_jzop�u6��wf��t��wms�1�q��sld�)��jm!c�o\�n��nuhЕ�ƭ|st�e��>�pl�qp�iwck���u�vf0uߒ��lvi�sn�Cgacul�wQ
E F  !� Fc.fd�Qv��� qw���Data� Acquisi��nF�|1�RR63�1`��TR�QDMCkM �2�P75H�]1�P583xP1��[71��59`�5�P57<PxP�Q����a(���Q��o pxP^!daq\�oA���@�� ge/�et�dms�"DMER9"؟,�pgdD����.�m���-��qaq1.<᡾xPmo��h����f{�u�`13��M�ACROs, Sksaff�@z����0E3�SR�Q(��Q6��E1�Q9ӡ�R�ZSh���PxPJ643�@7bؠ6�P�@�PRS�@����e �Q�UС P�IK�Q52 PT�LC�W��xP3 (��p/O��!�Pn� �xP5��03\�sfmnmc "MNMCq�<��Q��5\$AcX�FM��� ci,Ҥ�X����cdpql+�
�sk�SK�<xP�SH560,P���,�y�refp �"REFp�d�A�jlxP	�of�OFc�l<gy�to�TO_�x���ٺ���+j�e�u��caxis�2�xPE�\�e�q"I�SDTc��]�pr7ax ��MN��<u�b�isde܃h��\�w�xP! isb�asic��B� yP]��QAxes��R6������.�(B9a�Q�ess�� xP���2�D�@�z�atis���(�{������~��m��FM�c�u�{�
ѩ�MNIS��ݝ����x�����ٺ��x� j75���Devic�� �Interfacx�RȔQJ754��� xP�Ne`�� xP�ϐ2�б����{dn� "DNE�����
tpdnui�5UI��ݝ	bd��bP�q_rso�fOb
dv_aro��u�����stchkc��zp	 �(}onl��G!ffL+H�J( ��"l"/�n�b��<�z�hamp��T�eC�!i�a"�59�0�S�q��0 (�+P�`o�u�!2��xpc_2�pcchm��CH�MP_�|8бpev�ws��2쳌pcs|F��#C SenxPacro�U·�-�R6�Pd�xPk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GEM�,\i(��Dgesnd�5���H{�}Ha�@csy���c�Isu�xD��Fmd��I��7�4����u���AccuCal�P�4� ��ɢ�7ޠB0��6+6f�6��99\aFF q��S(�U��2�
X�p0�!Bd��cb_�Sa{UL��  �� �?�ܖto��otp�lus\tsrnPغ�qb�Wp��t����1��Tool (?N. A.)�[K�7�Z�(P�m���țbfcls� k9�4�"K4p��qtp{ap� "PS9|H�stpswo��0�p�L7��t\�q�� ��D�yt5�4�q��w��q��� �M�uk��rkey����s��}|t�sfeatu6�CEA��� cf)t\Xq`�����d�h5����LRC0�md�!�5!87���aR�(�����2V��8c?u3l\�pa3}H�&r-�Xuļ��t,�� �q " �q�Ot��~,���{�/ ��1c�}����y�p� r��5���S�XAg�-�xy���Wj874�- iRVis���Queu�� �@��-�6�1���(����u���tӑ�����
�tpvtsn "VTSN�3C�+�:� v\pRDV����^*�prdq\�Q�&�vstk=P�������nm&_�դ�c�lrqν���ge�t�TX��Bd���apoQϿ�0qstr�D[� ��t�p'Z�����npv��@�enl IP0��D!x�'�|���csc ߸��tvo/@��2�q���vb� ���q���!���h]����(� Cont�rol�PRAX:�P5��556�A@�59�P56.@56r@5A�J69$@�982 J552 IDVR7�hqA���16�H���La��� ��Xe�frlparm.f�7FRL�am��C9�@(F�����w6�{���A��QJ64�3�� 50�0LS�E
_pVAR $SGSYSC���RS_UNITS� �P�2�4tA�TX�.$VNUM_OLD 5�1�xP{�ƈ50+�"�` Funct���5tA� P}��`#@�`3�a0�c�ڂ��9���@H5 נ� �P���(�A�� ��۶}����ֻ�}��bPRb�߶~pp=r4�TPSPI�3�}�r�10�#;A� �t�
`���1���96�����%C�� Aفz��J�bIncr�	 ����\���1o5�qni4�MNIN�p	xP�`���!��H�our  �� 2�21 ~�AAVM��̳�0 ��TU�P ��J54s5 ��6162��VCAM  �(�CLIO= ��R6�N2��MSC "P� �STYL��C�28~ 13\��NRE "FH�RM SCH^��DCSU%OR�SR {b�04 ~�EIOC�1{ j 542 � �os| � egiCst�����7��1�MASK6�934"7 ��OOCO ��"3��8��2���� 0� HB��� 4�"39N� Re�� ��LCHK
%OPL�G%��3"%MHCMR.%MC  ; 4? ���6 dPI�5�4�s� DSW%M�D� pQ�K!637��0�0p"�1�Р"4� �6<27 CT�N K � 5 ����"7��<25�%/�T��%FRDM� �Sxg!��930 FB�( NBA�P� ( HLB  Men��SM$@jB( PVC� ��20v��2H�TC�CTM�IL��\@PAC c16U�hAJ`SAI N\@ELN��<29s�UECK �b��@FRM �b�O�R���IPL��R>k0CSXC ����VVFnaTg@HT�TP �!26 ���G�@obI�GUI"%IPGS|�r� H863 qbp�!�07r�!34 �r>�84 \so`!� Qx`CC3 Fb�21��!96 rb!531 ���!53R% E1!s3!��~�.p"�9js VATFUJG775"��pLR6^R�P�WSMjUCT�O�@xT58 F!890���1XY ta3!�770 ��88M5�UOL  GTSox
�{` LCM �r�| TSS�EfP6 |W�\@CPE `���0VR� l�QNL�"��@001 imrb�c3 =�b�0���0�`6 w�b-P�- R-�b8n@5EW�b9 �Ґa� ���b�`ׁ�b2 2'000��`3��`	4*5�`5!�c�#$��`7.%�`8 h6�05? U0�@B6iE"aRp7� !Pr�8 t�a@�tr2O iB/�1vp3�&vp5 Ȃtr9Σ�a�4@-p�r3 F��r5&�re`u��r�7 ��r8�U�p9? \h738�a�_R2D7"�1f���2&�7� �3 S7iC��4>w5Ip��Or60 C�L�1lbEN�4 I�pyL�`uP��@N�-PJ8�2N�8NeN�9 H�r`�E�b7]�|���q8�Вࠂ9 2���a`0�qЂ5�%U�097 0��@18�0���1 (�q�3 5R���0����mpU��0�0�7�*�H@(q�\P"R;B6�q124�b;�0�@���@06� x�3 pB/x�u ��~x�6 H606�a�1� ��7 6 ����p�b155� ����7jUU1632 �3 g���4*�65 2e 1"_��P�4U1`��ҢB1���`0'�17�4 �q��P�E18�6 R ��P�7 t��P�8&�3 (��90 B/�s1981����@202���6 3���A�RU�2� d��2 b2$h`��4�᪂2�4�&��19v Q�2��u�2d�Tpt2� ��H"�a2hP�$�5���!#U2�p�p
�2�p��B�@5�0-@��8 @�9��TX@�� �e�5�`rb26Af�2 ^R�a�2Kp��1y�bQ5Hp�`
�5�0@�0gqGA���a52ѐ��Z��6�60ہ5� Jׁ2��8�E��9�ESU5@ٰ\�q5hQT`S�2ޖ5�p\w�@۲�pJ �-P��5�p�1\t�H�4��PC2H�7j��phiw�@���P�x��559 ldu� P�D���Q�@������� �`.��Pt>��8�581�"6�q58�!AM۲T��A iC�a589`��@�x����5 �a��12׀0.�1����,�2����,�!P\hI8��Lp ��,�7���6�0840\� A?NRS 0C}A��0p��{��ran��FRA��Д�е� ��A%���ѹ�Ҍ� ����(����Ќ��� �З���������ь����$�G��1��ը����������� xS�`q�  X�����`64��M���iC/50T-H�������*��)p46���� C��N����mw75s֐� Sp��b46��v�����^�M-71?�7�������42������dC��-�а�70�r$�E��/h�����O$��rD���c7c7C�q��Ѕ���L��/��2\imm7c7�g������`���(�� e�����"������`�a r��c�T,����"��,�� ��x�<Ex�m77t����k���5�����)�;iC��-HS- � B
_�>���+����7U�]���Mh7�s��7�������-9?�/260L_������Qҡ������]�9pAA/@���q�S�������h6251��c��92���p����.�)92c0� g$�@�����)$��85$���pylH"O"�
�21���t?�350����p��`$�
�� �350!����0��9�U/0�\m9��M9A3���4%� s��3�M$��X%u���"him98J3����� i Ad�"m4~�103p�x� ����h794̂�&R���H�0����\� ���g�5AU��՜��0 ���*2��00��#06�АՃ�է!07{r ������� ��kЙ@����EP�#������?��8#!�;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?���CD25L�����0�"l�2BL 
#��B��\20�2_� r�re���X��1�� N����A@��z��`�C�pU��`��0�4��DyA�\�`f Q��sU���\�5�  ��� �p�^t��<$85����+P=�ab1l���1LT��lA8��!uDnE(�20T⧰J�1 e�bH85����b�Ռ�5[�16�Bs��������d2p��x��m6t! `Q����bˀ���b#�(�6iB;S�p�!� �3� ��b�s��-`�_�W8�_�����6I	$�X5�1�U815��R�p6S��� �/�/+q�!�q��`��6o��5m[o)�m6�sW��Q�?��se�t06p ��3%H�5��10p$����g/��JrH��  s��A�856�Ȝ��F�� ���p/2���h�܅�✐)�5���̑v��(��m	6��Y�H�ѝ̑m�Q6�Ҝ��a6�DM��F��-S�+��H2� ����Ҽ�� �r̑���✐��l���p�1���F���2�\t;6h T6H��� �Ҝ�'Vl���ᜐ��V7ᜐ/����;3A7��p~S��������4�`圐�V���*!3��2�PM[���%ܖO�chn��v�el5����Vq���_arp#��̑�.���?2l_hemq$�.�'�6415���5� ��?����F�����A5g�L�ј[���1��Ȝ�𙋹1����M7NU�М��eʾ�����uq$D;��-�4��3&H�f�c�Ĝ�h� ������u��� 㜐��ZS�!ܑ4���M-����S�$̑��� �� 0��<�����\07shJ�H�v �À�sF��S*󜐳� ��̑���vl�3�A�T�#��QȚ�Te��q�cpr����T@75j�5�dd�̑1�(UL�&� (�,���0�\�?���̑��a�� xStA���a�e�w�2��d(�	�2�C��A/����\�+p�����21s (ܱ�CL S�� ��B̺��7F���4?�<�lơ1L����c� ���u9�0����Ce/q��O���9�K��r9 (��,�Rs��ז�5�G�m2�0c��i��w�2 ��:�0`�$��2�2lҀ0�k�X�S� ,�ι2���O���1!41�w���2T@� _std��G�y� �ң�H� jdgm����w0 \� �1L���	�P�@~�W*�b��t 5��(����3�,���AE{������L��&�5\L��3�L�@|#~���~!���4�#@��O����h�L6A�������2璥����44�����[6\j4s��·���# ��ol�E"w�8Pk� ����?0xj�H1�1Rr��>��]�2a�2�Aw�P ��2��|41 �8��ˡ��{� �%�A<��� +�?�l��0�&0�"��|�`Am1�2� �ػ��3�HqB�� ��K�R��ˑb�W��� Fs���)�ѐ�!����a�1����5��16�16C��C����0\imBQ��d�P���b��\B5�-���DiL���O�_�<ѠPEtL�E�RH�Z�p�Pgω�am1l�� u���̑�b�<����<�$�T�̑�F���@�Ȋ�Dpb��X"�ἒ���p� ����^t��9�0\� j�971\kckrcfJ�F�s�����c���e "CTME��r�����!�a�`ma�in.[��g�`r#un}�_vc�#0 �w�1Oܕ_u����bctme��Ӧ�`ܑޅj735�- �KAREL UsKe {�U���J�P�1���p� Ȗ �9�B@��L�9��7�j[�atk208� "K��Kя��\��9��a��̹���N�cKRC�a�o ��kc�qJ�&s����� Grſ�fsD��:y��s���A1X\j|хrd�tB�, ��`.v�q�� �sǑIf�Wf�j52�TKQut_o Set��J�w H5K536(��932���91�58�(�9�BA�1(�74�O,A$�(TCP �Ak���/�)Y� ��\tpqtoo�l.v��v���!? conre;a#��Control �Re�ble��CNRE(�T�<�4�2����D�)���S�5524��q(g�� (򭂯�4X�cOux�\sfwuts�UTS`�i�栜���t�棂Č�? 6�T�!�SA OO+D6����@�����,!��6cp+� igt�t6i��!I0�TW8 ���la��vo58�o�bF� �򬡯i�Xh��!X�k�0Y!8\m6e��!6EC���v��6����������<16�A���A�6s�����U�g�T|ώ���r1"�qR��˔Z4�T��@���,#�eZp)g� ���<ONO0���uJ���tCR;��F�a� x�St�f��prds�uchk �1��2H&&?���t��*D%$ �r(�✑�娟:r���'�s�qO��<sc�rc�C�\At�trldJ"o�\�V�����Paylo�n�firm�l�!�87��7��A�3ad�! �?ވI�?p4lQ��3��3"�q��x pl�`���d7��l�calC�uDup���;��mov��<���initX�:s�8O��a�r4 ��r�67A4|�e Ge?neratiڲ����7g2q$��g R� (Sh��c �,|�bE��$Ԓ\��:�"��4��4X�4�. sg��5�ЌF$d6"e�!p "SHAP�TQ ongcr pGC��a(�&"� ��"GD�A¶��r6�"axW�/�$dataX<:s�"tpad��[q�%tput;a__O7@;a�o8�1�yl+s�Ar�?�:�#�?�5x�?�:c O�:y O�:�$IO�s`O%g�qǒ��?�@0\��"o�j9�2;!�Ppl.Co�llis�QSkip#��@5��@J��D���@\ވ�C@X�7ҥ�7�|s2��pt7cls�LS�DU��k?�\_ ets�`�< \�Q��@����`dcKqQ�FC�;��J,�n��` (���4eN����T �{���'j(�c�q����/IӸaȁ��̠H������зa�e�\mcclmt �"CLM�/��� moate\��lmp�ALM�?>p7qm!c?����2vm�q��8%�3s��_sv90�_x_msu�2L^va_� K�o�{in�8�(3r<�c_logpr��rtrcW񊬯 �v_3�~yc0��d�<�te���der$cCe� Fiρ�R��Q��?�l�enter ߄|��(Sd��1ثTX�+fK�r�a9�9sQ9+�5�r\�tq\� "FND�R���ST�Dn$LANG.�Pgui��D⠓0�S������sp�!ğ֙uf�ҝ�s����$�����e+�=���� �����������w�H�r\fn_�ϣ��$`�x�tcpma��-� TCP�����R638 R�Ҡ�V�38��M7p,�� �Ӡ�$Ӡ�8p0Р�VSl,�>�tk��99�a ��B3���PզԠ��D�2�����UI��t��� hqB���8��������p����re�ȿ��exe@4φ�B���e388�ԡG�rmpWX���var@�φ�3 N�����vx�!ҡ��~q�RBT $c�OPTN a�sk E0��1�R� MAS0�H59}3/�96 H50�Vi�480�5�H0Ԉ�m�Q�K��7�0�g�Pl�h0ԧ�2�OR�DP��@"��t/\mas��0�a�� "�ԧ�����k�գR����ӹ`m��b��&7�.f��u�d��}r��splayD��E���1w�UPDT� Ub��887 (&��Di{���v�Ӛ� �Ԛ⧔��#�B��㟳>��o  ����a�䣣��60q��B��|���qscan���B���ad@�������q`�䗣�#�p�К�`2�� vlv ��Ù�$�>�b����! S��Easy</К�Util���>��511 J���r��R7 ��Nor֠>��inc),<6Q
�� �`c��"4�[����986FVRx bSo����q�nd6� ���P��4�a\ (��
   �������d��K�rbdZ���men7����- Me`tyFњ�Fb�0�TUaN�577?i3R��\�5�u?��!� n���f������l\mh�Ц�ű8E|hmn�	��B<\O���e�1"�� l!��y���
��\|p����B���Ћmh�@��:. aG!���/�t�5�5�6�!X�l�.us���Y/k)ensubL���eK�h�� �B \1;5g?y?�?�?D���?*rm�p�?Ktbox O2K|?�G��C?A%ds���?1��#� �TR��/��P �4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ăd�Q3t.�P׀al��P+OP517F��IN0a��Q(}g���PESTf3ua@�PB�l�ig�h�6�a�q��P � x9S��`  n�0m�bumpP�Q969g�69�Qq��P0��baAp�@Q� B�OX��,>vche8�s�>vetu㒣^=wffse�3�Ā�]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q8<twaǂ tp�Q҄�Taror Re'cov�b�O�P�642����a�q���a⁠QErǃ�Qr!y�з`�P'�T�`�a�ar������	{'�paok971��71��`m���>�pjot���PXc��C�1�adb �-�ail��nagx���b�QR629�a�Q��b�P  ��
  �P���$$CL[q �����������$�PS_DIGsIT���"�!�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*���1:PRODU�CT�Q0\PGS�TK�bV,n��99�\����$FEAT_IN�DEX��~��� 搠IL�ECOMP ;���)��"��S�ETUP2 <����  �N !�_AP2�BCK 1=�  �)}6/E+%,/i/��W/�/ ~+/�/O/�/s/�/? �/>?�/b?t??�?'? �?�?]?�?�?O(O�? LO�?pO�?}O�O5O�O YO�O _�O$_�OH_Z_ �O~__�_�_C_�_g_ �_�_	o2o�_Vo�_zo �oo�o?o�o�ouo
 �o.@�od�o� ��M�q��� <��`�r����%��� ̏[�������!�J� ُn�������3�ȟW� �����"���F�X�� |����/���֯e��� ���0���T��x��� ���=�ҿ�s�ϗ�@,ϻ�9�b�� P/� 2) *.V1Riϳ�!�*����`������PC�|7�!�FR6:"�"c��χ��T��� ��Lը��ܮx��ﶏ*.F��>� �	�N�,�k��ߏ��STM �����Qа����!�iPen�dant Panel���H��F����4������GIF �������u����JPG&P��<�����	PANE�L1.DT��@������2��Y�G��
3 w�����//�
4�a/�O///�/��
TPEINSO.XML�/����\�/�/�!Cust�om Toolb�ar?�PAS�SWORD/��FRS:\R?? �%Passwo�rd Config�?��?k?�?OH� 6O�?ZOlO�?�OO�O �OUO�OyO_�O�OD_ �Oh_�Oa_�_-_�_Q_ �_�_�_o�_@oRo�_ voo�o)o;o�o_o�o �o�o*�oN�or� �7��m�� &���\�����y� ��E�ڏi������4� ÏX�j��������A� S��w�����B�џ f�������+���O�� �������>�ͯ߯t� ���'���ο]�򿁿 �(Ϸ�L�ۿpς�� ��5���Y�k� ߏ�$� ���Z���~�ߢߴ� C���g�����2��� V����ߌ���?�� ��u�
���.�@���d� �����)���M���q� ����<��5r �%��[� &�J�n�� 3�W���"/� F/X/�|//�/�/A/ �/e/�/�/�/0?�/T? �/M?�??�?=?�?�? s?O�?,O>O�?bO�? �OO'O�OKO�OoO�O _�O:_�O^_p_�O�_ #_�_�_Y_�_}_o�_��_Ho)f�$FIL�E_DGBCK �1=��5`��� ( ��)
SUMMA�RY.DGRo�\�MD:�o�o
`�Diag Sum�mary�o�Z
C?ONSLOG�o�o�a
J�aCon�sole log�K�[�`MEMCHECK@'�o��^qMemory� Data��W��)�qHAD�OW���P��s�Shadow C?hangesS�-c�-��)	FTAP=��9����w`q�mment TB�D׏�W0<�)�ETHERNET�̏�^�q�Z��aE�thernet �bpfigurat�ion[��P��DCSVRFˏ��Ïܟ��q%�� ve�rify all�ߟ-c1PY���DIFFԟ��̟a��p�%��diffc���q��1X�?�Q��� ����X=��CHGD��¯ԯi��px��� ����2`�G�Y�� ��� �GD��ʿܿ�q��p���Ϥ�FY�3h�O�a��� ��(�GD�������y��p�ϡ�0�UPDATES.������[FRS:\������aUpda�tes List����kPSRBWLOD.CM.��\���B��_pPS_ROBOWEL���_�� ��o��,o!�3���W� ��{�
�t���@���d� ����/��Se�� ���N�r � =�a�r� &�J���/� 9/K/�o/��/"/�/ �/X/�/|/�/#?�/G? �/k?}??�?0?�?�? f?�?�?O�?OUO�? yOO�O�O>O�ObO�O 	_�O-_�OQ_c_�O�_ _�_:_�_�_p_o�_ o;o�__o�_�o�o$o �oHo�o�o~o�o7 �o0m�o� �� V�z�!��E�� i�{�
���.�ÏR��� �������.�S��w� �����<�џ`���� ��+���O�ޟH�������8���߯n�����$FILE_��P�R���������� �M�DONLY 1=�4�� 
 � ��w�į��诨�ѿ�� �����+Ϻ�O�޿s� ��ϩ�8�����n�� ��'߶�4�]��ρ�� �߷�F���j����� 5���Y�k��ߏ��� B�����x����1�C� ��g������,���P� ��������?��L�u�VISBCK�R�<�a�*.VD�|�4 FR:\���4 Vis�ion VD file� :Lb pZ�#��Y� }/$/�H/�l/� /�/1/�/�/�/�/�/  ?�/1?V?�/z?	?�? �???�?c?�?�?�?.O �?ROdOO�OO�O;O �O�OqO_�O*_<_�O�`_�O�__%_�_�M�R_GRP 1>�4�L�UC4 w B�P	 ]��ol`�*u����RHB ���2 ��� ��� ���He �Y�Q`orkbIh�oJd�o�Sc�o�oL4���M���J��۴F�5U�aRǼ�%�o�o �D�C4ʿ�C���+�9��8g�=7���}?�?�1�9lq>���?����xq}E�� F@ �r�d�a}�J��NJk��H9�Hu���F!��IP�s�X~�`�.9�<�9�89�6C'6<,�6\b�}B%w�&@�_�BLɟ�A�e�+cA�ei@^��B+@�ATg�C�0��N��PA����� |�ݏx���%���p��A6Β@U��{�v�a����� ��П����ߟ��<��'�hzBH�P a�a`�Q�H�*-�o谯¯�U
6�P=��P=��o�o�B��P5���@�33@���4�m�,�/@UUU��U�~w��>u.�?! x�^��ֿ���3���=[z�=�̽�=V6<�=��=�=$q���~��@8�i�7G��8�D��8@9!�7�ϥ�@Ϣ���:t�@ D�� Cϟ�V��C��P��P'� 6��_V� m�o��To�� xo�ߜo������A� ,�e�P�b����� ��������=�(�a� L���p���������V� ������*��N9r ]������� �8#\nY� }�������/ ԭ//A/�e/P/�/p/ �/�/�/�/�/?�/+? ?;?a?L?�?p?�?�? �?�?�?�?�?'OOKO 6OoO�OHߢOl��ߐ� ���O�� _��G_bOk_ V_�_z_�_�_�_�_�_ o�_1ooUo@oyodo vo�o�o�o�o�o�o Nu�� �������;� &�_�J���n������� ݏȏ��%�7�I�[� "/�描�����ٟ�� �����3��W�B�{� f�������կ����� ��A�,�e�P�b��� �����O�O�O��O �OL�_p�:_������ ���������'��7� ]�H߁�lߥߐ��ߴ� ������#��G�2�k� 2��Vw�������� ���1��U�@�R��� v������������� -Q�u��� r��6��) M4q\n��� ���/�#/I/4/ m/X/�/|/�/�/�/�/ �/?ֿ�B?�f?0� BϜ?f��?���/�?�? �?/OOSO>OwObO�O �O�O�O�O�O�O__ =_(_a_L_^_�_�_�_ ���_��o�_o9o$o ]oHo�olo�o�o�o�o �o�o�o#G2k V{�h���� ���C�.�g�y�`� ���������Џ�� �?�*�c�N���r��� �����̟��)�� M�_�&?H?���?���? �?�?����?@�I�4� m�X�j�����ǿ��� ֿ����E�0�i�T� ��xϱϜ�������� �_,��_S���w�b߇� �ߘ��߼������� =�(�:�s�^���� �������'�9� � ]�o����~������� ������5 YD V�z����� �1U@yd ��v�����/Я */��
/�u/��/�/ �/�/�/�/�/??;? &?_?J?�?n?�?�?�? �?�?O�?%OOIO4O "�|OBO�O>O�O�O�O �O�O!__E_0_i_T_ �_x_�_�_�_�_�_o �_/o��?oeowo�oP� �oo�o�o�o�o+ =$aL�p�� �����'��K� 6�o�Z������ɏ�� 폴� ��D�/ / z�D/��h/ş���ԟ ���1��U�@�R��� v�����ӯ������ -��Q�<�u�`���`O �O�O���޿��;� &�_�J�oϕπϹϤ� �������%��"�[� F��Fo�ߵ����ߠo ��d�!���W�>�{� b������������ ��A�,�>�w�b��� �������������=��$FNO ����\��
F0�l q  FLAG�>�(RRM_C�HKTYP  r] ��d �] ���OM� _MI�N� 	���� ��  XT SSB_CFG ?\ �����OTP�_DEF_OW � 	��,IR�COM� >�$G�ENOVRD_D�O��<�lTH�R� d�dq_�ENB] qR�AVC_GRP s1@�I X( / %/7//[/B// �/x/�/�/�/�/�/? �/3??C?i?P?�?t? �?�?�?�?�?OOO�AO(OeOLO^O�OoR�OU�F\� ��,�B,�8�?���O�O�O	_|_���  DE_��Hy_�\@@m_B��=�vR/��I�O�SMT�G�SUoo|&oRHOSTC�s1H�I� ���zMSM�l[�bo�	127�.0�`1�o  e�o�o�o#z�o�FXj|�l60s	�anonymou�s�������QZao�&�&��o �x��o������ҏ� 3��,�>�a�O�� ��������Ο�U%�7� I��]����f�x��� �����ү����+� i�{�P�b�t������ ������S�(�:� L�^ϭ�oϔϦϸ��� ���=��$�6�H�Z� ����Ϳs�������� ��� �2���V�h�z� ��߰���������
� �k�}ߏߡߣ���� ����������C�* <Nq�_���� ��-�?�Q�c�eJ ��n����� ��/"/E�X/j/ |/�/�/�%'/ ?[0?B?T?f?x?� �?�?�?�?�??E/W/�,O>OPObO�KDaEN�T 1I�K P�!�?�O  �P �O�O�O�O�O#_�OG_ 
_S_._|_�_d_�_�_ �_�_o�_1o�_ogo *o�oNo�oro�o�o�o 	�o-�oQu8 n������� �#��L�q�4���X� ��|�ݏ���ď֏7����[���B�QUICC0��h�z�۟���1ܟ��ʟ+���2�,���{�!ROUTER|�X�j�˯!PCJOG̯���!192.�168.0.10���}GNAME �!�J!ROBO�T�vNS_CFG� 1H�I ��Auto-started�$/FTP�/���/ �?޿#?��&�8�J� �?nπϒϤ�ǿ��[� �����"�4ߵ&���� ������濜������� ���'�9�K�]�o�� �����������/ �/�/G���k��ߏ��� ����������1 T���Py���� �"�4�	H-|�Q cu�VD��� �/�;/M/_/q/ �/����/
/�/> ?%?7?I?[?*/?�? �?�?�/�?l?�?O!O 3OEO�/�/�/�/�?�O  ?�O�O�O__�?A_ S_e_w_�O4_._�_�_ �_�_oVOhOzO�O�_ so�O�o�o�o�o�o�_ '9Kno�o� ����o*o<oNo P5��oY�k�}����� pŏ׏����0����C�U�g�y���_�T_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
�FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@oG %j%@�_MOV�u����MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�a��ڿ�
��5� ۵MO�~q_DCd~�1PL�_NAME !�<u� �!De�fault Pe�rsonalit�y (from �FD) �4RR2�k! 1j)TEX�)TH��!�AX d�?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�Ox2-?�O�O�O__0_ B_T_f_x_�b<�O�_ �_�_�_�_�_o o2o�DoVoho&xRj" 1�o�)&0\�b, Ӗ9��b�a @oD�  �a?��c�a?�`�a�aA'��6�ew;�	l��b	 �xoJp��`��`	p �<; �(p� �.r� �K�K ���K=*�J���J���JV��k0q`q�P�x�|�� @j�@T;f�r�f�q�ac�rs�I��!�p����p�r� h}�3���´  ���>��ph�`z���꜖"�Jm�!� H�N��ac����dw��  _�  P� Q� }�� |  а��m�Əi}	'� �� �I� ��  ����:��È�È=̣��(�ts�a	����I  �n �@H�i~�ab�Ӌ�b��w��urN0�� � 'Ж�q�p@2?��@����r�q�5�C�pC0C�G@ C����`�
�A1q _  @B�V~�X�
nwB0h�A��p�ӊ�p�`���aDz���֏���Я�	�pv�( �� -��I��0-�=��A�a�we_q��`�p �?�f�f ��m��� ����Ƽuq@tݿ�>1�  P�apv(�`ţ� �=�qxst��?���`�x`�� <
6b<�߈;܍�<��ê<� <G�&P�ό�AO���c1��ƍ�?fff�?O�?&��qt@��.�J<?�`��wi4����dly �e߾g;ߪ�t��p� [ߔ�߸ߣ����� �`���6�wh�F0 %�r�!��߷�1ى�����E�� E�~O�G+� F�!� ��/���?�e�P���t�,��lyBL�cB��E nw4�������+��R ��s�����<����h�Ô�>��I�m0Xj���A�y��weC������Ƀ�#/*/c/N/wi�6����v/C�`� CCHs/`
=$4��<!��!��ܼ�'�3A��A�AR1A�O�^?�$�?���5p±
=�ç>����3�W
=�#�]�n;e�׬a@�����{����<��>(�B��u��=B�0�������	R��zH�F�G����G��H��U`E���C��+��}I#��I��HD��F��E��R�C�j=�>
�I��@H�!�H�( E<YD0w/O*OONO 9OrO]O�O�O�O�O�O �O�O_�O8_#_\_G_ �_�_}_�_�_�_�_�_ �_"oooXoCo|ogo �o�o�o�o�o�o�o 	B-fQ�u� ������,�� P�b�M���q�����Ώ ���ݏ�(��L�7� p�[������ʟ��� ٟ���6�!�Z�E�W�t��#1($1��9��K���ĥ%�����Ư!3�8�x��!4Mgs���,�IB+8�J��a���{�d� d�����ȿ���ڼ%%P8�P�=:G����S�6�h�z���R��Ϯ����������  %�� ��h�Vߌ� z߰�&�g�/9�$�������7����A�8S�e�w�  ��������������2 �F�$�&Gb���������!C���@���8������F� DzN��� F�P D�!������)#B�'�9K]o#?��W�@@v
��8��8��8�.
 v���! 3EWi{�����:� ��ۨ��1��$MSK�CFMAP  ���� ����(.�ONR�EL  ��!9��EXCFE�NBE'
#7%^!F�NCe/W$JOGO/VLIME'dO S"]d�KEYE'�%]�RUN�,�%��SFSPDT�Y0g&P%9#SIG�NE/W$T1MOT��/T!�_CE_�GRP 1p��#\x��?p��?�? �?�?�?O�?OBO �?fOO[O�OSO�O�O �O�O�O_,_�OP__ I_�_=_�_�_�_�_�_�oo�_:o�TC�OM_CFG 1�q	-�vo�o�o
�Va_ARC_b"��p)UAP_CP�L�ot$NOCHE�CK ?	+ �x�%7I [m���������!�.+NO_?WAIT_L 7%6S2NT^ar	+��s�_ERR_129s	)9�� ,ȍޏ��x���&��d�T_MO��t��,� z�*oq�9�P�ARAM��u	+��a�ß'g{��� =?�345678901��,�� K�]�9�i�������ɯۯ��&g������C��cUM_RSP�ACE/�|����$ODRDSP�c�#6p(OFFSET�_CART�o��D�ISƿ��PEN_FILE尨!�ai���`OPTION_�IO�/��PWOR�K ve7s# !��Vż�8� "�e8p�4�p�	 ���p���<���RG_D?SBL  ��P#���ϸ�RIEN�TTOD ?�C�� !l�UT_S/IM_D$�"����V��LCT �w}��6��a[�1�_�PEXE�j�RAATvШ&p%� ��2^3�j)TEX)TH}�)�X d3� ������%�7�I�[� m�����������@���!�3�E���2�� u���������������c�<d�ASe w���������Ǎ�^0OUa0o�(��(�����u2, ����O H @D� M [?�aG?��cc�D][�Z��;�	ls��xJ���������<w ��� ���ڐH(��H3k�7HSM5G�2�2G���Gp
1͜�'f�/-,�ڐCR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t�!�/ �/�"t�32����/6  ���P%�Q%��
%�|T��S62�q?'e	'� � �2�I� �  ���+==���г?�;	�h	�0�I�  �n @@�2�.��Ov;��ٟ�?&gN�]O  '�'�uD@!� C�C�A@F#H!�/�O�O sb�
���@�@"��@�e0@B�QqA�0Yv: �13Uwz$oV_�/z_e_��_�_	��( ?�� -�2�1 �1ta�Ua�c���:A�-���.  �?��ff���[o"o�_U�`oX�0A8���o�j�>�1  Po�V( ���eF0�f�Y���^L�?����xb�0@<
6b<���;܍�<����<� <�&�,/aA�;r�@|Ov0P?fff?�0�?&ip�T@�.�{r�J<?�` �u#	�Bdqt�Yc� a�Mw�Bo��7� "�[�F��j������� ُ����3�����,���(�E�� �E��3G+� F��a��ҟ�����@,��P�;���B�pAZ�>��B��6�<Oί D���P��t�=���a��s�����6j�h��<7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�%?��?���������#	Ę��P �N|F|CH���Ŀ�������@I�_�'��3A�A�AR�1AO�^?��$�?��������
=ç>�����3�W
=�s#� U��e���B���@��{�����<���(��B�u���=B0�������	�b�H�F��G���G���H�U`E����C�+��I�#�I��H�D�F��E���RC�j=[�
�I��@H��!H�( E<YD0߻��� ������� �9�$�]� H�Z���~��������� ����#5 YD} h������� 
C.gR�� �����	/�-/ /*/c/N/�/r/�/�/ �/�/�/?�/)??M? 8?q?\?�?�?�?�?�? �?�?O�?7O"O[OmO XO�O|O�O�O�O�O�O��O�O3_Q(���ٙ��b��gUU���W_i_2�3��8��_�_2�4Mgqs�_�_�RIB+�_��_�a���{�miGo5okoYo�o�}l��P'rP�nܡ ݯ�o=_�o�_�[R?Q�u���  �p���o� �/��S��z
uүܠ�������ڱ����એ�����   /�M�w�e��������l�2 F�$��Gb��t��a�`�p�S�C�y�@p�5�G��Y�۠F� Dz��� F�P �D��]����پ���ʯܯ� ��~�?_���@@�?��K�K���K���
 �|����� ��Ŀֿ�����0��B�T�fϽ�V� ����{��1��$P�ARAM_MEN�U ?3���  �DEFPULSE�r�	WAITT�MOUT��RC�V�� SHE�LL_WRK.$�CUR_STYLv��	�OPT�N�PTB4�.�C�R_DECSN�� �e��ߑߣ������� ����!�3�\�W�i��{���USE_P�ROG %��%������CCR����e����_HOST7 !��!��:����T�`�V��/��X����_TIME���^��  ��GDEBUG\�˴��GINP_FLMSK����Tfp����WPGA  �����)CH����TYPE������� ���� -? hcu����� ��//@/;/M/_/ �/�/�/�/�/�/�/�/�??%?7?`?��WO�RD ?	=	�RSfu	PNeSUԜ2JOK��DRTEy�]TR�ACECTL 1�x3��� ��`B &�`��`�>�6DT Qy�3�%@�0D �{ �c�a�:@V�@BR� 2ODOVOhOzO�O�O�O��O�O�O�O
__.Z
<TDT,Sb_t_�_ �Z]_�SM �R._@_*RXN\L�
o�[ "c�WBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟���`� �2�D�V�.I v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� j����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o��o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ����������*��$PGT�RACELEN � )�  ���(��>�_�UP z��e�m�u�Y�n��>�_CFG {�m�W�(�n����PЬ� ��DEF�SPD |��l'�P��>�IN�пTRL }���(�8��IPE_C�ONFI��~m�O�mњ���\��>�LID�����=�GRP 1���W��)�A ����&ff(�A�+33D�� D�]� CÀ A)@1��Ѭ(�d�Ԭ����0�0�� 	 �1��1��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P; t_�������  Dz (�
H�X~i� �����/�/�D///h/S/�/��
�V7.10bet�a1��  �A�E�"ӻ��A (�� ?!G�^�!>���"�����!���!BQ��!A\� �!���!*2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?O O:O%O7OpO[O�OO �O�O�O�O�O_�O6_ !_Z_E_~_i_�_�_�_ �_�_�_'o2o�_Vo AoSo�owo�o�o�o�o �o�o.R=vx1�/�#F@ �y �}��{m��y=�� 1�'�O�a��?�?�?�� ����ߏʏ��'�� K�6�H���l�����ɟ ���؟�#��G�2� k�V���z�������� o��ίC�.�g�R� d����������п	� ��-�?�*�cώ�� �Ϯ������B� ;�f�x�������DϹ� �߶��������7�"� [�F�X��|����� ������!�3��W�B� {�f��������� ��� ��/S>wb t������ =OzόϾψ� ���ϼ� /.�'/R� d�v߈߁/0�/�/�/ �/�/�/�/#??G?2? k?V?h?�?�?�?�?�? �?O�?1OCO.OgORO �OvO�O�O���O�O�O __?_*_c_N_�_r_ �_�_�_�_�_o�_)o Tfx�to��� /�o/>/P/b/ t/mo�|��� ����3��W�B� {�f�x�����Տ���� ���A�S�>�w�b� ���O��џ������ +��O�:�s�^����� ��ͯ���ܯ�@oRo do�o`��o�o�o��ƿ �o���*<N�Y� �}�hϡό��ϰ��� �����
�C�.�g�R� ��v߈��߬�����	� ��-��Q�c�N�ﲟ ���l�������� ;�&�_�J���n����� ������,�>�P�: L���������� ��(�:�3��0i T�x����� /�///S/>/w/b/ �/�/�/�/�/�/�/? ?=?(?a?s?��?�? X?�?�?�?�?O'OO KO6OoOZO�O~O�O�O �O�O*\&_8_r����_�_��$P�LID_KNOW�_M  ��� Q�TSV� ���P��?o"o4o �OXoCoUo�o R�S�M_GRP 1�T�Z'0{`�@�`)uf�e�`
�5�  �gpk'P e]o�����`�����SMR�cŅ�mT�EyQ}?  yR����������폯� ��ӏ�G�!��-��� ��������韫���ϟ �C���)������������寧���QST^�a1 1��)����P0� A  4��E2�D�V�h����� ��߿¿Կ���9�� .�o�R�d�vψ��Ϭ�(�����2�0� Q'�<3��3�/�A�S��4l�~ߐߢ߂�5���������6 
��.�@��7Y�k�}���8�������~�MAD  �)��PARN_UM  !�}o\+��SCHE� S��
��f���S��UP�Df�x��_CMP_�`H�� ��'�UER_C;HK-���ZE�*<RSr��_�Q_#MOG���_�X��_RES_G�� !���D�>1b U�y�����@/�	/���� +/�k�H/g/l/��� �/�/�/�	��/�/�/ �X�?$?)?���D? c?h?����?�?�?��V 1��U�ax�@�c]�@t@(@�c\�@�@D@�c[�*@��THR_INRr�J�bz�Ud2FMASS?O� ZSGMN>OqCM�ON_QUEUE� ��U�V P~P UX�N$ UhN�FV�@END�A��I�EXE�O�E��BE��@�O�COPTIO��G��@PROGR�AM %�J%��@�?���BTASK�_IG�6^OCFG� ��Oz��_�PD�ATA�c��[@Ц2=�DoVohozo �j2o�o�o�o�o�o�);M jINFO[��m��D� �������1� C�U�g�y���������@ӏ���	�dwpt�l� )�QE DIT� ��_i��^WE�RFLX	C�RG�ADJ �tZA	�����?נʕFA��?IORITY�GW}���MPDSPNQ�����U�GD��O�TOE@1�X�� (!AF:@E�� c�Ч!tc�pn���!ud|����!icm����?<�XY_�Q��X���Q)� *0�1�5��P��]� @�L���p�������� ʿ��+�=�$�a�H��ϗ�*��PORTT)QH��P�E���_CARTREP�PX��SKSTA��H�
SSAV�@��tZ	2500H863���_x�
�'�U�X�@�swP�tS�ߕߧ���URGeE�@B��x	WF��#DO�F"[W\��������WRUP_DELAY �X�>��R_HOTqX	B�%�c���R_NORMALq^R��v�SEMI�����9�_QSKIP'��tU;r�x 	7�1� 1��X�j�|�?�tU�� ������������ $J\n4��� �����4F X|j���� ���/0/B//R/�x/f/�/�/�/tU�$�RCVTM$��D]�� DCR'����Ў!BR�B�I-�Ce�?�7�{7���;����:��������Xs��%�#:�o?�� <
�6b<߈;����>u.�??!<�&�?h? �?�?�@>��?O O2O DOVOhOzO�O�O�O�O �O�?�O�O__@_+_ =_v_Y_�_�_�?�_�_ �_oo*o<oNo`oro �o�o�o�_�o�o�o�o �o8J-n��_ �������"� 4�F�X�j�U������ ď���ӏ���B� T��x���������ҟ �����,�>�)�b� M������������ï կ�Y�:�L�^�p��� ������ʿܿ� �� ��6�!�Z�E�~ϐ�{� �ϗ�����-�� �2� D�V�h�zߌߞ߰��� ������
���.��R� =�v��k������ ����*�<�N�`�r� ������������� ��&J\?�� ������"�4FXj|��!G�N_ATC 1��	; AT�&FV0E0��ATDP/6/�9/2/9�A�TA�,A�T%G1%B96}0�+++��,�H/,�!IO�_TYPE  �%�#t�REFPOS1 1�V+� x�u/� n�/j�/
=�/�/�/ Q?<?u??�?4?�?X?x�?�?�+2 1�V+�/�?�?\O�?�O�?�!3 1�O*O<O�vO�O�O_�OS4 1��O�O�O_�_t_|�_+_S5 1�B_�T_f_�_o	oBo�_S6 1��_�_�_5o�o�o�oUoS7 1�lo~o�o�oH3l>�oS8 1��%_���SM�ASK 1�V/ � 
?�M��XNO�S/�r������!MOTE  n��$��_CFG �����q���"PL_RA�NG�����POW_ER ������SM_DRYP_RG %o�%��P��TART ���^�UME_P�RO-�?����$_E�XEC_ENB � ���GSPD���Րݘ��TDB���
�RM�
�MT�_'�T����O�BOT_NAME� o����O�B_ORD_NU�M ?�b!�H863  a�կ����PC_TIMEO�UT�� x�S2�32Ă1�� �LTEACH PENDAN���w��-���Maintena�nce Consȡ��s�"���KCL/Cm��

����t�ҿ No Use-��Ϝ��0�NPO�򁋁���.�CH_�L������q	���s�MAVAILȶ����糅��SPACE1 2��, j�߂�D��s��߂� �{S�8�?�k�v�k�Z� ���ߤ��ߚ� �2� D���hߊ�|��`��� ������� �2� D��h��|���`���������y���2�� ��0�B���f������{���3 );M_�� ����/� /44FXj|*/� ��/�/�/?(??=?5Q/c/u/�/�/G? �/�/�?O�?$OEO,OZO6n?�?�?�?�? dO�?�?_,_�OA_b_I_w_7�O�O�O�O �O�_�O_(oIoo^oofo�o8�_�_�_ �_�_�oo6oEf)�{���G ��o� ���
M� ���*�<� N�`�r�������w��@�o�収���d.� �%�S�e�w������� ����Ǐَ���Θ8� +�=�k�}�������ů ׯ͟����%�'�X� K�]���������ӿ忀�����#�E�W�; `� @���@����x�����\�e� ����������R�d� ��8�j߬߾߈ߒߤ� ���������0�r�� ��X������������8����
�ύ��_MODE  ��{��S ��{|�2�0�����3��	S|)CWO�RK_AD��${��+R  �{��`� �� _INOTVAL���d����R_OPTION�� ��H VA�T_GRP 2���up(N�k|�� _�����/0/ B/��h�u/T� }/�/ �/�/�/�/�/?!?�/ E?W?i?{?�?�?5?�? �?�?�?�?O/OAOO eOwO�O�O�O�OUO�O �O__�O=_O_a_s_ 5_�_�_�_�_�_�_�_ o'o9o�_Iooo�o�o Uo�o�o�o�o�o�o 5GYk-��� u�����1�C� �g�y���M�����ӏ 叧�	��-�?�Q�c� ��������������ǟ�;�M�_�����$SCAN_TI�M��_%}�R ��(�#((��<04Jd d 
!D�ʣ��u�/���V��U��25�$��@�d5�P�g��]	���������d�d�x�  P���� ��  8�� ҿ�!���D��$�M�_�qσϕϧ� ���������ƿv��F�X��/� ;�ob���pm��t�_�DiQ̡  � l�|�̡ĥ���� ���!�3�E�W�i�{� ������������� �/�A�S�e�]�Ӈ� ������������ );M_q��� ����r��� j�Tfx���� ���//,/>/P/ b/t/�/�/�/�/�/�%�/  0��6��!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O*�O�O �O�O__+_=_O_a_ s_�_�_�_�_�_�_�_ oo'o9oKo�O�OJ �o�o�o�o�o�o�o  2DVhz�� �����
�7?  ;�>�P�b�t��� ������Ǐُ���� !�3�E�W�i�{�������ß �ş3�ܟ ��&�8�J�\�n������������ɯ��v��,� ��+�	12345�678�� 	�
 =5���f�x�������������
� �.�@�R�d�vψϚ� ៾���������*� <�N�`�r߄߳Ϩߺ� ��������&�8�J� \�n�ߒ������� �����"�4�F�u�j� |��������������� 0_�Tfx� ������ I>Pbt��� ����!/(/:/ L/^/p/�/�/�/�/�/�/�2�/?�#/�9?K?]?�iCz � Bp˚   刅h2��*�$S�CR_GRP 1��(�U8(�\�xd�@� � ��'�	 �3�1�2�4(1 *�&�I3�F1OOXOn}m��D�@��0ʛ)���HUK�L�M-10iA 7890?�90;��F~;�M61C D�P:�CP��1
\&V�1	�6F��CW�9)A7Y	(R�_�_�_�_4�_�\���0i^ �oOUO>oPo#G�/ ���o'o�o�o�o�oB�0�rtrAA�0*  @蠈Bu&Xw?��ju�bH�0{UzAF@ F�`�r��o�� ���+��O�:�s� �mBqrr����������B�͏b����7�"� [�F�X���|�����ٟ ğ���N���AO�0�B�CU
L���E�jqBq�>�q��$G@��@pϯ B����G�I
E�0EL_D�EFAULT  ��T���E��MIPOWERFL  
Ex*��7�WFDO�� *��1ERVE�NT 1����`(�� L!D?UM_EIP��>���j!AF_I�NE�¿C�!FIT������!o�:� ��a�!�RPC_MAIN�b�DȺPϭ�t�VI�S}�Cɻ����!�TP��PU�ϫ�d���E�!
PMON?_PROXYF߮�Ae4ߑ��_ߧ�f�����!RDM_S�RV�߫�g��)�!#R�Iﰴh�u�K!
v�M�ߨ�id����!RLSYN�C��>�8���!�ROS��4��4 ��Y�(�}���J�\��� ����������7�� ["4F�j|� ���!�Ei�o�ICE_KL �?%� (%SVCPRG1n >���3��3��"�4//�5./3/"�6V/[/�7~/�/���D�/�9�/�+ �@��/��#?�� K?��s?� /�?� H/�?�p/�?��/O ��/;O��/cO�? �O�9?�O�a?�O� �?_��?+_��?S_ �O{_�)O�_�QO �_�yO�_��Os� ���>o�o}1�o�o �o�o�o�o�o; M8q\���� �����7�"�[� F��j�������ُď ���!��E�0�W�{� f�����ß���ҟ� ��A�,�e�P���t���������ί�y_�DEV ���MC:��_!�OUT���2��REC 1q�`e�j� �	 �����˿��p�ڿ��
 �`e ���6�N�<�r�`ϖ� �Ϧ��Ϯ�������&� �J�8�n߀�bߤߒ� �߶�������"��2� X�F�|�j������� ��������.�T�B� x�Z�l����������� ��,P>`b t������ (L:\�d� ���� /�$/6/ /Z/H/~/l/�/�/�/ �/.��/?�/2? ?V? D?f?�?n?�?�?�?�? �?
O�?.O@O"OdORO �OvO�O�O�O�O�O�O __<_*_`_N_�_�_ x_�_�_�_�_�_oo 8oo,ono\o�o�o�o �o�o�o�o�o " 4jX����� �����B�$�f� T�v������������ ؏��>�,�b�P�r����p�V 1�}� 1P
�ܟ�o����TYPE\��HE�LL_CFG �.�F�͟  x	�����RSR�� ����ӯ������� ?�*�<�u�`������������  ��2�D���Q̊\�ҰM�o�p�)�d��2Ұd]�KϾ:�HK 1�H� u�������A� <�N�`߉߄ߖߨ��� ��������&�8��~=�OMM �H����9�FTOV_E�NB&�1�OW_?REG_UI����IMWAIT��\a���OUT�������TIM������VAL����_U�NIT��K�1�MO�N_ALIAS �?ew� ( he�#����������Ҵ ��);M��q� ���d�� %�I[m�< ������!/3/ E/W//{/�/�/�/�/ n/�/�/??/?�/S? e?w?�?�?F?�?�?�? �?�?O+O=OOOaOO �O�O�O�O�OxO�O_ _'_9_�O]_o_�_�_ >_�_�_�_�_�_�_#o 5oGoYokoo�o�o�o �o�o�o�o1C �ogy��H�� ��	��-�?�Q�c� u� �������ϏᏌ� ��)�;��L�q��� ����R�˟ݟ��� ��7�I�[�m��*��� ��ǯٯ믖��!�3� E��i�{�������\� տ�����ȿA�S� e�wω�4ϭϿ����� �����+�=�O���s� �ߗߩ߻�f������ �'���K�]�o��� >����������#� 5�G�Y��}����������n��$SMON�_DEFPRO ������� *S�YSTEM*  �d=��RECA�LL ?}�� �( �}
xyz�rate 61 �*.* virt�:\tmpbac�k\9 =>ins�piron:2260 Zas���  }.N3400 HZ����3copy f�rs:orderfil.dat<@�as��� *.mdb:9�Y���/�	/.@em=pQ992 �o/�/�/�'.&*.d B/T'V/�/�/?�-	��/�/�/n?�?�?� �W4G?Y?�?�?O�	2./@O,`OrO�O�O�)�IO�3XO�O�O,_�
-x.D:�<@O,�Om__�_�..Ua6_H_2 ]_�_ o o%O7O�O�Olo~o�o �O�O�OYo�o�o!_ 3_�_W_hz��_�_ B�_��
�o/oAo Sod�v�����oH��o ����+�O`� r������:��_�� ��'?��˟ݟn���x����	1844� Y�����!3����� a�s������E���Y� ���ϡ�3�F�£ݿ nπϒ�%&��?ϼ�^� ����&�8�����m�pߑߤ��
620Ư X������ �2Թ������n���߷	5512G�Y������!� 3�����a�s������� E���Y�����!�3� F�����n����6 HZ_�'�9� ��]n������� [��/#5�Y j/|/�/��D/��/ �/?1�Uf?x? �?��J?��?�?O�N�$SNPX_�ASG 1�����9A�� P 0 '�%R[1]@1�.1O 9?�#3% dO�OsO�O�O�O�O�O �O __D_'_9_z_]_ �_�_�_�_�_�_
o�_ o@o#odoGoYo�o}o �o�o�o�o�o�o* 4`C�gy�� �����	�J�-� T���c�������ڏ�� ���4��)�j�M� t�����ğ������ݟ �0��T�7�I���m� �������ǯٯ��� $�P�3�t�W�i����� ���ÿ����:�� D�p�Sϔ�wω��ϭ� �� ���$���Z�=� dߐ�sߴߗߩ����� �� ��D�'�9�z�]� ���������
��� �@�#�d�G�Y���}� ������������* 4`C�gy�� ����	J- T�c����� �/�4//)/j/M/ t/�/�/�/�/�/�/�/�?0?4,DPARAoM �9ECA_ �	��:P�4��0$HOFT_�KB_CFG  �p3?E�4PIN_�SIM  9K��6�?�?�?�0,@RV�QSTP_DSBº>�21On8J0SR� ��:� &� MULTIR�OBOTTASK�=Op3�6TOP�_ON_ERR � �F�8�APTN� �5�@�A�BRING_�PRM�O J0V�DT_GRP 1y�Y9�@  	�7 n8_(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 Dkhz���� ���
�1�.�@�R� d�v���������Џ�� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\������� ����ȯگ����"� I�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� tߛߘߪ߼������� ��(�:�a�^�p�� ���������� �'� $�6�H�Z�l�~��������������3VPRG_COUNT�6���A�5ENB��OM=�4J_U�PD 1��;8  
p2��� ��� )$6H ql~����� /�/ /I/D/V/h/ �/�/�/�/�/�/�/�/ !??.?@?i?d?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_�_�_Y?SDEBUG" � ��Pdk	�PSP_�PASS"B?~�[LOG ��+m�P�X�_�  �g�Q
M�C:\d�_b_M�PCm��o�o��Qa�o �vfSAV �m:dUb�U�\gSV�\TE�M_TIME 1]�� (�P��T���o	T1SVGgUNS} #'k��spASK_OPTION" �go�spBCCFG 3��| �b�{�}`����a&� �#�\�G���k����� ȏ������"��F� 1�j�U���y���ğ�� �ӟ���0��T�f��UR���S���ƯA� ����� ��D��nd� �t9�l���������ڿ ȿ�����"�X�F� |�jϠώ��ϲ����� ����B�0�f�T�v� xߊ��ߦؑ������ �(��L�:�\��p� ����������� � 6�$�F�H�Z���~��� ����������2  VDzh���� �����4Fd v������ //*/�N/</r/`/ �/�/�/�/�/�/�/? ?8?&?\?J?l?�?�? �?�?�?�?�?�?OO "OXOFO|O2�O�O�O �O�OfO_�O_B_0_ f_x_�_X_�_�_�_�_ �_�_oooPo>oto bo�o�o�o�o�o�o�o :(^Lnp �����O��$� 6�H��l�Z�|����� Ə؏ꏸ����2� � V�D�f�h�z�����ԟ ����
�,�R�@� v�d���������ίЯ ���<��T�f��� ����&�̿��ܿ�� &�8�J��n�\ϒπ� �Ϥ����������4� "�X�F�|�jߌ߲ߠ� ����������.�0� B�x�f��R������� �����,��<�b�P� ������x��������� &(:p^� ������  6$ZH~l�� ������/&/D/ V/h/��/z/�/�/�/��/�&0�$TBC�SG_GRP 2���%� � �1 
 ?�  /?A?+?e? O?�?s?�?�?�?�?�;�23�<d,� �$A?1	 H�C���6>���@E�5CL  B�p'2^OjH4J��B�\)LFY  A��jO�MB��?�IBl�O�O�@�JG_�@�  D	�15_ __$YC-P{_F_`_j\	��_�]@0�>�X�U o�_�_6oSoo0o~o�o�k�h�0	�V3.00'2	�m61c�c	*`�`�d2�o�e>�JC20(�a�i ,p�m�-  �0�����omvu1JCFG� ��% 1 �#0vz��rBrv�x����z � �%��I�4�m�X� ��|��������֏� ��3��W�B�g���x� ����՟������� �S�>�w�b�����'2 A ��ʯܯ������ E�0�i�T���x���ÿ տ翢����/��?� e�1�/���/�ϜϮ� �������,��P�>� `߆�tߪߘ��߼��� �����L�:�p�^� ������������  �6�H�>/`�r���� ������������  0Vhz8��� ���
.�R @vd����� ��//</*/L/r/ `/�/�/�/�/�/�/�/ �/?8?&?\?J?�?n? �?�?�?�?���?OO �?FO4OVOXOjO�O�O �O�O�O�O__�OB_ 0_f_T_v_�_�_�_z_ �_�_�_oo>o,obo Poroto�o�o�o�o�o �o(8^L� p������� $��H�6�l�~�(O�� ��f�d��؏���2�  �B�D�V�������n� ���ԟ
���.�@�R� d����v�������� Я���*��N�<�^� `�r�����̿���޿ ��$�J�8�n�\ϒ� �϶Ϥ�������ߊ� (�:�L���|�jߌ߲� �����������0�B� T��x�f������ �������,��P�>� t�b������������� ��:(JL^ ������ � 6$ZH~l� �^���dߚ // D/2/h/V/x/�/�/�/ �/�/�/�/?
?@?.? d?v?�?�?T?�?�?�? �?�?OO<O*O`ONO �OrO�O�O�O�O�O_ �O&__6_8_J_�_n_ �_�_�_�_�_�_�_"o oFo��po�o,oZo �o�o�o�o�o0 Tfx�H��� ����,�>��b� P���t���������Ώ ��(��L�:�p�^� ������ʟ���ܟ�  �"�$�6�l�Z���~� ����دꯔo��&� ЯV�D�z�h������� Կ¿��
��.��R��@�v�dϚτ�  ���� ��������$TBJOP_�GRP 2ǌ���  �?�������������x�JBЌ��9� �< �X�ƞ�� @���	� �C�� t�b�  C����>ǌ�͘Րդ�>���йѳ33=��CLj�fff?>��?�ffBG���Ќ�����t�ц�>;�(�\)�ߖ��E噙�;��h{CYj��  @h�~�B�  A�����f��C�  D�hъ�1��O��4�N����
:�/��Bl^��j�i��l�l����Aə�3A�"��D���Ǌ=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������<$�6�>B�\��T����Q�tsx�@g33@���C����y�1����>��Dh����������O<{�h�@i�  ��t��	� ��K&�j� n|���p�/��/:/k/�ԇ����!��	V3.0}0J�m61cIԃ*� IԿ��/�'� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�I�!CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;��;Q�UT,8�4` *���?�2���3\�X/�O��ESTPAR�S  ��	���H�R@ABLE 1%����0��
H�7Q 8��9
G
H
H�����
G	
H

H�
HYE��
H
H:
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_�^:BS _� �JGoYo ko}o�o�o�o�o�o�o �o1CUgy ����`#oRL�y�_ �_�_�_�O�O�O�O�O�X:B�rNUM  ����P���� V@P:B_CF�G ˭�Z�h�@���IMEBF_T�T%AU��2@�VE�RS�q��R {1���
 (�/����b� ����J� \���j�|���ǟ��ȟ ֟�����0�B�T�@��x�������2�_����@�
��MI_�CHAN�� � >��DBGLV����������ETHE�RAD ?��
O�������h������ROUT�!���!������SN�MASKD��U�255.���#������OOLOFS_�DI%@�u.�OR�QCTRL � ����}ϛ3rϧϹ��� ������%�7�I�[��:���h�z߯�APE?_DETAI"�G��PON_SVOF�F=���P_MON� �֍�2��S�TRTCHK ��^�����VTCOMPAT��O������FPROG �%^�%MULTIROBOTTݱx���9�PLAY&H���_INST_M�ް ������US8�q��LCK���QUICKME��=���SCREZ�}G�tps� @���u�z����_���@@n�.�SR_GR�P 1�^� �O����
��@+O=sa�� ��
m������ L/C1gU� y�����	/��-//Q/?/a/�/	1234567�0h�/�/@Xt�1����
 �}ipn�l/� gen.htm�? ?2?D?V?�`Panel� setupZ<}�P�?�?�?�?�?�? �??,O>OPObOtO �O�?�O!O�O�O�O_ _(_�O�O^_p_�_�_ �_�_/_]_S_ oo$o 6oHoZo�_~o�_�o�o �o�o�o�oso�o2D Vhz�1'� ��
��.��R�� v���������ЏG����UALRM��G ?9� �1�#� 5�f�Y���}������� џן���,��P���SEV  �����ECFG C��롽�A���   BȽ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �("� ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1`����(�:�'����71�߅�����J�3O���edit���MULTIROBOTTASKt� �'�9�D�=�g�y��� ������P�����	 -?��cu��� �L^�); M�q�������f��f//'/ 9/K/]/`�/�/�/�/ �/�/j/�/?#?5?G? Y?�/�/�?�?�?�?�? �?x?OO1OCOUOgO �?�O�O�O�O�O�OtO �O_-_?_Q_c_u__ �_�_�_�_�_�_�� )o;oMo_oqo�o�_�o �o�o�o�o�o%7 I[m� �� �����3�E�W� i�{������ÏՏ� ������A�S�e�w� ����*���џ���� �ooO�a�s����� ����ͯ߯���'� ��K�]�o��������� F�ۿ����#�5�Ŀ Y�k�}Ϗϡϳ�B��� ������1�C���g� yߋߝ߯���P����� 	��-�?�*�<�u�� ������������ )�;�M���������� ������l�%7 I[������ �hz!3EW i������� v////A/S/e/P����$UI_PA�NEDATA 1������!�  	�}�w/�/�/�/�/?? )?>?V�/i?{?�? �?�?�?*?�?�?OO OAO(OeOLO�O�O�O��O�O�O�O�O_&Y� b�>RQ?V_h_ z_�_�_�__�_G?�_ 
oo.o@oRodo�_�o oo�o�o�o�o�o�o *<#`G��}�-\�v�#�_�� !�3�E�W��{��_�� ��ÏՏ���`��/� �S�:�w���p����� џ������+��O� a���������ͯ߯ �D����9�K�]�o� �������ɿ���Կ �#�
�G�.�k�}�d� �ψ����Ͼ���n��� 1�C�U�g�yߋ��ϯ� ��4�����	��-�?� ��c�J������ ���������;�M�4� q�X����������� %7��[�� �����@� �3WiP�t �����/�// A/����w/�/�/�/�/ �/$/�/h?+?=?O? a?s?�?�/�?�?�?�? �?O�?'OOKO]ODO �OhO�O�O�O�ON/`/ _#_5_G_Y_k_�O�_ �_?�_�_�_�_oo �_Co*ogoyo`o�o�o �o�o�o�o�o-`Q8u�O�O}��@������)� >��U-�j�|������� ď+��Ϗ���B� )�f�M���������������ݟ��XS�K��$UI_PANELINK 1�U�  ��  ��}1�234567890s���������ͯդ �Rq����!�3�E�W� �{�������ÿտm��m�&����Qo�  �0�B�T�f�x�� v�&ϲ���������� ��0�B�T�f�xߊ�"� �����������߲� >�P�b�t���0�� ����������$�L� ^�p�����,�>�����`�� $�0,&� [�XI�m��� ����>P3 t�i��Ϻ�  -n��'/9/K/]/o/ �/t�/�/�/�/�/�/ ?�/)?;?M?_?q?�? �UQ�=�2"��?�? �?OO%O7O��OOaO sO�O�O�O�OJO�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5oGo�_ko}o�o�o �o�oTo�o�o1 C�ogy���� �B�	��-��Q� c�F�����|������ �֏�)��M���= �?��?/ȟڟ��� �"�?F�X�j�|��� ��/�į֯����� 0��?�?�?x������� ��ҿY����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z���� -���������
��. RdG��}� ���c���<�� `r������� �//&/8/J/�n/ �/�/�/�/�/7�I�[� 	�"?4?F?X?j?|?� �?�?�?�?�?�?�?O 0OBOTOfOxO�OO�O �O�O�O�O_�O,_>_ P_b_t_�__�_�_�_ �_�_oo�_:oLo^o po�o�o#o�o�o�o�o  ��6H�l~ a������� �2��V�h�K����� ��1�U
��.� @�R�d�W/�������� П������*�<�N� `�r��/�/?��̯ޯ ���&���J�\�n� ������3�ȿڿ��� �"ϱ�F�X�j�|ώ� �ϲ�A��������� 0߿�T�f�xߊߜ߮� =���������,�>� ��b�t�����+ ������:�L�/� p���e�����������  ��6���ۏ���$UI_QU�ICKMEN  }���}���RESTOR�E 1٩�  �
�8m3\n ���G���� /�4/F/X/j/|/' �/�/�//�/�/?? 0?�/T?f?x?�?�?�? Q?�?�?�?OO�/'O 9OKO�?�O�O�O�O�O qO�O__(_:_�O^_ p_�_�_�_QO[_�_�_ I_�_$o6oHoZoloo �o�o�o�o�o{o�o  2D�_Qcu�o �������.� @�R�d�v��������xЏ⏜SCRE� �?�u1�sc� u2�3��4�5�6�7��8��USER�����T���ksT'���4��5��6���7��8��� NDO_CFG ڱ�  �  � PD�ATE h���None�S�EUFRAME � ϖ��RTOL_ABRT�����ENB(��G�RP 1��	�?Cz  A�~�|��%|�������į֦��X�� UH�X�7�?MSK  K�S��7�N�%uT�%������VISCA�ND_MAXI��I�3���FAILO_IMGI�z �% �#S���IMREG�NUMI�
���S�IZI�� �ϔ�,�ONTMOU4'�K�Ε�&�����a��a���s�FR:\��� � M�C:\(�\LOGnh�B@Ԕ !{��Ϡ�����z �MCV����7UD1 �EX	��z ��PO64_t�Q��n6��PO!�LI�Oڞ�re�V�N�f@`��I�� =	_�SZ�Vmޘ��`�WA�Imߠ�STAT �k�% @��4�F��T�$#�x �2D�WP  ��P� G��=��������_JMP�ERR 1ޱ
�  �p2345678901��� 	�:�-�?�]�c����� ������������$�MLOW�ޘ�����g_TI/�˘'���MPHASE  �k�ԓ� ��SH�IFT%�1 Ǚ��<z��_� ���F/| Se������ �0///?/x/O/a/��/�/�/�/�/�����k�	VSFT1�[�	V��M+3 S�5�Ք p���ſA�  B8[0�[0�Πpg3a1Y2�_3Y�7ME��K�͗q	6e���&%���M���b��	���$��TDINEND3�4��4OH�+�G�1�OS2OIV I�{��]LRELEv�I��4.�@��1_AC�TIV�IT��B��A �m��/_��B�RDBГOZ�YBO�X �ǝf_[���b�2�TI�190.0.�P8�3p\�V254tp^�Ԓ	 �S��_�[b��r�obot84q_   p�9o[�pc�PZoMh�]�Hm�_Jk@1�o�ZA+BCd��k�,���P [�Xo}�o0); M�q����� ���>��aZ�b��_V