��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ����ALRM_�RECOV1   $ALMO�ENB��]ON�i�APCOUPwLED1 $[�PP_PROCE�S0  �1��GPCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y12 � u3�|4|GRG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WAx�471�:OFF_ �N�3DELHLO�Gn25Aa2?i1@N?�� -M��H W+0�$Y �$DB� 6COMW!2MO� 21\D�.	 \rVE��1$F��A{�$O��D�B�CTM�P1_F�E2�G1�_�3�B�2�XD��#
 d $�CARD_EXI�ST4$FSS�B_TYPuAH�KBD_S�B�1A�GN Gn $�SLOT_NUM�JQPREV,DB�U� g1G ;1_ED�IT1 � *1G=� S�0�%$EP�$�OP�AEToE_OKRUS�oP_CRQ$;4x�V� 0LACIw�1�RAPk �1x@M}E@$D�V��Q�Pv�A{oQLv� OUzR ,mAЧ0�!� B� LM�_O�^eR�"CAsM_;1 xr~$ATTR4�NP� ANN�@5I�MG_HEIGH|Q�cWIDTH4�VT� �UU0F_�ASPECQ$�M�0EXP��@A�X�f�CFT ?X $GR� � �S�!�@B@NFL�I�`t� UIREx 3dTuGITCHCj�`N� S�d_L�`2�C�"�`EDlpE
� J�4S�0� �zsa�!ip;G0 �� 
$WARNM��0f�!,P� �s�pN{ST� CORN�"�a1FLTR�uTRkAT� T�p H0ACCa1���{��ORI
`"S={R�T0_S�B�qHG�,I1 [ Thp�"3I9�TY�D(,P*2 �`w@� X�!R*HD�cJ* TC��2��3��4��U5��6��7��8���94nQCO�$ <� $6xK3 1w`�O_M�@�C t� � E#6NGP�ABA� �c��ZQ ���`���@nr���� ��P�0����x�p�PzPb26��4��"J�_R��B�C�J��3�JV P��tBS��}Aw��"~�@(�CP_*0wOFSzR @� �RO_K8���aIT<�3��NOM_�0�1Yĥ3�qPT� �� $���AxP��K}EX�� �0g0�I01��p�
$TF�a��C$MD3��T�O�3�0U� �� K�Hw2�C1|�	EΡg0wE{vF�vF�40CPp@�a2 m
P$A`PU�3N)#�dR*��AX�!sDETAI�3BUFV�p@1� |�p۶�pPIZdT� PP[�MZ��Mg�Ͱj�F[�SIMQSI�"0��A.�t���Pkx Tp�|zM��P�B�FAkCTrbHPEW7�`P1Ӡ��v��MCd�� �$*1JB8�p<�*1DECHښ��H��a� � ~+PNS_EMP��G$GP���,P_���3�p�@Pܤ��TC ��|r��0�s��b�0��� �B���!
���JR|� ��SEGFR���Iv �aR�TkpN&S,�PVF4��� &k�Bv�u �cu��aE�� !2��+�8MQ��E�SIZ�3�����T��P�����aRSINF����Ӏkq��������LpX�����F�CRCMu�3CClpG��p��� O}���b�1�������T2�V�DxIC��C����r����P��{� E�V �zF_��FR�pNB0�?���8���A�! �r� Rx����V�lp�2��aPR�t�,�g
�qRTx #�5�5H"2��uAR���`CX�'$LG�p��B�1 `s�P�t�aA�0{�Уb+0R���tME�`0!BupCrRA 3tCAZ�л�pc�OT�#FC�b�`�`FNp��8�1��ADI+�a %��b�{��p$�pSp�c�`S�P��a,Q�MP6�`Y�3��M�'�pU��aU � $>�TITO1��S�S�!��$�"0�D�BPXWO��!���$SK��2&�@DB�"�"@�;PR8� 
� ����# >�q1M$��$��+�L9!$?(�V�%@?R4�C&_?R4ENE���'~?(�� R�E�pY2(H v�OS��#$L�3$$3R��;3�MV�Ok_D@!V�RO�Scrr�w�S���CR�IGGER2FPA��S��7�ETURN�0B�cMR_��TUrː[��0EWM%���GN>`��RL�A���Eݡ�P�'&$P�t�'�@4a"��C�DϣV�DXQ���4�1��MVGO_A7WAYRMO#�a�w!� CS_)7  `IS#�  �� �s3S�AQ汯 4Rx�ZSW�AQ�p�@r1UW��cTNTV)�5RV
a���|c�éW�ƃ��JB��x0��S�AFEۥ�V_SV>�bEXCLUU�;���ONL��cY�g�~az�OT�a{�HI_V? ��R, M��_ *�0� ��_�z�2� p�QSGO  +�rƐm@��A�c~b���w@��V��i�b�fANNUNXx0�$�dIDY�UABc�@Sp�i�a+ �jr�f�!�pOGIx2,��$F�b�$ѐ�OT�@A $DUMMY��Ft���Ft±� 6U- 7` !�HE�|s��~bc�B@ SUF�FI��4PCA��Gs5Cw6dr� �DMSWU.{ 8!�KEYI��5�TM�1�s�qoA�vINޱw�X� , �/ D��HOST�P!4���<���<�0°<��p<�EM'����Z�� SBL� UL>��0  �	���E�� T�01 ϴ $��9USAMPLо�/����ĺ�$ I@갯 $SUBӄ��w0QS��8���#��SAV������c�S< 9�`�fP�$�0E!� YN_�B�#2 0�`DI��d�pO|�m��#$�F�R_IC� �?ENC2_Sd�3  ��< 3�9����� cgp����4��"��2�A��ޖ5���`ǻ�@Q@�K&D-!�a�AVE�R�q����DSP
���PC_�q��"�x|�ܣ�VALU3��HE�(�M�IP\)���OPPm �CTH�*��S" $T�/�Fb�;�d�����d D�;��16� H(rLL_DU ǀ�a�@��k���֠COT�"U�/��~@@NOAUTO70�$}�x�~�@s���|�C͠��C�� 2p�z�L�� �8H *��L � ���Բ@sv��`�  �� ÿ���Xq��cq��P�q���q��7��8���9��0���1�1� �1-�1:�1G�1�T�1a�1n�2|�2T��2 �2-�2:�U2G�2T�2a�2nʕ3|�3�3� �3�-�3:�3G�3T�3*a�3n�4|�a�����9 <���z�ΓKI����H硵Ba�FEq@{@: ,<��&a? P_P�?��>�����E@�@��QQ��;fp�$TP�$V�ARI����,�UP�2Q`< W�߃TD ��g���`������%����BAC�"= T2����$)�,+r³�p IFI��p�� q M�P"��l@``>>t ;��6����ST����@T��M ����0	�� i���F���������kR�t ����FORCE�UP�b܂FLUS

pH(N��� ��6b/D_CM�@E�7�N� (�v�P��REM� Fa��@(j���
K�	N����EFF/���@IN̆QOV��OV=A�	TROV �DT)��DTMX :e �P:/��Pq��vXpCLN _ �p��@ ��	_|���_T: �|�&PA�QDI���10��0�Y0RQm��_+qH���M���C9L�d#�RIV{�ϓnN"EAR/�IO�#PCP��BR��cCM�@N 1b 3�GCLF��!DY��(��a�#5T�D�G���� �%r�S9S� )�? P(q1�1�`_1"81�1�EC13D;5�D6�GRA���@������PW�ON<2EBUG�S�2�C`gϐ_E �A ��@a �/TERM�5B�5 O�ORIw�0C�51��SM_-`����0D�9TA�9Eܽ5p��UP��Fg� -QϒA�P|�3�@B$SEGGJv� EL�UUSEPNFI��pBx��1x@��4>DC$UF�P��$���Q�@C���G�0T�����SwNSTj�PATۡ<g��APTHJ�A�E*�Z%qB\`F�{E���F�q�pARxPY�aS�HFT͢qA�AX_�SHOR$�>��6 �@$GqPE���O#VR���aZPI@P@$�U?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi� [Y)��G�@R��i�e԰�i�R�!P�uAScYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UaP���P���WOR�@�M��k0SMT��G��GR��3�a�PA�@��p5�'�H� � j�A�T�OCjA7pP]Pp$OPd�O��C�%��p�O!��RE.pR�C�AO�?��Be5pR�EruIx'Q�G�e$PWR) IMdu�RR_$s��5�.�B Iz2H8�=��_ADDRH�H_LENG�B�q�q:��x�R��So�J.�SS��SK������ ��-�SE*���rmSN�MN1K	��j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ���p�Q� ��OUPW3��b_>�I��!q�a1 ��������|��� �����-���:���i+IOX2S=�D�e�x�]���L $��<p�!_OFF[r_�oPRM_��a�TTP_�H��M; (�pOBJ�"�p�G�$H�LE�C|��ٰN � 9�.*�AB_�T��
��S�`�S��LV��K�RW"duHITCOmU?BGi�LO�q����d� Fpk��GpSS� ���HW�h�wA��O.��`I�NCPUX2VISIO��!��¢.�á�<�á-� �IOL]N)�P 87�R'�^[p$SL�bd oPUT_��$dp��Pz �� F_�AS2Q/�$L D���D�aQT U�0]PA������PHY`G灱Z��P4�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp����x��ٶ��UJ���S����NE�WJsOG�G �DIS��b&�KĠ��3T |���AV��`_�CTR<!S^�FLAGf2&�;LG�dU �n�:���3LG_SIZ���ň��=���FD��I����Z �ǳ� �0�Ʋ�@s��-ֈ�-ր=�-���-��0-�ISGCH_��Dq��N?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHrܵ�I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn�a��_BWUFF1XY��PT�$�� �v���f�L6q1YY���P �����pOS1J�2�3���_�>0Z �  ��apiE�*��IDX�d	P�RhrO�+��A&+ST��R��Yz�<!� Y$EK&C K+���Z&m&KF�1[ L��o�0��]P L�6pwq�t^����w��~7�_ \ �`@��瀰�7��#�0C���] ��CLDP|��;eTRQLI�pjd.�094FLGz�0r1R3�DM�R7���LDR5<4R5ORG .���e2(`���V�8.�p�T<�4�d^ �q�P<4��-4R5S�`T00�m��0DFRCL�MC!D�?�?3I@�'��MIC��d_ Yd���RQm�q��DSTB	�  ؏Fg�HAX;b |�H�LEXCESZr���rBMup�a`�@�B;dKrB`��`a��F_A�J��$[�Ot�H0K�db \���ӂS�$MB��LI�Б}SREQUIR��R>q�\Á�XDEB�U���AL� MP�c��ba��P؃ӂ!B�M#ND���`�`d�҆��c�cDC1��IN@�����`@�(h?Nz��@q��o� p@�QP�ST8� e�rL�OC�RI�p�E�X�fA�p��A�AOwDAQP�f X��3ON��[rMF���� �f)�"I��%�e��T�v��FX�@IGG� g �q��"E��0��#���$R�a% ;#7y��Gx��VvCPi�ODATAw�pE:��y��RFЭ�NVh �t $MD�qI�ё)�v+�tń�tH��`�P�u�|��sAN�SW}��t�?�uD��)�b�	@Ði -�@CU��V�T0�eRR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2N�RIN��v�<��'NTE���kE����,��b����_Nl@��ڂ��~�ՆRm�7DIV�DH�@ـ:n�$V��'cv!$��$Z������~�[��o�H �$BEL�Tb��!ACCEL�+��ҡ��IRC��t����T/!���$PS�@#2L� q�Ɣ83������� ��PATH��������3̒Vp�A_�Q�.��4�B�Cᐈ�_M=Gh�$DDQ���G�$FWh��p���m�����b�DE��P�PABNԗROTSPEED����00�J�Я8��@����$USE_��P���s�SY��c�A �kqYNu@Ag��OsFF�q�MOUN�3NGg�K�OL�H�INC*��a��q��Bxj�L@�BENCS���q�Bđ���D��IN�#"I̒��4�\BݠV�EO�w�Ͳ23_UyPE�߳LOWLA���00����D��@�BwP��� �1RCʀ�ƶMOSIV�JRM�O���@GPERC7H  �OV�� ^��i�<!�ZD<!�c@��d@�P��V1�#P͑��L���EW�ĆĸUP������T�RKr�"AYLOA'a�� Q-�(�<�1�8�`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H�����b�DUM2(�S_�BCKLSH_C (���>�=�q�#�U��������2�t�]ACLA�LvŲ�1n�P�C�HK00'%SD�RT�Y4�k��y�1�q_�6#2�_UM$Pj�C�w�_�SCL��ƠLMT_J1_LO�"�@���q��E������๕�幘SPC`��7������PCo�B��H� �PU�m�C/@��"XT_�c�CN_b��N��e���SFu���V�&#����9�(�d��=�C�u�SH6# ��c����1�Ѩ�o�0�0͑
��_�PAt�h�_Ps�W�_10��4֠R�01D�VG�J� L��@J�OGW���ToORQU��ON*ɀMٙ�sRHљ��_	W��-�_=��C��TI��I�I�II�	F�`�JLA.�1[��VC��0�D�BO1�U�@i�B\JRK�U��	@DBL_�SMd�BM%`_D9LC�BGRV��0C��I��H_� �*COS+\�(LN�7+X>$C�9)�I�9)u*c,)�Z2 HƺMY@!�( "�TH&-�)THET=0�NK23I��"l=�A CB6CB=�C�A�B(261C�61�6SBC�T25GT	S QơC��aS$�" �4c#�7r#$DUD�EX�1s�t��B�6䆱�AQ|r�f$NE�DpIB U�\B5��	$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2��&�C�J�&!�VAHV�6H3�YLVhJVuKV��KV�KV�KV�KV�IHAHZF`RXM��wX�uKH�KH�KH�KH��KH�IO2LOAHOT�YWNOhJOuKO�KUO�KO�KO�KO�&�F�2#1ic%�d4GS�PBALANCE�_�!�cLEk0H_�%SP��T&�bc&�b>r&PFULC�hr��grr%Ċ1ky�U�TO_?�jT1T2Cy��2N&�v�ϰ ctw�g�p�0Ӓ~����T��O���� IN�SEGv�!�REV8�v!���DIF�鉳1l�w�1m�0OaB�q
����MIϰ�1��LCHWAR̭���AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|�n��ROBR�CR(����N��'�MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD���ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDX�Р  ��MOR^��t $-�U���)��r�B���  ����Gؒu � $SIMULT ৐~�� ���OBJ�E�` �ADJUS<>�1�AY_Ik���D_����C�_FIF�=�T� ��Ұ ��{��p� �����p�@:��D�FRI��ӥMT��RO� ��E�z��͐OPWO��ŀv0��SYS�BU�@ʐ$SOP�����#�U"��pPgRUN�I�PA��DH�D����_OUb�=��qn�$}�/IMAG��ˀ�0�P�qIM����IN��q���RGOVR!Dȡ:���|�P~���Р�0L_6p���i⦄�RB������ML���EDѐF� ��%N`M*���ⷀ˱�SL�`ŀw x �$OVSL�vS;DI��DEXm�g� e�9w�����V� ~�N���w����Ûǖ���M�\͐�q<�>�� x HˁE�^F�ATUS����C�0àǒ��BTMT����If���4����(�ŀy DˀEz�g���PE�r����8�
���EXE��V���E�Y�$Ժ ŀz �@ˁ��UP{�h�$�p��XN���9x�H��PG"��{ h $SUB��c�@_��01\�_MPWAI��P��&��LO��<�F�p��$RCVFAI�L_C�f�BWD�"�F���DEFSP>up | Lˀ`��D�� U�UNI��S���R`����_L�pP��̐ �	P�ā}��� B�~�о�|��`ҲN�`KE)T��y���P� $��~���0SIZE�] ଠ{���S<�O�R��FORMAT�/p � F���rEM2R��y�UX����@�PLI7�ā � $�P_S�WI����_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W ��U����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�aO�0\H��6@��� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�Hӱt��W�UpS����M��O㵐.'}q��C�g���@ʣ�ߑ��M��AÂ� � $sPY��$WH`'�NGp���H`��Fb`��Fb��Fb��PLM�@��	� 0h�H�{�X��	O��z�Z�eT�M���G� pS��C���O__0_B_�a��_%�� |S����@	 �v��v �@���w�vr��EM��% Z��fr�B�ː��ftPn��PM��QU� �U�Q��Af�wQTH=�HOL��oQHYS�ES�F,�UE��B��O#��  -�P0�|�gAPQ���ʠu���O��ŀ�ɂv�-�A;ӝGROG��a2D��E�Âv�_�ĀZ�INFO&��+����b�Ȝ�OI킍 ((@SLEQ/�#@������o���S`�c0O�0�01E�Z0NUe�_�AUT<�Ab�COPY���(��{��@M��N������1�P�
� ��RG4I�����X_�Pl�C$�����`�W���P��j@�G���E�XT_CYCtb����p��A`h�_NA�!$�\�<��RO�`]�� �s m��POR�㸅����SRVt�)l����DI �T_l� ��Ѥ{�ۧ��ۧ �ۧU5٩6٩7٩8���R�S�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,(@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#q�RQSK;IP�� ĕ�x�-O�`NT!���P_x���ǚ@�b�p 1�1�1Ǹ�?� � ?��>��>�&�>�3�z>�9�J2R;n쐖 4��EX� TQ����ށ�Q����[�KFд�KE�R;DCIf� �U`�X}�R�#%M!*�0��)��$RGEAR_�0IO�TJBFLG��igpERa��TC�݃������2TH2�N��� 1� ��Gq T�0 �����M���`I�b����REF�1��� l�h��ENsAB��lcTPE?@ ���!(ᭀ����Q �#�~�+2 H�W���2�Қ���"�4�F�X�j�3�қ{���P������j�4�Ҝ��@
��.�@�R�j�5�ҁ�u����������� )����6�Ҟ���(:Lj�7�ҟ�o�����j�8�Ҡ��"4F�j�SMSK�� � �+@��E�A��M�OTE�����`�@ "1��Q�IO�5�"%I��P��POWi@쐣  ������X�gpi�쐤��Y"$�DSB_SIGN�4A�Qi�̰C��>%S�232%�Sb�iDEVICEUS#|�R�RPARIT򱾈!OPBIT�Q���OWCONTR`��Qⱓ�RCU� �M�SUXTASK��3NB��0�$TAT�U�P�8�RS�@@쐦F�6�_�PC�}�$FREEF�ROMS]p�ai�GsETN@S�UPDl��ARB�#P%0����� !m$US�A���az9�L�ER1I�0f��pRY�5~"�_�@f�P�1�!�6WRK��D9�F9�~�FRIEND�Q�4bUF��&�A@TO�OLHFMY5�$�LENGTH_VT��FIR�pqC�@��E� IUFINt�R���RGI�1��AITI:�xGX���I�FG2�7G1`a����3�B�GPRR�DA��O_� o0e�I1�RER�đ�3&���T�C���AQJV �G(|�.2���F��1�! d�9Z�8+5K�+5��E��y�L0�4�X T�0m�LN�T�3Hz���89��%�4�3G��W$�0�W�RdD�Z���Tܳ��K�a3d��=$cV 2���1���I1H�02K2
sk3K3Jci�aI��i�a�L��SL��R$)Vؠ�BV�EVk�]V*R��� �,6Lc����9V2F{/P:B��P5S_�E��$rr�C��ѳ$A0��wP!R���v�U�cSk�� �{�X�6��� 0����VX`�!�tX`���0P�Ё�
�5S^K!� �-qR���!0���z�NJ A)X�!h�A�@LlA��^A�THIC�1��8�����1TFE���q>>�IF_CH�3A�aI0�����G1�x�������9�Ɇ_�JF҇PR(����RVAT�� ��-p��7@����DO��E��COU(��A�XIg��OFFS=E+�TRIG�SK���c���Ѽ�e�[�K�Hxk���8�IGMAo0�A-��ҙ�ORG�_UNEV��� ��S�쐮d ӎ$������GR3OU��ݓTO2��!�ݓDSP��JOG�'��#	�_P'�2O�R���>P6KEPFl�IR�0�PM�R&Q�AP�Q��E�0q�e���SYSG��"��;PG��BRK*Rd�r�3�-�������ߒ�<pAD�ݓJ�BS�OC� N�DU�MMY14�p\@S}V�PDE_OP3�SFSPD_OVR��ٰCO��"��OR-��N�0.�F�r�.��OV�SFc�2�f��F��!4��S��RA�"LCHD}L�RECOV��0�W�@M�յ�#RO3��_�0�� @�ҹ@VER�E�$OFS�@CV� 0BWDG�ѴC���2j�
�TR�!|��E_FDOj��MB_CM��U�B �BL=r0�w�=q�t�VfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�#�8$CA�{Й�>��8$HBK|1c��IO��.�:!aPPA"�N�3�^�F����:"�DVC_DB�C��d�w"����!"��1���ç�3����/ATIO� �q0��UC�&CAB �BS�PⳍP�Ȗ���_0c�SUBCPUq��S�Pa a� ��}0�Sb��c��r"ơ?$HW_C����:c��IcA�A-�l$�UNIT��l��A�TN�f����CYC=LųNECA��[��FLTR_2_F�I���(��}&��LPx&�����_SCT@SF_��F����G����FS|!�¹�CHA�A/����2��RS�D�x"ѡb�r�: _T��PRO��O�� KEM�_��8u�q u�q��D�I�0e�RAILAiC��}RMƐLOԠdC��:anq��wq��V��PR��SLQ�p�fC��30	��FUsNCŢ�rRINkP`+a�0 ��!RA� >R 
Я�ԯgWAR�BLFQ���A�����D�A�����LD@m0�aB9��nqBTIvrbؑ���PgRIAQ1�"AFS�P�!�����`%b����M�I1U�D�F_j@��y1°LM�E�FA�@HRDY4�4��Pn@RS@Q�0|"�MULSEj@xf�b�q �X���ȑ���$.A-$�1$c1Ó����� x~�EaG�0ݓ�q!AR����09>B�%��wAXE��ROB���W�A4�_�-֣SYЯ��!6��&S�'WR䩐�-1���STR���5�9�E�� !	5B��=QB90��@6������OT�0vo 	$�ARY8��w20���	%�FI���;�$LINK(�H��1�a_63��5�q�2XYZ@"��;�q�3@��1�2J�8{0B�{D0��� CFI��6G`��
�{�_J�p�6��3aOP_O42Y;5�QTBmA"2�BC
�z�DU"�6=6CTURN3�vr��E�1�9�ҍGFL��`���~ �@�5<:7��� 1�?0K�Mc�68Cb�vrb�4�ORQ��X� >8�#op������wq�Upf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W���T υ� ;����QH�!` �ҽ��U�Q�WkeK#keLcXER��	G!E	0��S�dAWaǢ�:D���7!�!AX�rB!{q��1u y-!y�pz�@z �@z6Pz\Pz� z 1v�y�y�+y �;y�Ky�[y�ky��{y��y�q�yDEBU��$�����L�!º2WG`  AB�!�,��SV���� 
w���m���w��� �1���1���A���A�� 6Q��\Q���!�m@�\�2CLAB3B�U������S  �ÐER���� �� $�@� Aؑ!p�PO��Z�q0w��^�_MRAȑ� �d  T�-�EcRR��TYz��B�I�V3@�cΑTOQ�d:`L� �d2��R]�X�C[! � p�`T}0i��_V1�r�a'�4��2-�2<����@P�8����F�$W��g�j�V_!�l�$�P�����c��q"�	��SFZN_CFG_!� 4��?º��|�ų����@�ȲW q����\$� �n����Ѵ��9c�Q��(�F�A�He�,�XED@M�(�����!s�Q��g�P{RV HELL�ĥ� 56�B�_BAS!�RSR(��ԣo �#S��[���1r�%��2ݺ3�ݺ4ݺ5ݺ6ݺ7rݺ8ݷ��ROOI�䰝0�0NLK!�CAqB� ��ACK��IN��T:�1�@�@� z�m�_PU!�CYO� ��OU��P� �Ҧ) ��޶��TPFWD_KARӑL��RE~��P��(��QUE�����P�
��CSTOPI_AL�����0&��8�㰑�0SEMl�bԲ|�M��d�TY|�SOK�}�DI����꣸(���_TM\�MOANRQ�ֿ0E+��|�$KEYSWITCH&	���{HE
�BEAT����E� LEҒ���U��FO�����O�_HOM�O�REF�PPRz��!�&0��C+�OA�E�CO��B�rIOcCM�D8׵�]�8��8�` � D�1����U��&�MH�»P��CFORC��� ���OM�  G� @V��|�U,3EP� 1-�`� 3-��4�p �SNPXw_ASǢ� 0Ȱ�ADD����$S�IZ��$VAR\ݷ TIP]�\�
2�A򻡐���]�H_� �"S꣩!Cΐ���FRIF⢞�S0�"�c���NF��V ܻ�` � x�`SI��TES�R6SSG%L(T�2P&��AxU�� ) STMTQ2ZPm 6BW�P*�SHOWb��S�V�\$�� ���A00P�a�6���@�J�T�5��	6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	 f0u�	�0u�	�@uP[Pu%121?U1L1Y1f1sU2�	2�	2�	2�	U2�	2�	2�	2U22%222?U2L2Y2f2sU3P)3�	3�	3�	U3�	3�	3�	3U33%323?U3L3Y3f3sU4P)4�	4�	4�	U4�	4�	4�	4U44%424?U4L4Y4f4sU5P)5�	5�	5�	U5�	5�	5�	5U55%525?U5L5Y5f5sU6P)6�	6�	6�	U6�	6�	6�	6U66%626?U6L6Y6f6sU7P)7�	7�	7�	U7�	7�	7�	7U77%727?U7,i7Y7Fi7s��'��VP�UP}D��  ��x|�԰��YSLOǢ� � z��и� ��o�E��`>�^t��А�ALUץ����CU����wFOqID_L��ӿuHI�zI�$FILE_���t�ĳ$`�JvSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_ �TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅�%L~�_Vj��+p�ޠ�� ` �GR�OU�pD��B�N�FLIC��RE�QUIREa�EB�UA��p����2��������c��{ \��APPR��iC���
�EN��CLOe��S_M� v�,ɣ�
���7� ���MC�&����g�_MG�q�C�� �{�9���|�BRKz�NOL��|ĉ R��_LI|��Ǫ�k�J����P
���ڣ������&���/���6��6��8������� ��8�%��W�2�e�PATH a�z�p�z�=�vӥ�ϰm�x�CN=�CA������p�IN�UCh��bq��CO�UM��!YZ������qE%����2������PAYL�OA��J2L3pR'_AN��<�L��F��B�6�R�{�R_F2�LSHR��|�LO�G��р��ӎ���ACRL_u�������.�r��H�p�$H{�^��FLEX
�s�}J�� :� /����6�2�����;�M�_�F16����n�@��������ȟ��Eҟ �����,�>�P�b� ��d�{�������������5�T��X ��v���EťmF ѯ�������&��/�A�S�e�D�Jx�� � ������j��4pAT����n�EL�  �%øJ���vʰJE��CTR�і��TN��F&��H�AND_VB[�
�pK�� $Fa2{�6� �rSW$#��U��� $$	Mt�h�R��08��@<b 35��^6A�p3�kƈ�q{9t�A�̈p��A���A�ˆ0��U���D*��D��P��G��ICST��$A��$AN��DYˀ�{�g4�5D� ��v�6�v��5缧�^�@��P����ՠ#�,�5�>�r�J�� &0�_�ER!V9��SQASYM��] ������x��ݑ���_SHl�������sT�( ����(�:�JA����S�cir��_VI��#Oh9�``V_UCNI��td�~�J�� �b�E�b��d��d�f ��n���������uNI���D��H��f����"CqEN� &a�DI��>�Obt2�Dpx�� ��2IxQA����q��-��s� �� ����� �^�OMME�h�rr/�TVpPT�P  ���qe�i����P��x ��yT�Pj� �$DUMMY9��$PS_��R�Fq�0$:� ����!~q� XX����K�STs�ʰ�SBR��M21_�Vt�8$SV_E�Rt�O��z���CLRx�A  O�r?p? �Oր � D ?$GLOB���#LO��Յ$�o���P�!SYSADqR�!?p�pTCHM0 � ,����oW_NA��/��e���r�SR��l (:]8:m� K6�^2m�i7m�w9m� �9���ǳ��ǳ���ŕ ߝ�9ŕ���i�L� ��m��_�_�_�TDџXSCRE�ƀӚ� ��STF����}�pТ6�1] _:v AŁ� T����TYP�r�K��u�!u���O�@I�S�!��tHD�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J��*��SE=�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� D�C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!&; SHI9F��|s�P�p��6�s���R���OS�URW�pRADIz��2�_�q�h�`g! �q)�LUza�$OUTPUTg_BM��IML��oR6(`)�@TILN<SCO�@Ce� ;��9��F��T�� a��o�>�3���$��w�2u�b�V�zu9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+Z�t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2� �2���5��`�? �PZA�BCS��  �$�2��J�
  �$$CLAS�����A��@<'@@VIRT��O�.@ABS�$�1 �<E� ?< *AtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d��v�����M@[�AXL�ր�&A�dC  �Ʃ�IN��ā��PR�E�����L�ARMRECOV� <I䂥�NG��� \K	 =�#�
J�\�M@PP7LIC�?<E��E�Han�dlingToo�l �� 
V7�.50P/28 �*A�b��
��_SW�� UPn*A� ��F0ڑ䢒��A@��� 20��*A����:����mFB 7DA5��� �'@	b�@����None엃���� ���Tg}*A4�`�x��P_��V�����g�UTO�B�ค����HGA�PON8@��LA��Uޖ�D 1<EfA���������^� Q 1שI Ԁ��Ԑ�:�i�pn����#B)B� ���\�H�E�Z�r�HTTHKY��$BI�[�m�� ���	�c�-�?�Q�o� uχϙϫϽ������� �_�)�;�M�k�q߃� �ߧ߹��������[� %�7�I�g�m���� ����������W�!�3� E�c�i�{��������� ������S/A_ ew������ �O+=[as �������K/ /'/9/W/]/o/�/�/ �/�/�/�/�/G??#? 5?S?Y?k?}?�?�?�? �?�?�?COOO1OOO UOgOyO�O�O�O�O�O �O?_	__-_K_Q_���(�TO4�s���DO?_CLEAN��e���SNM  9� �9oKo]ooo�o��DSPDRYRL�_%�HI��m@&o �o�o#5GYk }����"���p�FՆ �ǣ�qXՄ�ߢ��g�PLUG�GҠ�Wߣ��PRC*�`B`9��o��=�OB��oe�SEGF��K������o%o�����#�5�m���LAP�oݎ�������� ��џ�����+�=��O�a���TOTAL��.���USENU
ʀ׫ �X���R(��RG_STRIN�G 1��
��M��Sc�
~��_ITEM1 �  nc��.�@�R� d�v���������п� ����*�<�N�`�r��I/O SI�GNAL��T�ryout Mo{de�Inp���Simulate�d�Out���OVERR�` �= 100�I?n cycl����Prog Ab�or�����St�atus�	Heartbeat���MH Faul<B�K�AlerUم� s߅ߗߩ߻��������� �S���Q ��f�x������ ��������,�>�P��b�t�������,�WOR������V��
 .@Rdv��� ����*<N`PO��6ц ��o�����/ /'/9/K/]/o/�/�/��/�/�/�/�/�/�DEV�*0�?Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O|�O�OPALTB� �A���O�O__,_>_ P_b_t_�_�_�_�_�_��_�_oo(o:o�OGRI�p��ra�OLo�o �o�o�o�o�o* <N`r������`o��RB���o �>�P�b�t������� ��Ώ�����(�:��L�^�p����PREG�N��.������� �*�<�N�`�r����� ����̯ޯ���&�~���$ARG_���D ?	����i�� � 	$��	[}�]}���Ǟ�\��SBN_CONF�IG i��������CII_S�AVE  ���۱Ҳ\�TCELL�SETUP �i�%HOME_�IO�͈�%MO�V_�2�8�REP����V�UTOBA�CK
�ƽ�FRA:\��c �Ϩ���'`!���������� ����$�6�c�Z�l����Ĉ�������� �����!凞��M�_� q����2������� ��%�7���[�m�� ������@�������0!3E$���Jo��������INUI�@��ε��?MESSAG�����q��ODE_D$���O,0.��oPAUS�!�i�? ((Ol�� ������ /� //$/Z/H/~/l/�/��'akTSK  �q�����UPD�T%�d0;W_SM_CF°i��еU�'1GRP� 2h�93 |�B���A�/S�XSCR�D+11
1; ����/�?�?�? O O$O��߳?lO~O�O �O�O�O1O�OUO_ _ 2_D_V_h_�O	_X���GROUN0O�S_UP_NAL�h�s	�ĠV_ED� �11;
 �%�-BCKEDT-`�_`�!oEo%���Pa��o����������e2no_˔o�o�b���ee�o"�o�oED3�o�o� ~[�5GED4 �n#�� ~�j���ED5Z��Ǐ6�� ~���}���ED6 ����k�ڏ ~G���!�3�ED7��Z��~�� ~�V�şןED80F�&o��Ů}��8��i�{�ED9ꯢ�W�Ư
}3�����CRo�����3�տ�@ϯ����P�PNO_�DEL�_�RGE_�UNUSE�_�TL�AL_OUT �q�c�QWD_A�BOR� �΢Q��I�TR_RTN�����NONSe����CAM_PA?RAM 1�U3�
 8
SON�Y XC-56 �23456789�0�H � @����?���( �АV�|[r؀:~�X�HR5k�|U8�Q�߿�R57�����Aff��KO�WA SC310�M|[r�̀�d @6�|V��_� Xϸ���V��� ���$��6��Z�l��CE__RIA_I8557�F�1��R�|]��_LIO4�W=� ��P<~�F�<�GP 1�,���_GYk*�C*  ��C1*� 9� @� G� ЭCLC]� d� l�� s�R� ��[��m� v� � ��� �� C�� �b"�|W��7�HEӰ�ONFI� ��<G_PRI 1�+P�m®/���������'CHKPwAUS�  1E� ,�>/P/:/t/ ^/�/�/�/�/�/�/�/ ?(??L?6?\?�?"�O�����H�1_�MOR�� �>�PBZ?����5 	 �9 O�?$O@OHOZK�2	���=$9"�Q?55��C�P)K�D3P������a�-4�O__|Z
�OG_�7�PO��� ��6_��,xV�AD�B���='�)
m�c:cpmidb�g�_`��S:�)�����Yp�_)o�S`	�BBi�P�_mo8j�)�Koo�o9i+�)��og�o�o
�m�of�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`)ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCPU�eB��CF��;.<C����C5rSZE@D��nyDQ��D���>��D�;D�����F��>F�$�G}RB�7Gzր��SY��)!�vqG���Em�U)�.��)�)�1�<�q�G�x2��eҢ �� a�D�j��E�e��EX��EQ�EJP �F�E�F� �G�ǎ^F �E�� FB� �H,- Ge���H3Y���  �>�33 ����xV  n2xQ@F��5Y��8B� A�A�ST<#�
� ��_'�%��wRSMO�FS���~2�yT}1�0DE �O� c
�(�;�"� � <�6�z�R��X�?�j�C4��SZ�m� W��{�m�CR��B-G�C�`@$��q��T{�FPROG %i�����c�I��� �Ɯ�f�K�EY_TBL  �vM�u� �	
��� !"#�$%&'()*+�,-./01c�:�;<=>?@AB�C�pGHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������p����͓���������������������������������耇��������������������!j�LCK��.�j����STAT���_A�UTO_DO����W/�INDT_ENB߿2R��9�+��T2w�XSTOP�\߿2TRLl�LE�TE����_SCREEN i�kcsc��U���MMENU 1� i  < g\��L�SU+�U��p3 g������������ 2�	��A�z�Q�c��� ������������. d;M�q�� ����N% 7]�m��� /��/J/!/3/�/ W/i/�/�/�/�/�/�/ �/4???j?A?S?y? �?�?�?�?�?�?O�? O-OfO=OOO�OsO�O �O�O�O�O_�O_P_�Sy�_MANUAyL��n�DBCOU��RIG���DBN�UM�p��<���
��QPXWORK 1!R�ү�_oO�.o@oRk�Q_AWA�Y�S��GCP r��=��df_AL�P�db�RY�������X�_�p 1"�� , 
�^���o �xvf`MT�I^�rl@|�:sONTIM�כ����Zv�i
�õ�cMOTNEN�D���dRECOR/D 1(R�a��ua�O��q��sb �.�@�R��xZ���� ���ɏۏ폄���#� ��G���k�}�����<� ş4��X���1�C� ��g�֟��������ӯ �T�	�x�-���Q�c� u����������>�� ��)Ϙ�Mϼ�F�� �ϧϹ���:������� %�s`Pn&�]�o��ϓ� ~ߌ���8�J����� 5� ��k����ߡ�� J�����X��|��C� U����������0������	��dbTOL�ERENCqdB�ܺb`L�͐PCS_CFG )�k�)wdMC:\�O L%04d.C�SV
�pc�)sA� �CH� z�p�)~���hMRC_OUT *�[��`+P SGN �+�e�r��#��10-MAY-20 10:38*V�27-JANj2�1:4rv P;���)~��`pa�m���PJPѬV�ERSION �SV2.0�.�6tEFLOG�IC 1,�[ 	DX�P7)�PF.�"PROG_ENqB�o�rj ULSew� �T�"_WRS�TJNEp�V�r`dE�MO_OPT_S�L ?	�es
 	R575)s 7)�/??*?<?'�$TO  �-��?�&V_@pEX�Wd��u�3PATH ;ASA\�?�?\O/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C���SqqF�PMAqU� t/XrMSWR�.�i6.|S/�Z!D_N�O0__T_�C_x_g_�_�tSBL__FAUL"0�[^3wTDIAU 16M�6p�A1�234567890gFP?BoTo foxo�o�o�o�o�o�o �o,>Pb�SZ�pP�_ ���_ s�� 0`���� �)�;�M�_�q����������ˏݏ��|)U3MP�!� �^��TR�B�#+�=�PM�EfEI�Y_TEM=P9 È�3@�3�A v�UNI�.(Y�N_BRK 2�Y)EMGDI_�STA�%WЕNC�2_SCR 3��1o"�4�F�X�fv ���������#��ޑ14����)�;������ݤ5��� ��x�f	u�ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/߭P�b�t�� �� xߞ߰���������
� �.�@�R�d�v��� �����������*� <�N���r��������� ������&8J \n������ ��"`�FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/4? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O ?�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�O�O�o�o�o
 .@Rdv�� �������*� <�N�`�r����o���� ̏ޏ����&�8�J� \�n���������ȟڟ�����H�ETMO�DE 16���� ��ƨ
�R�d�v�נRROR�_PROG %fA�%�:߽�  ���TABLE  �A������#�L�R�RSEV_NUM�  ��Q���K�S���_AUT�O_ENB  ���I�Ϥ_NOh� �7A�{�R� W *���������	���^�+��Ŀֿ���HISO���I�}�_ALM 18A�� �;�����+�e�wωϛϭϿ�r�_H���  A����|��4�TCP_VER !A��!����$EXTL�OG_REQ�9�{�V�SIZ_�QԿTOL  ��D}z��=#׍�?XT_BWD���иr���n�_DI�� 9��}�z���<m���STEP����|4��OP_DO����ѠFACTO�RY_TUN�d�G�EATURE �:����l��Handlin�gTool �� � - CEn�glish Di�ctionary���ORDEA�A Vis�� M�aster���9�6 H��nalo�g I/O���H�551��uto �Software� Update � ��J��mati�c Backup~��Part&��ground E�dit��  8\�apCame�ra��F��t\j�6R�ell���LwOADR�omm���shq��TI" ��co��
! yo���pane��� 
!��ty�le selec]t��H59��nD�~��onitor��48����tr��R�eliab���a�dinDiagnos"����2��2 ual Che�ck Safet�y UIF lg�\a��hance�d Rob Se�rv q ct\���lUser F�rU��DIF��E�xt. DIO 6��fiA d��wendr Err YL@��IF�r�ನ  �П�90��F�CTN Menu�Z v'��74� T�P In��fac�  SU (�G=�p��k E�xcn g�3��High-Sper wSki+�  sO��H9 � mmuni]c!�onsg�te�ur� ����V��y��conn���2��EN��Inc=rstru����5.fdKA�REL Cmd.� L?uaA� O~�Run-Ti� 'Env����K� ��u+%�s#�S/W���74��Licen�seT�  (A�u* ogBook�(Sy��m)��"�
MACR�Os,V/Off�se��ap��MH�� ����pfa5�M�echStop �Prot��� d��b i�Shif����j545�!x�r ��#��,p�b ode Swiwtch��m\e�!�o4.�& pr�o�4��g��M?ulti-T7G����net.P{os Regi���z�P��t Fu9n���3 Rz1���Numx �����9�m�1�  Adju<j��1 J7�7�*� ����6tatu�q1EIKRD�Mtot��scove�� ��@By<- }uest1�$G�o� � U5\SNPX b"���<YA�"Libr��㈶�#�� �$~@h�p�d]0�Jts i?n VCCM����ĕ0�  �u!��2 �R�0�/I�08~��TMILIB�M� J92�@P�A�cc>�F�97�TgPTX�+�BRSQselZ0�M8 Rm��q%��692��Unexceptr �motnT  CcVV�P���KC�����+-��~K  I�I)�VSP CSXC�&.c�� e�"��� t�@We�w�AD Q�8bv9r nmen�@�KiP� a0y�0��pfGridAplay !� nh�@*��3R�1M-10iA�(B201 �`2�V"  F���sci�i�load��8�3 M��l����G�uar�d J85��0�mP'�L`���s�tuaPat�&]$C�yc���|0ori�_ x%Data'Pqu���ch�1���g`� j� RLJa�m�5���IMI �De-B(\A�cP"� #^0C  e�tkc^0assw�o%q�)650�Ap�U�Xnt��PvKen�CTqH�5�0�YELLOW� BO?Y��� Arc�0vis��C�h�WeldQci�al4Izt�Op�� ��gs�` 2@�a6��poG yRjcT1 NE�#HTf� xyWb��! �p��`gd`���p\� �=P��JPN ARCP*PR�A�� �OL�pSup̂fil�p��J�� n��cro�670�1�C~E�d��SS�pe.�tex�$ �P� �So7 t� ssa%gN5 <Q�BP:� 2�9 "0�QrtQCr��P�l0dpn������rpf�q�e�ppm�ascbin�4psyn�' pstx]08�HEL�NCL VIS �PKGS �Z@M�B &��B J8�@IPE GET_VAR FI?S_ (Uni� LU��OOL: ADD��@29.FD�TC4m���E�@DVp����`A�ТNO WT?WTEST �� ��!��c�FOR ^��ECT �a!� �ALSE ALA�`�CPMO-13�0��� b D: H�ANG FROM�g��2��R709� DRAM AV�AILCHECK�S 549��m�V�PCS SU֐L_IMCHK��P�0~x�FF POS� �F�� q8-12 CHARS��ER6�OGRA ���Z@AVEH�AME��.SV��Вאqn$��9�m "y��TRCv� SHA�DP�UPDAT �k�0��STATI���� MUCH ����TIMQ MOTN-003���@OBOGUI�DE DAUGH໱�b��@$tou�� �@C� �0��PA�TH�_�MOVE�T�� R64��V�MXPACK M�AY ASSERyTjS��CYCL`��TA��BE CO�R 71�1-�AN���RC OPTI�ONS  �`��A�PSH-1�`fi	x��2�SO��B��XO򝡞�_T��	�i�j�0j��du�byz �p wa��y�٠H�I������U�pb X?SPD TB/�F�_ \hchΤB0����END�CE�06�\Q�p{ sma'y n@�pk��L} ��traff#��	� ��~1fro�m sysvar/ scr�0R� ��Nd�DJU���H��!A��/��SET GERR�D�P7�����NDANT S�CREEN UNREA VM �P�D�D��PA���R~�IO JNN�0��FI��B��GRwOUNנD Y��Т٠�h�SVIP� 53 QS��DI�GIT VERS���ká�NEW�� �P06�@C�1IMCAG�ͱ���8� �DI`���pSSU�E�5��EPLAN� JON� DELL���157QאD��CALLI���Q��m���IPND}�IMG N9 PZ�{19��MNT/���ES ���`LocR Hol߀=��2�P�n� PG:��=�M��can����С�: 3D mE2view d X���ea1 �0b�po;f Ǡ"HCɰ��ANNOT AC�CESS M c�pie$Et.Qs �a� loMdFle�x)a:��w$qmo+ G�sA9�-'p~0̿�h0pa��eJ AUTO-�0��!�ipu@Т<ᡠIA�BLE+� 7�a F�PLN: L�p�l m� MD<�V�I�и�WIT H�OC�Jo~1Qu�i��"��N��US�B�@�Pt & r�emov���D�vAxis FT_7�PGɰCP:�O�S-144 � h� s 268QՐO�ST�p  CRA�SH DU��$P~��WORD.$��LOGIN�P��P�:	�0�046 i�ssueE�H�:� Slow st�c�`6�����z��IF�IMPR��SPOT:Wh4����N1STY��0V�MGR�b�N�CA�T��4oRRE�� �� 58�1��:N%�RTU!Pe -M .a�SE:�@pp���$AGpL��m@�all��*0a�OC�B WA���"3 �CNT0 T9DW�roO0alarm8�ˀm0d t�M��"0�2|� o�Z@O�ME<�� ��E%  ;#1-�SRE��M��st}0g   �  5KANJI~5no MNS@��INISITA7LIZ'� E�f�cwe��6@� dr�@� fp "��SC�II L�afai�ls w��SY�STE[�i�� � � Mq�1QGro8�m n�@vA�����&��n�0q��R�WRI OF L|k��� \ref"��
�up� de-r�ela�Qd 03�.�0SSchőb�etwe4�INDo ex ɰTPa�#DO� l� �ɰ�GigE�sope�rabil`p l�,��HcB��@]�lye�Q0cflxz�8Ð���OS {�����v4pfigi GL�A�$�c2�7H� wlap�0ASB� �If��g�2 l\�c�0�/�E�� �EXCE 㰁�P����i�� o0��G�d`]Ц�fq�l lsxt��EFal����#0�i�O�Y�n�CL�OS��SRNq1NT^�F�U��FqKP~�ANIO V7/�¥�1�{����DBa �0��ᴥ�ED��DET|�'� �b�F�NLINEb�B�UG�T���C"RL�IB��A��ABC? JARKY@���� rkey�`IL����PR��N��ITG+AR� D$�R �Er *�T��a�U�0��h�[�ZE V�� TASK p7.vr�P2" .�XfJ�srn�S谥d�IBP	c���B/��BUS��UNN�� j0-�{��cR�'���LOE�DIVS�CULs$cb����BW!��R~�W`�P�����IT(঱t�ʠ�OF��UNE�Xڠ+���p�FtE���SVEMG3`N�ML 505� D�*�CC_SAFE��P*� �ꐺ� PE�T��'P�`�F  �!���IR����c Ri S>� K��K��H GUNCHGz��S�MECH��IM��T*�%p6u���tPORY LE�AK�J���SP�EgD��2V 74\GRI��Q�g��oCTLN��TRe `@�_�p ���EN'�IN������$���r��T3)�i�STO��A�s�L��͐X	���q��Y� ��CTO2�J m��0F<�K����DU�S��O���3 9�J F��&���SSVGN�-1#I���RSRwQDAU�Cޱ� �T6��g��� 3�]���BR�KCTR/"� �q\�j5��_�Q�S�qI{NVJ0D ZO�P ݲ���s��г�Ui ɰx̒�a�DUAL�� J50e�x�RV�O117 AW�T�H!Hr%�N�247�%�52��|�&aol� ���R���at�Sd��cU���P,�LER��iԗQ0�ؖ  S!T���Md�Rǰt�_ \fosB�A�0@Np�c����{�U���ROP 2�b�pB>��ITP4M��b !AUt c0< � �plete�N@�� z1^qR635� (AccuCa�l2kA���I) �"�ǰ�1a\�Ps ��ǐ� bЧ0P������ig\cba?cul "A3p_ �1��ն���eta�ca��AT���PC��`�����_p�.�pc!Ɗ��:�cicrcB���5�tl��Bɵ�:�fm+�Ί��V�b�ɦ�r�upf�rm.����ⴊ�x�ed��Ί�~�ped�A�D �}b�ptl�ibB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆Ϙ���c�Ӳ�5�1j>�����tcȐ�Ϣ	�r����mm 1���T�sl^0��T�m�ѡ�#�rm3��u8b Y�q�std}��3pl;�&�ckv�=߆r�vf�䊰��9�v1i����ul�`�04fp�q �.f���� daq; i Da�ta Acqui+si��n�
��4T`��1�89���22 DMCM oRRS2Z�75���9 3 R710,�o59p5\?T "��1 (D�T� nk@���� ����E Ƒȵ��Ӹ��etdmm ��ER�����gE��1�q\mo?۳�=( G���[(

�2�` �! �@JMAC�RO��Skip/Offse:�a���V�4o9� &qR6C62���s�H��
 6Bq8����9~Z�43 J77� =6�J783�o `��n�"v�R5�IKCBq2 PT�LC�Zg R�3; (�s, �������03�	зJ���\sfmnmc? "MNMC�����ҹ�%mnf�FM�C"Ѻ0ª etm�cr� �8����� ,pD�p   874\prdq>�,jF0���axi�sHProcess Axes e�wrol^PRA
��Dp� 56 J81�j�59� 56o6�� ���0w�690 998� [!IDV�1��2(x2��2ont �0�
����m2����?C��etis "ISD��9�� F/praxRAM�P�8 D��defB�,��G�isbasicHB�@޲{6�� W708�6��(�Acw:������D
�/,��AMOX�� ��DvE ��?;T��>Pi� RACFM';�]�!PAM�V �W�Ee�U�Q'
bU�75�.�ceN�e� nterfa�ce^�1' 5&!5�4�K��b(Dev am±�/�#���/<�Tazne`"DNEWE����btpdnui� �AI�_s2�d_rsono���bAs�fjN��bdv_arFvf�xhpz�}w��shkH9xstc��gAponlGzv{�ff��r���z��3{q'Td>pcOhampr;e�p� ^5977��	܀�4}0��mɁ�/�����l�f�!�pcchmp�]aMP&B�� �m�pev�����p�cs��YeS�� M/acro�OD��16Q!)*�:$�2U"_,x��Y�(PC ���$_;������o��J�g�egemQ@GEM�SW�~ZG�gesn�dy��OD�ndda��S��syT�Kɓ�Csu^Ҋ���n�m��<�L��  ���9:�p'ѳ޲��spotplusp���`P-�W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\f�eatu 0FEA�WD�oolo�s�rn'!2 p���a؝As3��tT.� (?N. A.)��!�e!�J# (j�,`��oBIB�oD -��.�n��k9�"K���u[-�_���p� "PSEqW����?wop "sEЅ� &�:�J������y�|� �O8��5��Rɺ��� ɰ[��X������ـ%�(
ҭ�q HL �0k�
�z�a!�B�Q�"(g�Q����� ]�'�.�����&���<�0!ҝ_�#��tpJ�H� ~Z��j�����y���� ��2��e������Z�� ��V��!%���=�]�p͂��^2�@iRV� Kon�QYq͋JF0B� 8ހ�`�	(^>�dQueue���X�\1�ʖ`�+F1tpv�tsn��N&��ftupJ0v �RDV�	�f��J1 Q���v��en��kvst�k��mp��btk�clrq���get����r��`kack�XZ��strŬ�%�st0l��~Z�np:!�`����q/�ڡ6!l��/Yr�mc�N+v�3�_� ����.�v�/\jF���� �`Q�΋ܒ�N50 (FRA��+�����fraparm���Ҁ�} 6�J6�43p:V�ELSE�
#�VAR $�SGSYSCFG�.$�`_UNITS 2�DG~°@�4�Jgfr��4A�@FRL-��0ͅ�3ې���L �0NE�:�=�?@�8 �v�9~Qx304��;�BPRSM~QA��5TX.$VNUM_OL��5��DJ�507��l� Functʂ"qwAP��琉�3 H�ƞ�kP	9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TP�PR���QA�prnaSV�ZS��AS8D�j510U�-�`cAr�`8 ��ʇ�DJR`�jYȑH  ��Q �PJ6�a2�1��48AA�VM 5�Q�b0 �lB�`TUP xb?J545 `b�`�616���0V�CAM 9�CwLIO b1�s5 ���`MSC8��
rP R`\s�STYL MNI�N�`J628Q  �`NREd�;@�`�SCH ��9pDCSU Mete�`�ORSR Ԃ�a0�4 kREIO�C �a5�`542�b9vpP<�nP�a�`�R�`7�`�M?ASK Ho�.r�7 �2�`OCO :��r3��p�b�p���r0X��a�`13\�mn�a39 HR�M"�q�q��L�CHK�uOPLG� B��a03 �q.��pHCR Ob�pC�pPosi�`fP6� is[rJ554��òpDSW�bM�D8�pqR�a37 }Rjr30 �1�s4 �R6�m7��52�r5 �2.�r7 1� P6����Regi�@T^�uFRDM�uSaq�%�4�`930�uS�NBA�uSHLB�̀\sf"pM�N{PI�SPVC�oJ520��TC�`�"MNрTMIL��IFV�PAC �W�pTPTXp6�.%�TELN N� Me�09m3�UECK�b�`U�FR�`��VCOR^��VIPLpq89q�SXC�S�`VVF��J�TP �q��Rw626l�u S�`�Gސ�2IGU�I�C��PGSt�\ŀH863�S�q������q34sŁ6�84���a�@b>�3� :B��1 T��9�6 .�+E�51 �y�q53�3�b1 ̛��b1 n�jr9 <���`VAT ߲�q�75 s�F��`�sA�WSM��`TOP u�ŀR52p���a�80 
�ށXY �q���0 ,b�`8855�QXрOLp}��"pE࠱tp�`LCyMD��ETSS�挀6 �V�CPEs oZ1�VRCd3�
�NLH�h��0011m2Ep��3 f��p���4 /165CR��6l���7PR���008 tB��9 o-200�`U0�p�F�1޲1 ��޲2 L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�J�?7 rbcfA�L��8\PC����"�32�m0u�n�K�Rٰn�5� 5EW
n�99 z��40 kB���3 ��6ݲ�`00�iB/��6�u��7�u��8 µ������s�U0�`�t �1 0�5\rb��2 E@���K���j���5˰��60��a�HУ`:Ł63�jAF�_���F�7 ڱ݀H�8�eHЋ�&�cU0��7�p���1u��8u��9 c73������D7� r��5t�97 ��E8U�1��2��1�)1:���h��1np�"���8(�U1��\pyl��,࿱v ��B�854��1V���D�-4��im��1�<����>br�3pr�48@pGPr�6 B����$�p��1����1�`͵�155ض157 �2��62�S����B��1b��2����1Π2"�2���B6`�1<c�4 7B�5i DR��8_�B/���187 uJ�8 ;06�90 rBn��1 (��202 /0EW,ѱ2^��2��90�U2�p�2��S2 b��4��2�a�"RB����9\�U�2�`w�l���4 6	0Mp��7������b�,s
5 ��3����<pB"9 3 ����l�`ڰR,:7 �2��V�2��5���2^H��a^9���qr�����n�5����5᥁""�8a�Ɂ}�5B���5����`UA���� ���86 �6 S�0�5�p�2�#�52�9 �2^�b1
P�5~�2`���&P*5��8��5��u�r!�5��ٵ544��%5��R�ąP nB^,z�c (�4���L���U5J�V�5��1�1^��%�����5 b21��gA���58W82� r�b��5N�E�589�0r� 1�95  �"������c8"a��|�L ���!J"5|6���^!��6��B�"8P�`#��+�8%�6B��AME�"1 iCN��622�Bu�6V���d� 4��84�`A�NRSP�e/S� C�5� �6� ��� \� �6� �V� 3�t��� T20CA�R��8� Hf� 1D�H�� AOE� ��� ,|�� a�0\�� �!64K���ԓrA� �1 (M{-7�!/50T� [PM��P�Th:1�C��#Pe� �3�0� 5>`M75T"� �D�8p� �0Gc� u�4|��i1-710i�1B� Skd�7j�?6�:-HS,� �RN�@��UB�f�X�=m7C5sA*A6an���!X/CB�B2.6A �0 ;A�CIB�A�2�QF1�U�B2�21� /70�S� �4����Aj1��3p���r#0 B2\m*A@C��;bi"�i1K�u"A~AAU� imm7c7��ZA@HI�@�Df�A�D5*A��E� 0TkdR1�35�Q1�"*�@�Q�1�QC )P�1*A�5*A�EA�5XB�4>\77
B7=Q �D�2�Q$B�E7�C�D%/qAHEE�W7�_|` jz@� 2�0�Ejc�7�`�E"l7�@7@�A
1�E�V~`�W2%Qr�R9ї@0L_�#�����"A���b��H3s=rA/2�R5nR 4�74rNUQ1ZU�A�sw\m9
1M92L2��!F!^Y�ps� 2c1i��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHsXBSt62�q`s������ ��Pxq3530_*A3I)�2�db�u0�@� '4TX�m0�pa3i1A3s0Q25�c��st�r�VR1%e�q0
��j1 ��O2 �A�UEiy�@.�‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?P Q��qA!Pvs� 5	1 5aU���?PŅ���ဝQ9A6�zS*�7�qb5�1����Q��'00P(��V7]u�a itE1���ïp?7� �!?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ�޵y00\ry�"R�2BL�tN  ���� �1DAp�2�qeR�5���_b�3�X]1m1l�cqP1�a�E�Q� 5�F����!5���@M-16Q�� f���r���Q�e� ��� PN�L�T_�1��i1��945�3��@�e�|�b1l>F1u*AY2�
�R8�Q����RJ�J13�D}T� 85
Qg� /0��*A!P�*A�Ð�d����2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt]1 ^u�ajrI�B����~`�|I�b��yI�\m�Qb�I�uz�A�c3Apa\9q� B6S��S��m���}�85`N�N�  �(M�� �f1���6����161j��5�s`�SC���U��A����5\se�t06c����10��y�h8��a6��6x��9r�2HS �� �Er���W@}�a��IlB���Y�ٖ�m�u �C����5�B��B��h`�F���X0���A :���C�M��AZ��@��4�6i����� e�O�-	���f1��F  �ᱦ�1F�Y	���GT6HL3��U66~`Ȗ��U�dU�9D20Lf0��Qv� ��fjq ��N������0v
� ���i	�	��72l�qQ2������� \�chngmove�.V��d���@2l_arf	�f ~��6������9C��Z���~���kr41@ S���0��V��t�����U�p7nu�qQ%�A]��V�1\"�Qn�BJ�2W� EM!5���)�#:��64��F�e50S �\��0�=�PV�� �e������E������m7shqQSH"U��)��9�!A���(���� �,p�ॲTR11!��,�60e=��4F�����2��	 R-����������@�Ж��4���LS0R�)"�!lOA��Q�X) %!� 16�
U /��2�"2�E�9p���2>X� SA/i��'�
7F�H�@!B�0�� �D���5V��@2cV E��p��T��pt갖��1L~E�#�F�Q��9�E�#De/��RT��59���	�A�EiR���|����9\m20챃20��+�-u�19r4 �`�E1�=`O9`� �1"ae��O�2��_\$W}am41�4�3��/d1c_std ��1)�!�`_T��r~�_ 4\jdg�a �q�PJ%!~`-�r�+�bgB��#c300D�Y�5j�QpQb1�`bq��vB��v25�Up�����qm43�  �Q<W�"PsA��e ����t�i�P�W .��c�FX.�e4�kE14�44�~o6\j4�443sxj��r�j4up�� �\E19�h�PA�T�= :o�APf��coWol!\�2a��2A;_	2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a�:88J9X�l5�m�1a첚��*���(85�&�������P6���R,52&A����,fA9IfI50\u�z�OV
�v��}E�֖J���Y>� 16�r�C�Y��;��1��L ���Aq�&ŦP1��vB�)e�m�����1pĻ �1Dp�27��F�KAREL �Use S��FC�TN��� J970�FA+�� (�Q޵0�p%�)?�Vj9F?(��j�Rtk208 C"Km�6Q�y�j��iæPr�9�s#��v��krcfp�RCF�t3���Q��kcctme�!ME�g����^6�main�dV�� ��ru��kDº��c���o����J�dt��F �»�.vrT�f�����E%�!��\5�FRj73B�K����UER�HJ�O  �J�� (ڳF���F �q�Y�&T��p�F�z��19�tkvBr���V�Bh�9p�E�y�<�k�������;�v���"CT��f����)�
І ��)�V	�6���!� �qFF��1q���=��� ��O�?�$"���$���je���TCP A�ut�r�<520 �H5�J53E19�3��9��96�!8���9��	 �B574V��52�Je�(�� Se%!Y�����u���ma�Pqtool��ԕ������co�nrel�Ftro�l Reliab�le�RmvCU!��H51����� a�551e"�CNRE¹I�c�&���it�l\sfut?st "UTա��"X�\u��g@�i�D6Q]V0�B,Eѝ6A� �Q�)C���X���Yf�I�1|6s@6i��T6IU��vR��d�
$e%1��2�C58�E6��8�Pv�iV�4OFH58SOeJ� mnvBM6E~O58�I �0�E�#+@�&�F�0 ���F�P6a���)/++��</N)0\tr1x�����P ,pɶ��rmaski�ms�k�aA���ky'd�h�	A	�P�sDisp_layIm�`v��~��J887 ("A��+Heůצprd�s��Iϩǅ�h�0p�l�2�R2��:�Gt�@��PRD�TɈ�r��C�@Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��Px^@�P�firmQ� ���Pp�2�=bk�6�r��3��6��tppl��PL���O�p<b�ac�q	��g1J�U�d0�J��gait_9e���Y�&��Q���	�S�hap��erat�ion�0��R6�7451j9(`sGen�ms�42-f�Ár�p�5����2�rsgl�E��p�G���qF�205p�5S���ՁN�retsap�BP�O��\s� "GC�R�ö? �qngda�G��V��st2axU��Aa]��b�ad�_�btpu�tl/�&�e���tp�libB_��=�2.p����5���cird��v�slp��x�hex��v�re?�Ɵx�gkey�v�pm���x�us$�6�gcr��F������[�q27�j92�v�ollismqSk�9O��>�� (pl.���t��p!o��29$Fo8���cg7no@�tptwcls` CLS�o�b�\�km�ai_
�!s>�v�o	�t�b��x�ӿ�E�H��6~�1enu501�[�m��utia|$c�almaUR��Ca�lMateT;R5	1%�i=1]@-��/V�� ��Z�� �fq1�9 "K9E�L����z2m�CLMTq��S#��et �LM�3!} �F�c�ns�pQ�c���c_mo4q��� ��c_e���F��su��ޏ �_ �x@�5�G�join�@i�j��oX���&cW0v	 ���N�ve��C�clm�&Ao# �|$�finde�0�STD ter� FiLANiG���R��
��8n3��z0Cen���r,������J��� �� ���K��Ú�=�К�_Ӛ��r� "FNDR�� 3��}f��tguid��`��N�."��J�tq��  �������������J����_������c���	m�Z��\fndr.��n#>
B2�p��Z�CP Ma�����38A��� c
��6� (���N�B ������� 2�$�	81��m_���"ex�z5�.Ӛ��c���bSа�ef�Q��	��RBT~;�OPTN � +#Q�*$�r*$��*$r *$%/s#C�d/.,P�/|0*ʲDPN���$���$*�Gr�$ko Exc�'IF�$�MASK�%93 {H5�%H558�$_548 H�$4-1��$��#1(�$�0 E�$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3��9j0"M�49�4 � ��4�4tp�sh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E�\���5�A�4��3a�dq\�5K979�":E�ajO l "�DQ^E^�3i�Dq� ��4ҲO ?R�? ��q�5��T��3rAq�O�Lst�5~��7�p�5��REJ#�2�@a�v^Eͱ�F���4��.��5y N� �2il�(in�4��31 aJH1�2Q4�251ݠ��4rmal� �3) �REo�Z_�æOx�����4��^F�?onor Tf��7_ja�UZҒ4l��5rmsAU�Kkg���4�$HCd\�fͲ�e�ڱ�4�REM���4y�ݱ"u@�RER593�2fO��47Z��5lity,�U��e"DGil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe�=$��^�
E��u�IAymptm�U��BU��vste�y\�3��me� b�DvI�[�Qu�:F�U�b�*_�
E,�su$��_ Er��oxx���4huse�E-�?�sn�������FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��� b���(��1�� �c��Y�R�� �>�P� ��W��������'��0ɵ�[��͂����  � ,N@� �A��bumpšf��B*�Box%��7Aǰ�60�BBw���MC� u(6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`���)���\bbk968� "�4�ω�bb��9va69����etbŠ��X�����#ed	�F��u�f�& �sea"������'�\��,���b�ѽ"�o6�H�
�x�$�f���!y���Q[�!� tperr�f�d� TPl0o� R/ecov,��3D���R642 � 0���C@}s� N@��(NU�rro���yu2�r��  �
�  ����$$�CLe� �������������$~z�_DIGIT��.������ .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ oo$j��+c:PRODUCTM��0\PGSTKD��V&ohozf99���D���$F�EAT_INDE�X��xd���  
�`IL�ECOMP ;����#��`�cS�ETUP2 <��e�b�  �N �a�c_AP2�BCK 1=�i  �)wh0?{%&c����Q� xe%�I�m�� �8��\�n����!� ��ȏW��{��"��� F�Տj���w���/�ğ S���������B�T� �x������=�үa� �����,���P�߯t� �����9�ο�o�� ��(�:�ɿ^���� �ϸ�G���k� �ߡ� 6���Z�l��ϐ�ߴ� ��U���y����D� ��h��ߌ��-���Q� ��������@�R��� v����)�����_��� ��*��N��r� �7��m�@&�3\�i
pP� 2#p*.V1Rc�*��`� /��PC/|1/FR6:/"].��/+T�`�/ �/F%�/�,�`r/?��*.F�8?	�H#&?e<�/�?;STM �2�?�.K �?��=iPen�dant Panel�?;H�?@O�7�.O�?y?�O:GIF �O�O�5�OoO�O_:JPG _J_�56_�O�_�_�	PANE�L1.DT�_@�0�_�_�?O�_2�_�So�WAo�_o�o�Z3 qo�o�W�o�o�o)�Z4�o[�WI���
TPEINSO.XML��0�\���qCust�om Toolb�ar	��PAS�SWORDy�FRS:\L�� �%Passwo�rd Config���֏e�Ϗ�B 0���T�f�������� ��O��s������>� ͟b��[���'���K� �򯁯���:�L�ۯ p�����#�5�ʿY�� }��$ϳ�H�׿l�~� Ϣ�1�����g��ϋ�  ߯���V���z�	�s� ��?���c���
��.� ��R�d��߈���;� M���q������<��� `������%���I��� �����8����n ���!��W�{ "�F�j| �/�Se��/ �/T/�x//�/�/ =/�/a/�/?�/,?�/ P?�/�/�??�?9?�? �?o?O�?(O:O�?^O �?�O�O#O�OGO�OkO }O_�O6_�O/_l_�O �__�_�_U_�_y_o  o�_Do�_ho�_	o�o -o�oQo�o�o�o�o @R�ov��; �_���*��N� �G������7�̏ޏ m����&�8�Ǐ\�� ���!���E�ڟi�ӟ ���4�ßX�j����� ���įS��w�������B�#��$FIL�E_DGBCK �1=��/���� ( ��)
SUMMA�RY.DGL����MD:������Diag Sum�mary��Ϊ
C?ONSLOG������D�ӱCon�sole log�E�ͫ��MEMCHECK:�!ϯ����X�Memory� Data��ѧ��{)��HAD�OW�ϣϵ�J����Shadow C?hangesM�'��-��)	FTAP7Ϥ�3ߨ���Z��mment TB�D��ѧ0=4)�ETHERNET��������T�ӱE�thernet �\�figurat�ionU�ؠ��DCSVRF�߽߫������%�� ve�rify all���'�1PY���DIFF�����[����%��diff]������1R�9�K���� ���X=��CHGD������c��r�����2ZAS� ��GD����k��z��FY�3bI[� �/"GD����s/����/*&UPDATES.� ��/��FRS:\��/�-ԱUpda�tes List��/��PSRBWLOD.CM(?���"�<?�/Y�PS_ROBOWEL��̯�? �?��?&�O-O�?QO �?uOOnO�O:O�O^O �O_�O)_�OM___�O �__�_�_H_�_l_o �_�_7o�_[o�_lo�o  o�oDo�o�ozo�o 3E�oi�o�� �R�v���A� �e�w����*���я `���������O�ޏ s������8�͟\�� ���'���K�]�쟁� ���4���ۯj����� �5�įY��}���� ��B�׿�x�Ϝ�1� ��*�g�����Ϝ��� P���t�	�ߪ�?��� c�u�ߙ�(߽�L߶� �߂���(�M���q�  ���6���Z���� ��%���I���B������2�����h�����$FILE_� P�R� ��������M�DONLY 1=�.�� 
 � ��q��������� �~%�I�m �2��h� �!/�./W/�{/
/ �/�/@/�/d/�/?�/ /?�/S?e?�/�??�? <?�?�?r?O�?+O=O �?aO�?�O�O&O�OJO �O�O�O_�O9_�OF_�o_
VISBCK�L6[*.VD�v_�_.PFR:\��_�^.PVis�ion VD file�_�O4oFo\_ joT_�oo�o�oSo�o wo�oB�of�o �+����� ��+�P��t���� ��9�Ώ]�򏁏��(� ��L�^�������5� ��ܟk� ���$�6�ş�Z��~�����
M�R_GRP 1>�.L��C4 w B���	 W������*u����RHB ���2 ��� ��� ���B� ����Z�l���C���D�ি����Ŀ��J�8�LJ�4�F�5U��R��
���ֿ �Gn�E��.�E88�-���?:u�{@ �����@A�A�!��f�?h!A��%r��E�� F�@ ������ھ���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6\b��+�&�(�a�hL߅�p�A��A��� ��v���r������
� C�.�@�y�d����� ����������?�Z��lϖ�BH�� ��Ζ�������
0�PJ��P�T���ܿ� �B���/ ��O@�33:��.�\gN�UUU�U���q	>u.�?!rX��	�-�=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!��7�:����D��@ D�� CYϥ��C������'/0-��P/����/ N��/r��/���/�? ?;?&?_?J?\?�?�? �?�?�?�?O�?O7O "O[OFOOjO�O�O�O �O�гߵ��O$_�OH_ 3_l_W_�_{_�_�_�_ �_�_o�_2ooVoho So�owo�o�i��o�o �o��);�o_J �j������ �%��5�[�F��j� ����Ǐ���֏�!� �E�0�i�{�B/��f/ �/�/�/���/��/A� \�e�P���t������� �ί��+��O�:� s�^�p�����Ϳ��� ܿ� ��OH��o�
� ��~ϷϢ�������� ��5� �Y�D�}�hߍ� �ߞ��������o�1� C�U�y��߉��� ���������-��Q� <�u�`����������� ����;&_J \���������� ڟ�F�j4�� �������!/ /1/W/B/{/f/�/�/ �/�/�/�/�/??A? ,?e?,φ?P�q?�?�? �?�?O�?+OOOO:O LO�OpO�O�O�O�O�O �O_'__K_�o_�_ �_�_l��_0_�_�_�_ #o
oGo.okoVoho�o �o�o�o�o�o�o C.gR�v�� ���	���<� `�*<��`���� �ޏ��)��M�8�q� \�������˟���ڟ ���7�"�[�F�X��� |���|?֯�?����� 3��W�B�{�f����� ÿ���������A� ,�e�P�uϛ�b_���� �Ϫ_��߀�=�(�a� s�Zߗ�~߻ߦ����� ��� �9�$�]�H�� l������������ #��G�Y� �B����� ��z�������
ԏ:� C.gRd��� ���	�?* cN�r���� �/̯&/�M/�q/ \/�/�/�/�/�/�/�/ ?�/7?"?4?m?X?�? |?�?�?�?�?��O!O 3O��WOiO�?�OxO�O �O�O�O�O_�O/__ S_>_P_�_t_�_�_�_ �_�_�_o+ooOo:o so^o�o�op��o��  ��$��o�o �~������ �5� �Y�D�}�h��� ����׏����
� C�.�/v�<���8��� ���П����?�*� c�N���r�������� ̯��)��?9�_�q� ��JO�����ݿȿ� �%�7��[�F��j� �ώ��ϲ�������!� �E�0�i�T�yߟߊ� �߮��߮o�o��o>� t�>��b���� �������+��O�:� L���p����������� ��'K6oZ �Z�|�~���� �5 YDi�z ������/
/ /U/@/y/@��/�/�/ �/���/^/???Q? 8?u?\?�?�?�?�?�? �?�?OO;O&O8OqO \O�O�O�O�O�O�O�O�_�O7_��$FN�O ����VQ�
�F0fQ kP FL�AG8�(LRRM�_CHKTYP � WP��^P��WP�{QOM�P_�MIN�P�����P�  XNPS�SB_CFG �?VU ��_���S ooIU�TP_DEF_O/W  ��R&h�IRCOM�P8o��$GENOVRD7_DO�V�6�fl�THR�V d�ed�kd_ENBWo �k`RAVC_GR�P 1@�WCa X"_�o_1U <y�r���� �	��-��=�c�J� ��n��������ȏ� ���;�"�_�F�X���.ibROU�`FVX�P�&�<b&�8�?��埘��������  Da?�јs���@@g�B�7�p�)�ԙ���`WSMT�cG�mM����� �LQHOST�C�R1H���PĹ�at�SM���f�\���	1�27.0��1��  e��ٿ���� �ǿ@�R�d�vϙ�0��*�	anonymous���������F��s[�� � �����r����ߨߺ� ����-���&�8�[� I�π����� �1�C��W�y���`� r������ߺ������� %�c�u�J\n� ��������M� "4FX��i�� ����7//0/ B/T/���m/��/ �/�/??,?�/P? b?t?�?�/�?��?�? �?OOe/w/�/�/�? �O�/�O�O�O�O�O=? _$_6_H_kOY_�?�_ �_�_�_�_'O9OKO]O __Do�Ohozo�o�o�o �O�o�o�o
?o}_ Rdv���_�_o o!�Uo*�<�N�`� r��o������̏ޏ� ?Q&�8�J�\���>��ENT 1I��� P!􏪟  ����՟ğ����� ��A��M�(�v���^� ����㯦��ʯ+��  �a�$���H���l�Ϳ �����ƿ'��K�� o�2�hϥϔ��ό��� ��������F�k�.� ��R߳�v��ߚ��߾߀��1���U��y�<�?QUICC0��b�t����1�����%��2&���u�!?ROUTERv�R��d���!PCJO�G����!19�2.168.0.�10��w�NAME� !��!RO�BOTp�S_C�FG 1H�� ��Aut�o-starte�d�tFTP� ������  2D��hz��� �U��
//./A�#����~/�� ��/�/�/�/� ?2? D?V?h?�/?�?�?�? �?�?�?���@O? dO�/�O�O�O�O�?�O �O__*_MON_�Or_ �_�_�_�_	OO-O�_ A_&ouOJo\ono�o�o =o�o�o�o�oo�o 4FXj|�_�_�_ o�7o��0�B� T�#x���������� e�����,�>��� ��ŏ���Ο��� ���:�L�^�p��� ��'���ʯܯ� �O� a�s�����l������� ��ƿؿ����� �2� D�g��zόϞϰ��� �#�5�G�I��}�R� d�v߈ߚ�iϾ����� ���)߫�<�N�`�r����XST_ERR� J5
���PDUSIZ  ��^J����>��W�RD ?t���  guest}��%�7�I��[�m�$SCDMN�GRP 2Kt;�������V$�K�� 	P01.14 8���   y�����B    �;����� ��������
 �������������~����C�.gR|��� � i  � � 
��������� +��������
���l .Vr���"�l��� m
d�������_GROU��L.�� �	�����07EQUPD � 	պ�J�T�Ya ����TT�P_AUTH 1�M�� <!i?Pendany���6�Y!KAREL:*��
-�KC///A/ �VISION SCETT�/v/�" �/�/�/#�/�/
??�Q?(?:?�?^?p>�C?TRL N�����5�
�FF�F9E3�?�F�RS:DEFAU�LT�<FAN�UC Web S_erver�:
� ����<kO}O�O�O�O��O��WR_CON�FIG O�� ��?��IDL_�CPU_PC@��B��7P�BH�UMIN(\��<TGNR_IO��������PNPT_SI�M_DOmVw[T�PMODNTOL�mV �]_PRTY��X7RTOLNK 1P����_o!o�3oEoWoio�RMAS�TElP��R�O_gCFG�o�iUO�|�o�bCYCLE�o��d@_ASG 19Q����
 ko, >Pbt����������sk�bN�UM����K@�`I�PCH�o��`RTRY_CN@oR���bSCRN����Q���� �b�`�bR���Տ��$J2�3_DSP_EN�	����OBP�ROC�U�iJO�GP1SY@��8�?�!�T�!�}?*�POSRE�~zVKANJI_�` ��o_�� ��T�L�6�͕����CL_L�GP<�_���EYLO�GGIN�`����LANGUA�GE YF7R�D w���LG��U��?⧈�x� ������=P��'0���$ NMC�:\RSCH\0�0\��LN_DISP V��
�ј������OC�R.RD�zVT=#�K@9�B?OOK W
{��`i��ii��X������ǿٿ�����"��6	h������e�?�G_BUF/F 1X�]��2	աϸ������� ����!�N�E�W߄� {ߍߺ߱�����������J���DCS� Zr� =����^�+�ZE������|��a�IO 1[
{G ُ!� �!� 1�C�U�i�y������� ��������	-A Qcu�����z��EfPTM  �d�2/ASew �������/ /+/=/O/a/s/�/�/���SEV���.�TYP�/0??y͒�RS@"�|�×�FL 1\
������?�?�?�?0�?�?�?/?TP6���">�NGNA�M�ե�U`�UPSF��GI}�𑪅mA�_LOAD�G �%�%DF_�MOTN���O�@MAXUALRM<���J��@sA�Q����(WS ��@C �]m�-_����MP2�7�^
{k ر�	�!P��+ʠ�;_/��Rr�W�_�WU�W�_�� �R	o�_o?o"ocoNo so�o�o�o�o�o�o�o �o;&Kq\� x������� #�I�4�m�P���|��� Ǐ���֏��!��E� (�i�T�f�����ß�� ӟ���� �A�,�>� w�Z�������ѯ���� د���O�2�s�^� ������Ϳ���ܿ��'��BD_LDXD�ISAX@	��ME�MO_APR@E {?�+
 �  *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT�� Q�c�Ϝ߇��ߧ��� ��w����>�)�b�t� [����{������� ���:���I�[�/��� ���������o����� 6!ZlS�� s����2� AS'�w��� �g��.//R/d/��_MSTR �`�-w%SCD 1am͠L/�/H/�/�/ ?�/2??/?h?S?�? w?�?�?�?�?�?
O�? .OORO=OvOaO�O�O �O�O�O�O�O__<_ '_L_r_]_�_�_�_�_ �_�_o�_�_8o#o\o Go�oko�o�o�o�o�o �o�o"F1jU g������� ��B�-�f�Q���u�𮏙�ҏh/MKCF/G b�-㏕"�LTARM_��c�L�� �σQ�N�<�METP�UI�ǂ���)N�DSP_CMNT�h���|�  d�.��ς�ҟܔ|�_POSCF�����PSTOL 1e�'�4@�<#�
 5�́5�E�S�1�S�U� g�������߯��ӯ� ��	�K�-�?���c�u������|�SING_?CHK  ��;�/ODAQ,�f��Ç���DEV 	�L�	MC:!�HOSIZEh��-��TASK %6��%$123456�789 �Ϡ��T�RIG 1g�+ l6�%���ǃ��0���8�p�YP[� ���EM_INF �1h3� �`)AT&F�V0E0"ߙ�)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ�����ԁH�����A���A�I�q�,��|����  ���ߵ�����J��� n������W������� ����"����X�� /����e���� ��0�T;x�= �as��/�,/ c=/b/�/A/�/�/ �/�/��?��� ^?p?#/�?�/�?s?}/ �?�?O�?6OHO�/lO ?1?C?U?�Oy?�O�O 3O _�?D_�OU_z_a_��_�ONITORG ?5�   �	EXEC1TɃ�R2�X3�X4�XQ5�X���V7�X8�X9Ƀ�RhBLd�RLd �RLd�RLd
bLdbLd "bLd.bLd:bLdFbLcU2Sh2_h2kh2whU2�h2�h2�h2�hU2�h2�h3Sh3_h�3�R�R_GRP?_SV 1in����(ͅ�
�Å���ۯ_MOx�_�D=R^��PL_N�AME !6���p�!Defa�ult Pers�onality �(from FD�) �RR2eq �1j)TUX)TsX��q��X dϏ 8�J�\�n��������� ȏڏ����"�4�F�@X�j�|������2'� П�����*�<�N�`�r��<�������� ү�����,�>�P�tb� �Rdr 1o�y� �\�, ��3���� @D��  ��?�����?x䰺��A'�6�����;�	lʲ	� �xJ������ �< ��"�� �(pK��K ��K=�*�J���J���JV���Zό����rτ́p@j�@T;f��f��ұ]�l���I��p�����������b��3���´  �
`�>�����bϸ�z��w꜐r�Jm��
� B�H�˱]Ӂt��q�	� p��  P�pQ�p�>�p|  Ъ�g����c�	'� �� ��I� ��  ����:��È
�È=����"�s��	�ВI�  �n @@B�cΤ�\��ۤ��t�q�y߁rN���  �'�����@2��@�����/��C��C�C�@� C������
��A�W�@<�*P�R�
h�B�b�A��j�����:����Dz۩��߹������j��( ?�� -��C�`��'�7�����q��Y����� �?�ff ��gy �����q�:a��
>+�  PƱj�(����7	����|�?���xZ�p<
6b�<߈;܍��<�ê<� �<�&Jσ�A�I�ɳ+���?ff�f?I�?&�k�@��.��J<?�`�q�.�˴ fɺ�/��5/���� j/U/�/y/�/�/�/�/��/?�/0?q��F �?l??�?/�?+)��?�?�E�� E��I�G+� F� �?)O�?9O_OJO�OXnO�Of�BL޳B� ?_h�.��O�O��%_�O L_�?m_�?�__�_�_x�_�_�
�h�Îg>��_Co�_`goRodo�o�GA�ds�q�C�o�o�o|����$]Hq�m��D��pC����pCHmZZ7t����6q�q��ܶN'�3�A�A�AR1�AO�^?�$��?�K�0±
�=ç>�����3�W
=�#�\W��e��9������{����<���(�B��u��=B�0�������	L��H�F�G����G��H��U`E���C��+���I#��I��HD��F��E��R�C�j=��
�I��@H�!�H�( E<YD0q�$��H� 3�l�W���{������� �՟���2��V�A� z���w�����ԯ���� ����R�=�v�a� �����������߿� �<�'�`�Kτ�oρ� �ϥ��������&�� J�\�G߀�kߤߏ��� ��������"��F�1� j�U��y������� �����0��T�?�Q�t���(�1��3/�E�����5�������q3�8�x����q4Mgs�&IB+2D�a���{�^ ^	������u%P2P7Q4_A���M0bt��R�������/   �/�b/P/�/ t/�/ *a)_3/�/�/�%1a?�/?;?8M?_?q?  �?�/��?�?�?�?O 2 �F�$�vGb��/�A��@�a�`�qC��C@�o�O2���O�F� DzH@��� F�P D�!��O�O�ys<O!_�3_E_W_i_s?��W�@@pZ.t2�2!2~
 p_�_�_�_	oo -o?oQocouo�o�o�o��o��Q ��+���1��$MSK�CFMAP  ��5� ��6�Q�Q"~�cONR�EL  
�q3�bEXCFE�NB?w
s1uXqF�NC_QtJOGO/VLIM?wdIpMr]d�bKEY?w�u]�bRUN�|�u��bSFSPDT�Y�avJu3sSIG�N?QtT1MOT��Nq�b_CE_�GRP 1p�5s\r���j����� T��⏙������<� �`��U���M���̟ ��🧟�&�ݟJ�� C���7�������گ��������4�V�`TC�OM_CFG 1�q}�Vp�����
�P�_ARC_\r�
jyUAP_CP�L��ntNOCHE�CK ?{ 	r��1�C� U�g�yϋϝϯ����������	��({NO_?WAIT_L�	u6M�NTX�r{�[�m�_ERRY�29sy3� &�������r�c� �촯T_MO��t��,�  ��$�k�3�P�ARAM��u{��V[��!�u?��� =9@345678901��&��� E�W�3�c�����{������� �����=�UM_RSP�ACE �Vv��$ODRDSP����jxOFFSET�_CARTܿ�D�IS��PEN_FILE� �q��c����OPTION_�IO��PWOR�K v_�ms �P(�R�Q
�j.j	 ��Hj&�6$� RG_DS�BL  �5Js��\��RIENTkTO>p9!C��P�q=#�UT__SIM_D
r��b� V� LCT ww�bc��U)+$�_PEXE�d&R�ATp �vju�p��2�X�j)TUX)T�X�##X d -�/�/�/??1?C? U?g?y?�?�?�?�?�?��?�?	OO-O?O�H2 �/oO�O�O�O�O�O�O�O�O_]�<^O;_M_ __q_�_�_�_�_�_�_`�_o���X�OU[��o(��(����$o�, ���IpB` @D��  Ua?�[cAa?��]a]�DWcUa쪞�l;�	lmb�`�xJ�`�����a�<� ��`� ���b, H(��H3�k7HSM5G��22G���Gpc
��
�!��,'|, CR�>�>q��GsuaT�3���  �4spBpyr�  ]o�*SB_�����j]��t3�q� ��r�na �,���6 W ��PQ�|N�M�,k��!�	'� � ���I� � � ��%�=�̡ͭ���ba	����I  �n �@��~���p������ �N U�[�'�!o�:q�pC\�C�A@@sBq�|��� m�O
�A\��h@ߐE�n����Z�B\���A���p� �-�qbz�P��t��_������( �� -��@恊�n�ڥ[A]Ѻ�b�4�'!��(p �?�ff� ��
����!OZ�R��8��z�:��>΁  Pia��(�ವ@���ک�a�c��dF#?����x�����<
6b<�߈;܍�<��ê<� <�#&�o&�)�A�lc�ΐI�*�?fff?��?&c���@�.�uJ<?�`��Yђ^�nd��]e ��[g��Gǡd<���� 1��U�@�y�dߝ߯� �����߼�	���-�������&��"�E��� E��G+� Fþ������������&��J�5��bB��AT�8�ђ��0�6� ��>���J�n�7���[m�0��h�y�1��>�M��I
�@��A�[��C-�)<��?����( /�YĒ��Jp���vav`CH/����x��}!@I�Y��'�3A�A�A�R1AO�^??�$�?�����±
=ç>�����3�W
=�#����+e���ܒ�����{�����<��.�(�B�u���=B0�������	�*H��F�G���G���H�U`E����C�+�-I�#�I��H�D�F��E��RC�j=U>�
I��@H��!H�( E?<YD0/�? �?�?�?�?O�?3OO WOBOTO�OxO�O�O�O �O�O�O_/__S_>_ w_b_�_�_�_�_�_�_ �_oo=o(oaoLo�o �o�o�o�o�o�o�o '$]H�l� ������#�� G�2�k�V���z���ŏ ���ԏ���1��U� g�R���v�����ӟ��������-��(��3������a�����Q�c�,!3ǭ8�}���,!4M�gs����ɢIB+�կ篴a���{���A�/�e�S�(��w��P!�P�������7��ӯ����R9�Kτ�oχ�,�ϥ�  ���χ� ���)��M������ ����{߉ߛ������ߤ�������  )�G�q�_����~��2 F�$�&'Gb���n�[Z,jM!C�s�@j/��A�S���F� D�z��� F�P D��W����)�����������x�?���@@
J9�E�E��E��
 v� �������*<N`�*P ����˨�1��$�PARAM_ME�NU ?-���  �DEFPULS�El	WAIT�TMOUT�R�CV� SH�ELL_WRK.�$CUR_STY�L�,OPT��/PTB./("C��R_DECSN ���,y/�/�/�/�/ �/�/?	??-?V?Q?�c?u?�?�USE_PROG %�q%�?�?�3CCR������7_HOSoT !�!�44O�:T̰�?PCO)A�RC�O�;_TIMqE�XB�  �?GDEBUGV@���3GINP_FL'MSK�O�IT`��O��EPGAP �L̳�#[CH�O�HTY+PE����?�? �_�_�_�_�_oo'o 9obo]ooo�o�o�o�o �o�o�o�o:5G Y�}����������1�Z��EW�ORD ?	7]�	RS`�	P�NS�$��JO�E!>�TEs@WVT�RACECTL �1x-�� ��Ӱ��Ɇ_DT Qy-��~�D � ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�T�(�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_j��_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ�_��� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��������//"#��$PGTRACE�LEN  #! � ���" �8&_UP _z���g!o �S!h 8!_CFoG {g%Q#�"!x!�$J �#|"D�EFSPD |��,!!J �8 I�N TRL }ʇ-" 8�%�!PE�_CONFI� ~>g%�g!�$��%�$LID�#��-74GRP 1��7Q!�#!A ���&ff"!�A+33D�� �D]� CÀ SA@+6�!�" d�$�9�9*1*0� 	� +9�(�&�"�? #´	C�?�;B@3A�O�?OIO3OmO"!>�T?�
5�O��O�N�O =��=#�
�O_�O_ J_5_n_Y_�O}_�_y_x�_�_�_  Dzco" 
oBo�_Roxo co�o�o�o�o�o�o �o>)bM��;�
V7.10b�eta1�$ � A�E�r�ϻ�A " �p?!{G��q>���r���0�q�ͻqB7Q��qA\�p�q��4�q�p�"�B�@�2�D�V�h�w��p�?�?)2{ȏw� ׏���4��1�j�U� ��y�����֟���� ��0��T�?�x�c��� ����ү����!o�,� ۯP�;�M���q����� ο���ݿ�(��L��7�p�+9��sF@ �ɣͷϥ�g%��� ���+�!6I�[߆��� ���ߵߠ��������� !��E�0�B�{�f�� ������������ A�,�e�P���t����� �������=( aL^����� ��'9$]�� ���ϖ������� /<�5/`�r߄ߖߏ/ >�/�/�/�/�/?�/ 1??U?@?R?�?v?�? �?�?�?�?�?O-OO QO<OuO`O�O�O�O�O ���O_�O)__M_8_ q_\_n_�_�_�_�_�_ �_o�_7oIot�� �o�o���o�o�o(/ !L/^/p/�/{*o� �������� A�,�e�P�b������� ���Ώ��+�=�(� a�L���p������Oߟ 񟠟� �9�$�]�H� ��l�~�����ۯƯ�� �#�No`oro�on��o �o�o�oԿ���8 J\ng����vϯ� ��������	���-�� Q�<�u�`�r߫ߖ��� ��������;�M�8� q�\��������z��� ���%��I�4�m�X� ��|����������� :�L�^���Z������ �����$�6�H� Swb��� ����//=/(/ a/L/�/p/�/�/�/�/ �/?�/'??K?]?H? �?��?�?f?�?�?�? O�?5O OYODO}OhO �O�O�O�O�O�O&8 J4_F_����_�_ ��_�_"4-o�O *ocoNo�oro�o�o�o �o�o�o)M8 q\������ ���7�"�[�m��? ����R�Ǐ���֏� !��E�0�i�T���x� �������_$_V_ ��2�l_~_�_�����R��$PLID_KNOW_M  �T?������SV ��U.͠�U��
� �.�ǟR�=�O������mӣM_GRP S1��!`0u��T�@ٰo�ҵ�
 ���Pзj��`��� !�J�_�W�i�{ύϟπ����������߱�MR�����T��s�w� s��ߠ޴߯߅� �ߩ߻�����A��� '��������� ������=���#��� ������}������S��{ST��1 1��U�# ���0�_ A .��,>Pb �������� 3(iL^p������2�*���<-/3 /)/;/M/4f/x/�/�/5�/�/�/�/�6??(?:?7 S?e?w?�?8�?�?��?�?MAD  �d#`PARNUM  qw�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a�OT>_CMP_��B@��P@'˥TER�_CHK'U��0˪?R$_6[RSl�¯���_MOA@�_�U_��_RE_RES_G ��>�oo8o +o\oOo�oso�o�o�o �o�o�o�o�W �\�_%�Ue Baf �S� ����S0� ���SR0��#��S �0>�]�b��S�0}���<���RV 1�����^rB@c]��t�_(@c\����_D@c[�$���RTHR_INRl��DA��˥d,�MASmS9� ZM�MN8��k�MON_QUEUE ���˦��Vx� RDNPUbQqN{�P[��END���_ڙEXE�ڕ�@�BE�ʟ��OPT�IOǗ�[��PROGRAM %���%��ۏ�O��TA�SK_IAD0�OCFG ���tO��^ŠDATA���Ϋ@��27�>�P� b�t���,�����ɿۿ������#�5�G���IWNFOUӌ���� ���ϭϿ�������� �+�=�O�a�s߅ߗ� �߻��������^�jč�� yġ?PDIT �ίc���WERFL
��
�RGADJ �&n�A����?�����@���IORITY�{�QV���MPDSQPH�����Uz��ޝ�OTOEy�1��R� (!AF�4�E�P]���!�tcph���!�ud��!icqm��ݏ6�XY_ȡ��R��ۡ)�� *+/ ۠� W:F�j�� ����%7�[B�*��POSRT#�BC۠�����_CARTR�EP
�R� SKS�TAz��ZSSAV����n�	2500H863���r�T$!�R���Áq�n�}/�/�'� U�RGE�B��rYW�F� DO{�rUVW�V��$�A�WRUP�_DELAY ��R��$R_HOT�k��%O]?�$R_?NORMALk�L?<�?p6SEMI?�?|�?3AQSKIP!��n�l#x 	 1/+O+ OROdOvO9H n��O�G�O�O�O�O�O _�O_D_V_h_._�_ z_�_�_�_�_�_
o�_ .o@oRoovodo�o�o �o�o�o�o�o*< Lr`���n��$RCVTM�v����pDCR!��LЈqC`N��C���C��Q?��>r�ߝ<|�{4M�g��&��/���Z��t����?l4�{�4Oi���O <
6b<�߈;܍�>�u.�?!<�&{�b�ˏݏ�� 8�����,�>�P�b� t���������Ο��� ݟ��:�%�7�p�S� �����ʯܯ� �� $�6�H�Z�l�~����� ��ƿ���տ���2� D�'�h�zϽ��ϰ��� ������
��.�@�R� d�Oψߚ߅߾ߩ��� ������<�N��r� ������������ �&�8�#�\�G����� }�����������S� 4FXj|��� ������0 T?x�u��� �'//,/>/P/b/ t/�/�/�/�/�/�/� ?�/(??L?7?p?�? e?�?�?��?�? OO $O6OHOZOlO~O�O�O �?�?�O�O�O�O __ D_V_9_z_�_�?�_�_ �_�_�_
oo.o@oRo�dovo�X�qGN_A�TC 1�� �AT&FV�0E0�kAT�DP/6/9/2{/9�hATA�n�,AT%G�1%B960�i�+++�o,�aH�,�qIO_TY�PE  �u�s�n_�oREFPOS�1 1�P{ x�o�Xh_�d_ �����K�6�o� 
���.���R����{{/2 1�P{����؏V�ԏz����q3 1��$�6�p��ٟ|���S4 1������˟���n���%�S5 1�<�N�`������<���S6 1�ѯ���/�����ѿ>O�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASKw 1�P  
9ߜG��XNOM����a~߈ӁqMOTE�  h�~t��_CFG ������рrPL_RANG����Q��POWER ���e��SM�_DRYPRG �%i�%��J��T?ART �
�X�UME_PRO'��9��~t_EXEC_ENB  �e��GSPD�����蜩c��TDB���R�M��MT_!�T����`OBOT�_NAME �i���iOB_O�RD_NUM ?�
�\qH?863  �T���������bPC_TIMEOUT��{ x�`S232���1��k L�TEACH PE�NDAN �ǅ��}���`Mai�ntenance Cons�R}�m
�"{�dKCL/!Cg��Z ��n�� No Us�e}�	��*NPqO��х��ӽ(CH_L��������	�mMAVAIL��{���ՙ�SPACE�1 2��| �d��(>��&����p��M,8�?�ep/eT/�/�/�/ �/�W//,/>/�/b/ �/v?�?Z?�/�?�9�e �a�=??,?>?�?b? �?vO�OZO�?�O�O�Os�2�/O*O <O�O`O�O�_�_u_�_�_�_�_[3_#_5_ G_Y_o}_�_�o�o�o �o�o[4.o@o Rodovo$�o�o��@��"�	�7�[5K ]o��A���菀	�̏�?�&�T�[6 h�z�������^�ԏ�� �&��;�\�C�q�[7��������͟{�� �"�C��X�y�`���[8����Ưدꯘ� �0�?�`�#�uϖ�}ϼ��[G �i�� �ϋ
G� ����$�6�H�Z�l� ~ߐ��8 ǳ���������d(���M� _�q�������� ���?���2�%�7�e� w��������������� �����!�RE�W�� ��������p?Q `�� @0��ߖrz	�V_��� ��
/L/^/|/2/d/ �/�/�/�/�/�/?�/ �/�/*?l?~?�?R?�? �?�?�?�?�?�?2O�?�
��O[_MO�DE  �˝IS ���vO,*Aϲ�O-_��	M_�v_#dCWORK_�AD�M,�$bR  ��ϰ�P{_��P_INTVAL��@����JR_OPoTION�V �E�BpVAT_GR�P 2�����(y_Ho � e_vo�o�oYo�o�o�o �o�o*<�bOo NDpw����� �	���?�Q�c�u� ����/���ϏᏣ��� �)�;���_�q����� ����O�ɟ���՟ 7�I�[�m�/������� ǯٯ믁��!�3��� C�i�{���O���ÿտ ���ϡ�/�A�S�e� 'ωϛϭ�oρ����� ��+�=���a�s߅� Gߕ߻����ߡ��� '�9�K�]��߁��� ��y����������5��G�Y��E�$SCAN_TIM�AYue�w�R �(ӿ#((�<0.a�aPaP
Tq>��Q��oa�����OOE2/���d;D2BaR��WY���^���^R^	r � P��� �  8�P�	<�D��G Yk}���������Qp�/@/R//)P;��o\T��Qpg-�t�_DiKT|��[  � l v%������/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OWW�#�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_olO~Od+No`o ro�o�o�o�o�o�o�o &8J\n�������u�  0�"0g�/�-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ����$o��˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�����Do������ ��ҿ�����,�>� P�b�tφϘϪϼ���`������w
�  5 8�J�\�n߀ߒߜկ� ��������	��-�?�Q�c�u����� ��-����� � 2�D�V�h�z��������������������& ��%	�12345678^�" 	��/� `r��������(: L^p����� �� //$/6/H/Z/ l/~/��/�/�/�/�/ �/? ?2?D?V?h?�/ �?�?�?�?�?�?�?
O O.O@Oo?dOvO�O�O �O�O�O�O�O__*_ YON_`_r_�_�_�_�_ �_�_�_ooC_8oJo \ono�o�o�o�o�o�o �oo"4FXj�|������� ��	��s3�E�W��{�Cz  Bp���   ��2����z�$SCR_�GRP 1�(��U8(�\x�^ @ > 	!��	  ׃���"�$� ���-��+��R�w����D~�����#�����O���M-�10iA 890�9905 Ŗ5 M61C >4��J*ׁ
� ����0�����#�1�	�"�z�������¯Ҭ ���c��� O�8�J��������!�����ֿ��B�By���������A��$�  @��<� �R�?��d���Hy�u�O����F@ F�` �§�ʿ�϶������� %��I�4�m��<�l�`�߃ߕߧ߹�B��� \����1��U�@�R� ��v������������;���*<=�
�F���?�d�<�>HE�����@�:��� B���ЗЙ����EL_DEFA�ULT  ���_�B��MIPOWERFL  �$1 oWFDO $���ERVENT �1�����"��pL!DUM_�EIP��8��j!AF_INE <�=�!FT����!��4 ���[!RPC�_MAIN\>�8J�nVISw=y���!TP��PU��	d�?/!�
PMON_PR'OXY@/�e./�/�"Y/�fz/�/!RDM_SRV�/r�	g�/#?!R dC?�h?o?!
p�M�/�i^?�?!?RLSYNC�?8��8�?O!ROS�.L�4�?SO" wO�#DOVO�O�O�O�O �O_�O1_�OU__._ @_�_d_v_�_�_�_�_�o�_?oocoiICE_KL ?%y� (%SVCPRG1ho8��e��D�o�m3�o�o�`4 D�`5(-�`6PU�`7x}�`���l9��{�d:?� �a�o��a�oE��a�o m��a���aB���a j叟a���a�5� �a�]��a����a3� ���a[�՟�a�����a ��%��aӏM��a��u� �a#����aK�ů�as� ��a��mob�`�o�` 8�}�w�������ɿ�� �ؿ���5�G�2�k� VϏ�zϳϞ������� ���1��U�@�y�d� �߯ߚ��߾������ �?�*�Q�u�`��� ����������;� &�_�J���n������������sj_DEV� y	�M{C:L!`OUT",?REC 1�Z� �d   	 	������

 �Z�{ 0H6lZ�~� ����� //D/ 2/h/z/\/�/�/�/�/ �/�/�/?�/,?R?@? v?d?�?�?�?�?�?�? �?OO(ONO<OrOTO fO�O�O�O�O�O�O_ &__J_8_Z_\_n_�_ �_�_�_�_�_�_"oo Fo4oVo|o^o�o�o�o �o�o�o�o0T Bxf����( ���,��P�>�`� ��h���������Ώ� �(�:��^�L���p� ������ܟ���� � 6�$�Z�H�~���r��� ��دƯ����2�� &�h�V���z�����Կ �ȿ
�����.�d� RψϚ�|ϾϬ����� ����<��`�N�p� �߄ߺߨ�������� �8�&�\�J�l��joV 1�w P�l�	� � ��F��
TYP�EVFZN_C�FG �x��d7�GR�P 1�A�c �,B� A� D;� B���  �B4RB2�1HELL:�4(
 X���>�%RSR���� E0iT�x� �����/�Sew�  ��%w������#����)�A�2#�d�����HK 1��� ���m/h/z/�/�/ �/�/�/�/�/
??E? @?R?d?�?�?�?�?��?OMM ����?���FTOV_EN�B ���+�HOW_?REG_UIO��IMWAITB\�JKOUT;F���LITIM;E��ΆOVAL[OMC_U�NITC�F+�MO�N_ALIAS �?e�9 ( he�s_(_:_L_^_�� _�_�_�_�_j_�_�_ oo+o�_Ooaoso�o �oBo�o�o�o�o�o '9K]n�� ��t���#�5� �Y�k�}�����L�ŏ ׏������1�C�U� g����������ӟ~� ��	��-�?��c�u� ������V�ϯ��� ���;�M�_�q���� ����˿ݿ����%� 7�I���m�ϑϣϵ� `�������ߺ�3�E� W�i�{�&ߟ߱����� �ߒ���/�A�S��� w����X������ ����=�O�a�s��� 0������������� '9K]��� �b���#� GYk}�:�� ����/1/C/U/  /f/�/�/�/�/l/�/ �/	??-?�/Q?c?u? �?�?D?�?�?�?�?O �?)O;OMO_O
O�O�O �O�O�OvO�O__%_�7_�C�$SMON�_DEFPRO ����`Q� *S�YSTEM*  �d=OURECA�LL ?}`Y �( �}4xco�py fr:\*�.* virt:�\tmpback��Q=>192.1�68.4�P46:8736 �R�_�_,�_�K}5�Ua�_�_`�V�_goyo�o}9�T�s:orderf?il.dat.l@o�Vo�o�o}0�Rmdb:+o�o�Q�ob t�c�_2o?U� �
�o��Sod�v�����
xyzra?te 61 +�=� O����������504 *�ҏc�u� ���o�o56�ٟ��� "��5�џb�t���r�6����emp:�2164 W����:��.��*.d��Ʈ`ϯ`�r�����1 +� =�O�����)�Ҳ ��ҿc�uχϚ���5� ͧ�������"���̨ ��b�t߆ߙ����Q� U�����
������N� ��h�z��ϱ�:��� ����
�߸�A���d� v�����.�;������� ����O�`r� ���2������ '��K�\n����� 8�����#� G/j/|/����3/E/�W/�/�/�/��w1356?��/b?t?�?� �458�?�?�?" �?58�?bOtO�O���?|���p6088 WO �O�O�O��O�I�O`_ r_�_�/��;_M_�_�_ o?'?�T�_�_couo �o�?�?5O�G�o�o�o O"O�o�H�obt� ��/�/:dV���/��8 �g�y� ���o�o9T���	� ��@ҏc�u�������$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1����?���%֟ ��&�	��\�?�f� ��u��������ϯ�� "��F�)�;�|�_��� ����ֿ��˿��� B�%�f�I�[Ϝ�Ϧ� �ϵ�������,��6� b�E߆�i�{߼ߟ��� ��������L�/�V� ��e��������� ���6��+�l�O�v� �������������� 2V9K�o� ������& R5vYk��� ��/��<//F/ r/U/�/y/�/�/�/�/ ?�/&?	??\???f? �?u?�?�?�?�?�?�? "OOFO)O;O|O_O�O �O�O�O�O�O_�O_ B_%_f_I_[_�__�_ �_�_�_�_�_,oo6o boEo�oio{o�o�o�o �o�o�oL/V �e������ ��6��+�l�O�v��������PARAM� ����� ��	��P�����OFT_K�B_CFG  �ヱ���PIN_S_IM  ����C�U�g�����RVQSTP_DSB,��򂣟����SR ��/�� & � ULTIROB?OTTASK������TOP_ON_ERR  ����PTN �/�@�A�	�RING_PR�M� ��VDT_GRP 1�ˉ�  	������ ������Я����� *�Q�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߣߠ߲������� ����0�B�i�f�x� ������������� /�,�>�P�b�t����� ����������( :L^p���� ��� $6H Z�~����� ��/ /G/D/V/h/ z/�/�/�/�/�/�/? 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�__\_��VPRG_�COUNT��8@���RENBU��U�M�S��__UPD� 1�/�8  
s_�oo*oSoNo `oro�o�o�o�o�o�o �o+&8Jsn �������� �"�K�F�X�j����� ����ۏ֏���#�� 0�B�k�f�x������� ��ҟ������C�>� P�b���������ӯί������UYSDOEBUG�P�P�)��d�YH�SP_PA�SS�UB?Z�L�OG ��U��S)�#�0�  ���Q)�
MC:�\��6���_MPC ���U���Qñ8�� �Q�SAV ������ǲ&��ηSV;�TEM_TIME 1��[� (m��&�����}YT1SVGU�NS�P�U'�U����ASK_OPT�ION�P�U�Q�Q���BCCFG ��[u� n�A�a�`a�gZo��߃� ���߹�������:� %�^�p�[����� ���� �����6�!�Z� E�~�i���������&�������&8�� nY�}�?��� � ��(L: p^������ �/ /6/$/F/l/Z/ �/~/�/�/�/�/�/�/ �/2?8 F?X?v?�? �??�?�?�?�?�?O *O<O
O`ONO�OrO�O �O�O�O�O_�O&__ J_8_n_\_~_�_�_�_ �_�_�_o�_ o"o4o joXo�oD?�o�o�o�o �oxo.TBx ��j����� ���,�b�P���t� ����Ώ��ޏ��(� �L�:�p�^������� ʟ��o��6�H� Z�؟~�l�������د ���ʯ ��D�2�h� V�x�z���¿���Կ 
���.��>�d�Rψ� vϬϚ��Ͼ������� *��N��f�xߖߨ� ��8���������8� J�\�*��n����� ��������"��F�4� j�X���|��������� ����0@BT �x�d���� �>,Ntb� �����/�(/ /8/:/L/�/p/�/�/ �/�/�/�/�/$??H? 6?l?Z?�?~?�?�?�? �?�?O�&O8OVOhO zO�?�O�O�O�O�O�O 
__�O@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<o^o�oro�o �o�o�o�o�o  J8n$O���� �X���4�"�X��B�v��$TBCS�G_GRP 2��B�� � �v� 
 ?�  ������׏�� �����1��U�g�z����ƈ�d, ����?v�	 HC{��d�>����~e�CL  B����Пܘ������\)��Y  A��ܟ$�B�g�B�Bl��i�X�ɼ���X��  D	J���r������C����үܬ���D�@v�=�W�j�}� H�Z���ſ���������v�	V�3.00��	mw61c�	*X�0P�u�g�p�>���v�(:�� ��p͟�w  O����p������z�JCFG [�B��� ��V��������=��=�c�q�K� qߗ߂߻ߦ������ ��'��$�]�H��l� ������������#� �G�2�k�V���z��� �����������p *<N���l�� �����#5G Y}h���� v�b��>�// /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?d?R? t?v?�?�?�?�?�?O �?*OO:O`ONO�OrO �O�O��O�O�O_&_ _J_8_n_\_�_�_�_ �_�_�_�_�_�_oFo 4ojo|o�o�oZo�o�o �o�o�o�oB0f T�x����� ��,��P�>�`�b� t�����Ώ������ �&�L��Od�v���2� ����ȟʟܟ� �6� $�Z�l�~���N����� دƯ�� �2��B� h�V���z�����Կ¿ ����.��R�@�v� dϚψϪ��Ͼ����� ��<�*�L�N�`ߖ� �ߺߨ����ߚ��� ����\�J��n��� ��������"���2� X�F�|�j��������� ������.TB xf������ �>,bP� t�����/� (//8/:/L/�/�ߚ/ �/�/h/�/�/�/$?? H?6?l?Z?�?�?�?�? �?�?�?O�?ODOVO hO"O4O�O�O�O�O�O �O
_�O_@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<oro`o�o �o�o�o�o�o�o& �/>P�/��� ������4�F� X��(���|�����֏ ����Ə0��@�B� T���x�����ҟ���� ��,��P�>�t�b� ������������� �:�(�^�L�n����� ��2d�����̿� $�Z�H�~�lϢϐ��� �����Ϻ� ��0�2� D�zߌߞ߰�j����� �����
�,�.�@�v� d����������� ��<�*�`�N���r� ������������& J\�t��B ������F 4j|��^��p��/�  2 �6# 6&J/6"��$TBJOP_G�RP 2����  ?i�X,i#�p,� ��x�J� �6$�  �_< �� �6$� @2 �"	 ߐC�� �&b � Cق'�!�!>�c��
559>�0�+1�33=�{CL� fff?+0?�ffB� J1�%�Y?d7�.��/>��2\)?0�5����;��hC=Y� �  @� �!?B�  A�P?�?��3EC�  Dp�!�,�0*BOߦ?��3JB��
:���Bl�0��0�$�1��?O6!Aə�A�ДC�1D�G6��=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH��1ts�A@333@?1� C�� �@�_�_&_8_>��D��UV_0�LP�Q30<'{�zR� @�0�V �P!o3o�_<oRifoPo ^o�o�o�oRo�o�o�o �oM(�ol�pP~��p4�6&�q�5	V3.00��#m61c�$�*(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�N�aF���F�^�lF���F�:�
F�)F���3G�G���G��G,I�R�CH`�C��dTDU�?D���D��DE(�!/E\�E���E�h�E��ME��sF�`F+'\FD���F`=F}�'�F��F��[
F���F���M;S@;Q�*�|8�`rz@/&�
8�6&<��1�w��^$ESTPARS�  *({ _#HR���ABLE 1̒p+Z�6#|�Q� (� 1�|�|�|�5'T=!|�	|�
|�|�T˕6!|�|�|����RDI��z!�ʟܟ� ��$���O ������¯ԯ�����	S��x# V���˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �U-����ĜP�9�K� ]�o��-�?�Q�c�u����6�NUM  V�z!� > � Ȑ����_CFGG �����!@b �IMEBF_TT�����x#��a�VER腣b�w�a�R 1=�p+
 (3�6"	1 ��  6!���� ������ �9�$�:�H� Z�l�~����������� ����^$��_���@x�
b MI_CWHANm� x� k�DBGLV;0o��x�a!n ETHER_AD ?�� �y�$"�\&n oROUT��!p*�!*�SNM�ASK�x#�255.h�fx^$�OOLOFS_D�I��[ՠ	ORQCTRL �p+ ;/���/+/=/O/ a/s/�/�/�/�/�/���/�/�/!?��PE_�DETAI��P�ON_SVOFF��33P_MON ��H�v�2-9ST�RTCHK ����42VTCOMPATa8�24:0�FPROG %��%MULTI?ROBOTTO!O<06�PLAY��L:_INST_MPe GL7YDUS���?�2LCK�LPKQ?UICKMEt �O��2SCRE�@>�
tps��2 �A�@�I��@_Y����9�	SR_GRP� 1�� ���\�l_zZg_�_ �_�_�_�_�^�^�o j�Q'ODo/ohoSe� �oo�o�o�o�o�o�o !WE{i�������	1?234567���!���X�E1�V[
� �}ipnl�/a�gen.htmno��������ȏ~��Panel _setup̌}�?���0�B�T�f�  ��񏞟��ԟ��� o����@�R�d�v��� ���#�Я����� *���ϯůr������� ��̿C��g��&�8� J�\�n�����϶��� ������uϣϙ�F�X� j�|ߎߠ����;��߀����0�B��*NU�ALRMb@G ?�� [���� �������� ��%�C��I�z�m�������v�S�EV  �����t�ECFG �Ձ=]/BaA$ �  B�/D
  ��/C�Wi{�� ����� PRց; �To\�o�I�6?K0(% ����0����� //;/&/L/q/\/�/0�/�/l�D �Q��/I_�@HIST� 1ׁ9  �(  ��(/�SOFTPART�/GENLINK�?current�=menupag�e,153,1 �Ec0p?�?�?�?/C�s� >?P=962n?��?
OO.O�?�?�136c?|O�O�O�OAOSO �?�O__0_�O�O_L u_�_�_�_:_�/�_�_ oo)o;o�__oqo�o �o�o�oHo�o�o%7I~��a81�ou ������o�� �)�;�M��q����� ����ˏZ�l���%� 7�I�[��������� ǟٟh����!�3�E� W����������ïկ �v���/�A�S�e� Pb������ѿ��� ���+�=�O�a�s�� �ϩϻ�������ߒ� '�9�K�]�o߁�ߥ� ���������ߎ�#�5� G�Y�k�}������ ���������1�C�U� g�y���v��������� ��	�?Qcu ��(���� )�M_q�� �6���//%/ �I/[/m//�/�/�/ D/�/�/�/?!?3?�/ W?i?{?�?�?�?���� �?�?OO/OAOD?eO wO�O�O�O�ONO`O�O __+_=_O_�Os_�_ �_�_�_�_\_�_oo 'o9oKo�_�_�o�o�o �o�o�ojo�o#5 GY�o}�������?��$UI_�PANEDATA 1������  	�}�0�B�T�f�x��� )����mt�ۏ ����#�5���Y�@� }���v�����ן���� ���1��U�g�N���.��� �1��Ï ȯگ����"�u�F� ��X�|�������Ŀֿ =������0�T�;� x�_ϜϮϕ��Ϲ������,ߟ�M��j� o߁ߓߥ߷������ `��#�5�G�Y�k��� ������������� ��C�*�g�y�`��� ������F�X�	- ?Qc����߫� ���~;" _F��|��� ��/�7/I/0/m/ �����/�/�/�/�/�/ P/!?3?�W?i?{?�? �?�??�?�?�?O�? /OOSOeOLO�OpO�O �O�O�O�O_z/�/J? O_a_s_�_�_�_�O�_ @?�_oo'o9oKo�_ oo�oho�o�o�o�o�o �o�o#
GY@} d��&_8_��� �1�C��g��_���� ����ӏ���^��� ?�&�c�u�\������� ϟ���ڟ�)��M� ����������˯ݯ 0�����7�I�[�m� ���������ٿ�ҿ ���3�E�,�i�Pύπ�φ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#������� � �$�6��Z�A�~�e� w����������� 2��V�h�O�����v��p��$UI_PA�NELINK 1��v�  ��  ���}1234567890����	- ?G ���o��� ��a��#5�G�	����p&���  R���� �Z��$/6/H/Z/ l/~//�/�/�/�/�/ �/�/
?2?D?V?h?z? ?$?�?�?�?�?�?
O �?.O@OROdOvO�O O �O�O�O�O�O_�O�O�<_N_`_r_�_�_�0,���_�X�_�_�_ o 2ooVohoKo�ooo�o �o�o�o�o�o�� ,>r}������ ������/�A� S�e�w��������я ���tv�z���� =�O�a�s�������0S ��ӟ���	��-��� Q�c�u�������:�ϯ ����)���M�_� q���������H�ݿ� ��%�7�ƿ[�m�� �ϣϵ�D�������� !�3�Eߴ_i�{�
�� �����߸������/� �S�e�H���~�� R~'�'�a��:�L� ^�p������������� �� ��6HZl ~���#�5���  2D��hz� ����c�
// ./@/R/�v/�/�/�/ �/�/_/�/??*?<? N?`?�/�?�?�?�?�? �?m?OO&O8OJO\O �?�O�O�O�O�O�O�O [�_��4_F_)_j_|_ __�_�_�_�_�_�_o �_0ooTofo��o�� �o��o�o�o, >1bt���� K����(�:�� ��{O������ʏ܏ �uO�$�6�H�Z�l� ��������Ɵ؟��� �� �2�D�V�h�z�	� ����¯ԯ������ .�@�R�d�v������ ��п���ϕ�*�<� N�`�rτ��O�Ϻ�Io ���������8�J�-� n߀�cߤ߇����߽� ���o1�oX��o|� ������������ �0�B�T�f������ ��������S�e�w�, >Pbt��'� ����:L ^p��#��� � //$/�H/Z/l/ ~/�/�/1/�/�/�/�/ ? ?�/D?V?h?z?�? �?�???�?�?�?
OO .O��ROdO�߈OkO�O �O�O�O�O�O_�O<_ N_1_r_�_g_�_7O�M�m�$UI_�QUICKMEN�  ���_AobREST�ORE 1��  �A|��Rto�o�im�o �o�o�o�o:L ^p�%���� ��o����Z�l� ~�����E�Ə؏��� � �ÏD�V�h�z��� 7�������/���
�� .�@��d�v������� O�Я�����ßͯ 7�I���m�������̿ ޿����&�8�J�� nπϒϤ϶�a����� ��Y�"�4�F�X�j�� �ߠ߲������ߋ����0�B�T�gSCR�E`?#m�u1sco`u2���3��4��5��6ʏ�7��8��bUS#ERq�v��Tp���Sks����4��5��6��7��8��`N�DO_CFG m�#k  n` `PDATE ����None�bSEUFRAM/E  �TA�n��RTOL_ABRqTy�l��ENB��~��GRP 1�ci�/aCz  A� ����Q�� $6BHRd��`U������MSK  h�����Nv�%�U��%���bVIS�CAND_MAXλI��FA?IL_IMG� �P�ݗP#��IMR_EGNUM�
,�[SIZ�n`��A�,VONTM�OU��@����2��a��a�����FR�:\ � �MC:\�\L�OG�B@F� �!�'/!+/O/�Uz MCV��8#UD1r&EX�{+�S�PPO6�4_��0'fnm6PO��LIb��*�#V���,fy@�'�/� =	�(wSZV�.����'�WAI�/STAOT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_J�MPERR 1��#k
  �2345678901dF �ψO{O�O�O�O�O�O _�O*__N_A_S_�_<
� MLOWc>
 ��_TI�=�'�MPHASE'  ��F��P�SHIFT�1 9�]@<�\�Do �U#oIo�oYoko�o�o �o�o�o�o�o6 lCU�y��� �� ��	�V�-�e�2����	VSF�T1�2	VMN�� �5�1G� ����%A�  B8*̀̀�@ pكӁb˂�у��z�ME@Ľ?�{��!c>&%��aM1��k�0��{ �$`0TDINGEND��\�O� �z����S��w��P���ϜREL�E�Q��Y���\�_ACTIV��:�R�A ��e����e�:�RD� ���Y?BOX �9�دV�6��02����190.0.��83��2�54��QF�	 ��X�j��1�?robot���   p��<���5pc��̿ �����7�����-�f�ZABC�����, ]@U��2ʿ�eϢω� �ϭϿ����� ��߀V�=�z�a�s߰�E�Z��1�Ѧ