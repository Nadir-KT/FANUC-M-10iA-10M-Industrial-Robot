��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �� �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1���|URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y12 � u3�|4|�RG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�&�ASBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�:OF�F_ N�3DELHLOGn25Aa2�?i1@N?�(� -M�H W+0�$=Y $DB� 6�COMW!2MO�� 21\D.	 \vrVE�1$F��A{$O��D�B~�CTMP1_F�E�2�G1_�3�B�2��GXD�#
 �d $CARD�_EXIST4�$FSSB_TY�PuAHKBD_YS�B�1AGN Gn� $SLOT�_NUMJQPREV,DBU� g1� �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��AETE_OK�RUS�P_CR�Q$;4�V� 0LACIw1�RAP�k �1x@ME@$D�V�Q�Pv�Ah{oQL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa4 hq;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I�9�TY�D,P*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6��U7��8��94�� ;CO�$ <� �$6xK3 1w`O_M|�@�C t � �E#6NGP�ABA� �c��ZQ���`����@nr��� ��P`�0���p� �v�p�PzPb26����"MJ�_R��BC�1J��3�JVP���tBS��}Aw��"�tP�_*0OFSzR @� RO_K8���a�IT�3��NOM_��0�1ĥ3�ACPT �� $���2AxP��K}EX�� ��0g0I01��p�
$�TFa��C$MD3&��TO�3�0U� ��/ �Hw2�C%1|�EΡg0wE{`vF�vF�40CPp@��a2 
P$A`PqU�3N)#��dR*�AX�!sDET;AI�3BUFV��p@1 |�p۶�pkPIdT� PP[�EMZ�Mg�Ͱj�F[�SIMQSI�"0�ȪA.�����lw 	Tp|zM��P�B��FACTrbHPE�W7�P1Ӡ��v��M]Cd� �$*1�JB�p<�*1DEC�Hښ�H���b� �� +PNS_E;MP��$GP���B,P_��3�p�@Pܤ��TC��|r��0�s ��b�0�� �B���!
����JR� ��SEGKFR��Iv �aR��TkpN&S,�PVF����� & k�Bv�u�cu��aE�� �!2��+�MQ��E�SI!Z�3����T��P������aRSINF �����kq���������LX�����F�C3RCMu�3CClpG� �p���O}���b�1��������2�V�DxIC��C���r����P��L{� EV �zF�_��F�pNB0��?������A�! �r�Rx����V�lp �2��aR�t�,�g��}RTx #� 5�5"2��uAR���`�CX�$LG�p��B@�1 `s�P�t�aA�0�{�У+0R���tM�E�`!BupCrRA 3tAZ�л�pc��OT�FC�b�`�`F�Np���1��ADI +�a%��b�{��p $�pSp�c�`S�P�L�a,QMP6�`Y�3���M'�pU��aU�  $>�TITO1�S�S�!��$�"0�DBPXWO��z!��$SK���2��DB�"��"@�PR8� 
p� ���# >�6q1$��$��+ЅL9$?(�V�%�@?R4C&_?R4E3NE��'~?(��� RE�pY2(H� �OS��#$L�3$$3R��;43�MVOk_D@!V�ROScrr�w�S���~CRIGGER2F�PA�S��7�ETUsRN0B�cMR_���TUː[��0EW5M%���GN>`��FRLA���Eݡ�P��&$P�t�'��@4a��C�DϣV�D�XQ��4�1��MVGO�_AWAYRMO�#�aw!� CS_�)  `IS #� �� �s3S�AQ汯 4Rx�ZSW�AQȉp�@1UW��cTNT	V)�5RV
a���|c�éWƃ��JB��x0���SAFEۥ�V_�SV�bEXCLUtU�;��ONL��bcYg�~az�OT�a{�HI_V? ��S<, M�_ *�0� r��_z�2� �"vPSGO  +�r Ɛm@�A�c~b���w@♐V�i�b�fANNcUNx0�$�dIDY�	UABc�@Sp�i�a�+ �j�f�Ca�pOGuIx2,��$F�b̫$ѐOT�@A $DUMMY��Ft��Ft±� 6U�- ` !�HE��|s��~bc�B@ SoUFFI��4P�CA�Gs5Cw6�Cq��DMSWU.{ 8��KEYI��5�TM�1�s�qoA�vINޱw�X� , �/ D��HOST�P!4���<���<�0°<��p<�EM'����Z�� SBL� UL>��0  �	���w�CaT�01 ϴ $��9USAMPLо�/����ĺ�$ I@갯 $SUBӄ��w0QS��8���#��SAV������c�S< 9�`�fP�$�0E!� YN_�B�#2 0��DI��d�pO|�m��#$�F�R_IC� �?ENC2_Sd�3  ��< 3�9����� cgp����4��"��2�A��ޖ5���`ǻ�@Q@�K&D-!�a�AVE�R�q����DSP
���PC_�q��"�x|�ܣ�VALU3��HE�(�M�IP\)���OPPm �CTH�*��S" $T�/�Fb�;�d�����d ����ET6� H(rLL_DU ǀ�a�@��k���֠COT�"U�/��q~@@NOAUTO70�$}�x�~�@s���|�C͠��C�� 2�!z�L�� �8H *��L � ���Բ@sv��`�  �� ÿ���Xq��cq��P�q���q��7��8���9��0���1�1� �1-�1:�1G�1�T�1a�1n�2|�2T��2 �2-�2:�U2G�2T�2a�2nʕ3|�3�3� �3�-�3:�3G�3T�3�a�3n�4|&q����9 <���z�ΓKI����H���ͰFEq@{@�: ,��&a? P_P?��>���%��E�@��C`QQ���;fp$TP~�$VARI���r��\@P2Q`< W�߃TD��g���`���������BAC��"= T2����$)�,+r³�p IFI@��p�� q M�P"�Ɛ�Fl@``>�t ;��6����ST����T��M ����0	��i��� F���������kRt �����FORCEUP��b܂FLUS
pH�(N��� ��6bD_CM�@E�7N� p(�v�P��REM� Fa��@j��ʥ
K�	N���EF1F/���@IN�QsOV��OVA�	�TROV DT<)��DTMX:e  �P:/��Pq�v,XpCLN _�p���@ ��	_|��_T�: �|�&PA�QDI���1��L0�Y0RQm�_+qdH���M���CL�d�#�RIV{�ϓN"E�AR/�IO�PC�P��BR��CM؍@N 1b 3GC3LF��!DY�(�lq�#5T�DG����� �%�&�FSS� )�? P(q1�1��`_1"811R�EC13D;5D6O�GRA���@��i���PW�ON2EBUG�S�2��Ͱgϐ_E A� ��?�����TERM�5B�5?��ORIw�0�C�5݁�SM�_-`���0D�5EG�.�TA�9E�5n� S�UP��Fg� -QϒA�P|�3�@B$SEGGJv� EL�UUSEPNFI��pBx��1x@��4>DC$UF�P��$���Q�@C���G�0T�����SwNSTj�PATۡ<g��APTHJ�A�E*�Z%qB\`F�{E���F�q�pARxPY�aS�HFT͢qA�AX_�SHOR$�>��6 �@$GqPE���O#VR���aZPI@P@$�U?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi� [Y)��G�@R��i�e԰�i�R�!P�uAScYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UaP���P���WOR�@�M��k0SMT��G��GR��3�a�PA�@��p5�'�H� � j�A�T�OCjA7pP]Pp$OPd�O��C�%��p�O!��RE.pR�C�AO�?��Be5pR�EruIx'Q�G�e$PWR) IMdu�RR_$sp�5�.�B Iz2H8�=��_ADDRH�H_LENG�B�q�q:��x�R��So�J.�SS��SK������ ��-�SE*���rmSN�MN1K	��j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ���p�Q� ��OUPW3��b_>�I��!q�a1 ��������|��� �����-���:���i+IOX2S=�D�e���^���L $x��p�!_OFF[r�_�PRM_��^�aTTP_�H��wM (�pOBJ�"l�pG�$H�LE�C���ٰN � \9�*�AB_�T��b
�S�`�S��LV���KRW"duHITC�OU?BGi�LO�q����d� Fp�k�GpSS� ���HQWh�wA��O.��`�INCPUX2VISIO��!��¢.��á<�á-� �IO�LN)�P 87�R�'�[p$SL�b�d PUT_��$�dp�Pz �� F�_AS2Q/�$ALD���D�aQT U�0�]P�A������PH�YG灱Z��5�UO� 3R `F���H�@Yq�Yx�ɱvpP�S�dp���x��ٶ1 ��UJ��S����NEΊWJOG�G �DI�S��r�KĠ��3T� |��AV��`_�C�TR!S^�FLAG�f2r�LG�dU ��n�:��3LG_SIZ��ň��=���FD��I����Z  �ǳ��0�Ʋ�@s��-� ��-�=�-���-��0-�ISCH_��Dq���N?���V��EE !2�C��n�U����r�`L�Ӕ�DAU�ՃEA��Ġt����G�Hr��OGBO}O)�WL ?`��� ITV���0\�R;EC�SCRf 0��a�D^�����MARG��`!P�)�T�/ty�$?I�S�H�WW�I�ܩ�T�JGM��MN�CH��I�FNKEuY��K��PRG���UF��P��FWDv��HL�STP���V��@�����RS"S�H�` �Q�C�T1� ZbT�R ���U����@��|R��t�i���G��8PPO��6�F�1�Mޘ�FOCU��RG�EXP�TUI��IЈ�c��n��n ����ePf���!p6�ePr7�N���CANAI��jB��VAIL��C�Lt!;eDCS_H!I�4�.��O�|!"�S Sn�y�0I�BUFF1�XY��PT�$ �� �v��fă�`1�A�rYY��P ���\��pOS1�2��3���_�0Z �  ��aiE�*�.�IDX�dP�RhraO�+��A&ST���R��Yz�<! Y$EK&CK+����Z&m&��1[ L ��o�0��]PL�6pwq��t^����tL6�_ \ ����瀰��7��#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3b�DM�R7��LDR5<4R5ORG.���e2 (`���V�8.��T<�4�d^ �q�<4��-4
R5S�`T00m��0D}FRCLMC!D`�?�?3I@�� MIC���d_ d���RQzm�q�DSTB	��  �Fg�HAX�;b �H�LEXC#ESZr�rBMup�a`��B;d��rB`�j�`a��F_A�J���$[�O�H0K�db� \��ӂS�$MB既LIБ}SREQUIR�R>q�\Á�X�DEBU��DI�+ML� MP�c�ba���P؃ӂ!B0ND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@qܮ�o� �SPS�T8� e�rLO�C�RI�p�EXfA�p��A�AOD�AQP�f X��ON��[rMF�����f )�"I��%�e��T��ѻFX�@IGG� g �q��"E�0�h�#���$R�a%;#�7y��Gx��VvCPi�D'ATAw�pE:�y��[�Eѭ�NVh t_ $MD�qIёA)�v+�tń�tH�`��P�u�|��sANSAW}��t�?�uD��)�r�	@Ði �@CU��V�T0�A�oARR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2��RIN��v�<ZN�NTE���kE�`��,�V�����_N�l��ڂ��kDׄRmn�DIViFDH�@tـn�$V���'c!$��$Z �����~�[���oH �$BE�LTb��!ACCE�L+��ҡ��IR!C�t����T/!���$PS�@#2L  �Ė83������� ��PATH������"��3̒Vp�A_�Q��.�4�B�Cᐈ�_{MGh�$DDQ�<��G�$FWh��p`��m�����b�DE���PPABNԗROTSPEED����00J�Я8��@��̐?$USE_��P��s�SY��c�A- >qYNu@Ag���OFF�q�MOUfN�NGg�K�OL�H�INC*��a��q��Bj�L@�BENCS���q�Bđ���D��IN#"I̒��4�\Bݠ�VEO�w�Ͳ23_�UPE�߳LOWL����00����D����BwP��� �1RC<ʀƶMOSIV�JR�MO���@GPERoCH  �OV� �^��i�<!�ZD<!��c��d@�P��V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�̒<�p1Ӣ`0 ��RTI$Qx�0 MO���МB R �0J��D��s�H�����b�DUM2(�S�_BCKLSH_C̒��>�=�q�#�U���ԑ���2�t�]ACLALvŲ�1n�P�CHK00'%SD�RTY4�k��y�1�q9_6#2�_UM$Pj�9Cw�_�SCL��Ơ�LMT_J1_LDO��@���q��E������๕�幘SP�C��7������PC�o���H� �PU�m�C�/@�"XT_�c�CN�_��N��e���SFu���V�&#����9��̒��=�C�u�SH 6#��c����1�Ѩ�o�`0�͑
��_�PAt�&h�_Ps�W�_10��@4�R�01D�VG�J� 1L�@J�OGW����TORQU��ON *�Mٙ�sRHљ��_W��-�_=��C���I��I�I�II�F�`�JLA.�1[�VC��0�D�BO�1U�@i�B\JR�KU��	@DBL�_SMd�BM%`_sDLC�BGRV�`�C��I��H_8� �*COS+\�(LN�7+X>$C� 9)I�9)u*c,)�1Z2 HƺMY@!�(� "TH&-�)THE{T0�NK23I���"=�A CB6CB=�C�A�B(261C��616SBC�T25GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t��Bȿ6���AQ|r�f$N	E�DpIB U�\B5��$!��!A�%E(G8%(!LPH$U�2׵�2SXpCc%pCr%@�2�&�C�J�&!�VAHQV6H3�YLVhJVuKUV�KV�KV�KV�KV�IHAHZF`RXM��TwXuKH�KH�KH�KUH�KH�IO2LOAH�O�YWNOhJOuKO��KO�KO�KO�KO�&F�2#1ic%�d4G�SPBALANC�E_�!�cLEk0H_�%SP��T&�bc&|�br&PFULC�h`r�grr%Ċ1ky��UTO_?�jT13T2Cy��2N&�v� ϰctw�g�p�0Ӓ~����T��O���� I�NSEGv�!�REqV�v!���DIF�f�1l�w�1m�0�OB�q
����MI�ϰ1��LCHWA�R����AB&u�$MECH,1� :�,@�U�AX:�P��Y�8G$�8pn 
Z���|���ROBR�CR�̒��N�x&�M�SK_�`f�p P+ Np_��R����΄ݡ�1��ҰТ΀�ϳ��΀"�IN�q��MTCOM_C|@j�q  L���p��$NORE�³5���$�r �8� GR�E�SD��0ABF�$XY�Z_DA5A���D�EBU�qI��Q�su �`$�COD��G ��k�F�f��$BUFIND�XР  ��MO�R��t $-�U ��)��r�B��Ӱ���Gؒu � ?$SIMULT ���~�� ���OBJE|�` �ADJUS>��1�AY_Ik��Dp_����C�_FIF�=�T� ��Ұ�� {��p� �����p�@�ŝD�FRI��ӥT&��RO� ��E�{�=͐OPWO�ŀ�v0��SYSByU�@ʐ$SOP�ȸ��#�U"��pPR�UN�I�PA�DpH�D����_OU��=��qn�$}�I�MAG��ˀ�0Pf�qIM����IN��q���RGOVRDȡ:���|�P~���Р�0L_6p���i��SRB���0��M���EDѐF� ��N�`M*���a��˱S�L�`ŀw x �$OVSL�vSDI��DEXm�g�eĐ9w�����V� ~�N ���w����Ûǖȳ�}M�{ ��q|<��� x Hˁ�E�F�ATUS����C�0àǒ��BT�M����If���4p����(�ŀy Dˀ!Ez�g���PE�r��p���
���EXE���V��E�Y�$Ժ ŀz3 @ˁ��UP{�h�3$�p��XN����9�H� �PG�"�{ h $S#UB��c�@_��01�\�MPWAI��PL����LO��<�F�p��$RCVFA�IL_C�f�BW�D"�F���DEFS}Pup | Lˀ�`�D�� U�UN!I��S���R`���_L�pP��̐���ā}��� B�~����|��`ҲN�`KET���y���P� $�~z���0SIZE���ଠ{���S<�OR~��FORMAT/p` � F���rEMR��y�UX������PLI7�ā � $�P_SW�I���͐�_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W �U����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�!O�0\H��6@�@�U�� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�Hӱt@�W�UpS��хDM��O㵐.'}q��Cg@���@ʣ�ߑ�R�M�A�Â� � $P9Y��$WH`'�NGp���H`��Fb��0Fb��Fb��PLM����	� 0h�H�{�X��O���z�Z�eT�M����# pS��C��O@__0_B_�a��_%�� |S����@	�v ��v �@���w�v��9EM��% yR�frJ�B�ː��ftP��PM��QU� ��U�Q��Af�Q�TH=�HOL��Q7HYS�ES�,��UE��B��O#��  ��P0�|�gAQ�(��ʠu���O��ŀ��ɂv�-�A;ӝR#OG��a2D�E��Âv�_�ĀZ�INF�O&��+����b�vR�OI킍 ((@SLEQ/�#� �����o���S`c0QO�0�01EZ0sNUe�_�AUT�Ab�COPY��Ѓ�{��@M��N�����1h�P�
� ��RGI������X_�Pl��$�����`�W��P���j@�G���EX_T_CYCtb����p����h�_N�A�!$�\�<�R�O�`]�� � 9m��POR�ㅣ\���SRVt�)��6��DI �T_l����Ѥ{�ۧ��ۧ �ۧ5*٩6٩7٩8��R�iS�B쐒��$�)F6���PL�A�A^�TAR��@E `��Z�����<��d� �,(@FLq`h��@Y�NL���M�C���GPWRЍ�쐔e�ODELAѰ�Y�p�AD#qX� �QSwKIP�� ĕ�Zx�O�`NT!���P_x���ǚ@�b �p1�1�1Ǹ�?�  �?��>��>�&�>��3�>�9�J2R�;쐖 4��EX� TQ����ށ�Q����[�KFд�8�RD�CIf� �U`�X}�R�#%M!*�0�)�~�$RGEAR_0sIO�TJBFLG�L�igpERa��TC݃�������2TH2N<��� 1�b��uGq T�0 ����M���`Ib����REF�1�� yl�h��ENAB��lcTPE?@���! (ᭀ����Q�#�~��+2 H�W���2�Қ����"�4�F�X�j�3�қ{��������
j�4�Ҝ��
��.�(@�R�j�5�ҝu������������j�6�Ҟ���(:Lj�7�ҟo�����
j�8�Ҡ��"x4Fj�SMSK������a��E�A~��REMOTE������@ "1��Q&�IO�5"%I��P��POWi@쐣  �����X�gpi������Y"$DSB_SIGN4A�Qi�̰�C���tRS232�%�Sb�iDEVI�CEUS#�R�RP�ARIT�!OP�BIT�Q��OWCONTR��Qⱬ��RCU� M�SU_XTASK�3NB���0�$TATU�PK��S@@쐦F��6�_�PC}�$F�REEFROMS8]p�ai�GETN@S��UPDl�ARB��S�P%0���� !>m$USA���a8z9�L�ERI�0f�&�pRY�5~"_�@f�qP�1�!�6WRK�D9�F9ХFR�IEND�Q4bUFx��&�A@TOOLHF�MY5�$LEN�GTH_VT��FCIR�pqC�@�E� �IUFIN�R����RGI�1�AITI:�xGX��I�FG2�7G1a����3��B�GPRR�DA��Oa_� o0e�I1RER�0đ�3&���TC���AQJV�G|�.2���F��1�!d�9Z�8 +5K�+5��E�y�L0�4��X �0m�L
N�T�3Hz��89��%��4�3G��W�0�W�RdD�Z��Tܳ���K�a3d��$cV �2���1��I1TH�02K2sk3K3Jci�aI�i�a�0L��SL��R$Vؠ�B%V�EVk��A bQ*R
��� �,6Lc����9V2F{/P:B��PS_�Et�$rr�C��γ$A0��wPR���v�U�cSk�� {��w�"�1��� 0����VX`�!�tX`���0P�Ё�
�5S^K!� �-qR���!0���z�NJ A)X�!h�A�@LlA��^A�THIC�1��8�����1TFE���q>>�IF_CH�3A�aI0�����G1�x�������9�Ɇ_�JF҇PR(����RVAT�� ��-p��7@����DO��E��COU(��A�XIg��OFFS=E+�TRIG�SK���c���Ѽ�e�[�K�Hxk���8�IGMAo0�A-��ҙ�ORG�_UNEV��� ��S�쐮d ӎ$������GR3OU��ݓTO2��!�ݓDSP��JOG�'��#	�_P'�2O�R���>P6KEPFl�IR�0�PM�R&Q�AP�Q��E�0q�e���SYSG��"��;PG��BRK*Rd�r�3�-�������ߒ�<pAD��ݓJ�BS�OC� N�DU�MMY14�p\@S}V�PDE_OP3�SFSPD_OVR��ٰCO��"��OR-��N�0.�F�r�.��OV�SFc�2�f��F��!4��S��RA�"LCHD}L�RECOV��0�W�@M�յ�#RO3��_�0�� @�ҹ@VER�E�$OFS�@CV� 0BWDG�ѴC���2j�
�TR�!|��E_FDOj��MB_CM��U�B �BL=r0�w�=q�t�VfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�#�8$CA�{Й�>��8$HBK|1c��IO��.�:!aPPA"�N�3�^�F����:"�DVC_DB�C��d�w"����!"��1���ç�3����/ATIO� �q0��UC�&CAB �BS�PⳍP�Ȗ���_0c�SUBCPUq��S�Pa a� ��}0�Sb��c��r"ơ?$HW_C����:c��IcA�A-�l$�UNIT��l��A�TN�f����CYC=LųNECA��[��FLTR_2_F�I���(��}&��LPx&�����_SCT@SF_��F����G����FS|!�¹�CHA�A/����2��RS�D�x"ѡb�r�: _T��PRO��O�� KEM�_��8u�q u�q��D�I�0e�RAILAiC��}RMƐLOԠdC��:anq��wq��V��PR��SLQk�fC�ѷ 	��FUsNCŢ�rRINkP`+a�0 ��!RA� >R 
Я�ԯgWAR�BLFQ���A�����D�A�����LD@m0�aB9��nqBTIvrbؑ���PgRIAQ1�"AFS�P�!�����`%b����M�I1U�D�F_j@��y1°LM�E�FA�@HRDY4�4��Pn@RS@Q�0|"�MULSEj@xf�b�q �X���ȑ���$.A-$�1$c1Ó����� x~�EaGvpݓ�q!AR����09>B�%��wAXE��ROB���W�A4�_�-֣SYЯ��!6��&S�'WR䩐�-1���STR���5�9�E�� !	5B��=QB90��@6������OT�0vo 	$�ARY8��w20���	%�FI���;�$LINK(�H��1�a_63��5�q�2XYZ@"��;�q�3@��1�2J�8{0B�{D0��� CFI��6G`��
�{�_J�p�6��3aOP_O42Y;5�QTBmA"2�BC
�z�DU"�6=6CTURN3�vr��E�1�9�ҍGFL��`���~ �@�5<:7��� 1�?0K�Mc�68Cb�vrb�4�ORQ��X� >8�#op������wq�Upf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W���T υ� ;����QH�!` �ҽ��U�Q�WkeK#keLcXER��	G!E	0��S�dAWaǢ�:D���7!�!AX�rB!{q��1u y-!y�pz�@z �@z6Pz\Pz� z 1v�y�y�+y �;y�Ky�[y�ky��{y��y�q�yDEBU��$�����L�!º2WG`  AB�!�,��SV���� 
w���m���w��� �1���1���A���A�� 6Q��\Q���!�m@�\�2CLAB3B�U������S  �ÐER���� �� $�@� Aؑ!p�PO��Z�q0w��^�_MRAȑ� �d  T�-�EcRR��TYz��B�I�V3@�cΑTOQ�d:`L� �d2��]�X�C[! � p�`T}0i��_V1�r�a'�4��2-�2<����@P�8����F�$W��g�j�V_!�l�$�P�����c��q"�	��SFZN_CFG_!� 4��?º��|�ų����@�ȲW �oV ��\$� �n���Ѵ��9c�Q���(�FA�He�,�XEDM�(�����!s��Q�g�P{RV HE�LLĥ� 5�6�B_BAS!�R�SR��ԣo �#S���[��1r�%��2�ݺ3ݺ4ݺ5ݺ6�ݺ7ݺ8ݷ��ROaOI䰝0�0NLK!ưCAB� ��AC-K��IN��T:�1��@�@ z�m�_PUf!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KA1Rӑ��RE~��qP��(��QUE������P
��CSTOPI_AL�����0�&���㰑�0SEM�l�b�|�M��d�TYf|�SOK�}�DI������(���_TM>\�MANRQ�ֿ0�E+�|�$KEY?SWITCH&	����HE
�BEAiT����E� LEҒ���U��FO�����O_HOM�On�REF�PPRzP��!&0��C+�OA��ECO��B�r�IOCM�D8׵��]���8�` � DH�1����U��&�MHx�»P�CFORC��n� ��OM�  � @V��|�U,3P� 1-�`� �3-�4��NPXw_ASǢ� 0Ȱ�ADD����$S�IZ��$VAR\ݷ TIP]�\�
2�A򻡐���]�H_� �"S꣩!Cΐ���FRIF⢞�S0�"�c���NF��V ܻ�` � x�`SI��TES�R6SSG%L(T�2P&��AxU�� ) STMTQ2ZPm 6BW�P*�SHOWb��S�V�\$�� ���A00P�a�6���@�J�T�5��	6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	 f0u�	�0u�	�@uP[Pu%121?U1L1Y1f1sU2�	2�	2�	2�	U2�	2�	2�	2U22%222?U2L2Y2f2sU3P)3�	3�	3�	U3�	3�	3�	3U33%323?U3L3Y3f3sU4P)4�	4�	4�	U4�	4�	4�	4U44%424?U4L4Y4f4sU5P)5�	5�	5�	U5�	5�	5�	5U55%525?U5L5Y5f5sU6P)6�	6�	6�	U6�	6�	6�	6U66%626?U6L6Y6f6sU7P)7�	7�	7�	U7�	7�	7�	7U77%727?U7,i7Y7Fi7s�?&��VP�UP}D��  ��x|�԰��YSLOǢ� � z��и� ��o�E��`>�^t��А�ALUץ����CU����wFOqID_L��ӿuHI�zI�$FILE_���t�ĳ$`�JvSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_ �TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅�%L~�_Vj�7+p�ޠ�� ` �GR�OU�pD��B�N�FLIC��RE�QUIREa�EB�UA��p����2��������c��{ \��APPR��iC���
�EN��CLOe��S_M� v�,ɣ�
���7� ���MC�&����g�_MG�q�C�� �{�9���|�BRKz�NOL��|ĉ R��_LI|��Ǫ�k�J����P
���ڣ������&���/���6��6��8��Y����� ��8�%��W�2�e�PATH a�z�p�z�=�vӥ�ϰm�x�CN=�CA������p�IN�UCh��bq��CO�UM��!YZ������qE%����2������PAYL�OA��J2L3pR'_AN��<�L��F��B�6�R�{�R_F2�LSHR��|�LO�G��р��ӎ���ACRL_u�������.�r��H�p�$H{�^��FLEX
�s�}J�� :� /����6�2�����;�M�_�F16����n�@��������ȟ��Eҟ �����,�>�P�b� ��d�{�������������5�T��X ��v���EťmF ѯ�������&��/�A�S�e�D�Jx�� � ������j��4pAT����n�EL�  �%øJ���vʰJE��CTR�і��TN��F&��H�AND_VB[�
�pK�� $Fa2{�6� �rSWi��4r�U��� $$Mt�h�R��08�� @<b 35��^6A�p3�k��q{9t�A�̈p��A��A�ˆ0��U���UD��D��P��G���IST��$A��$AN��DYˀ�{�g4�5 D���v�6�v��5缧�^�@��P���Հ�#�,�5�>�
�K�� &0�_�ER!V9��SQASYM��] ������x��ݑ���_SHl�������sT�( ����(�:�JA����S�cir��_VI��#Oh9�``V_UCNI��td�~�J�� �b�E�b��d��d�f ��n���������uN!���2�H����3��"CqEN� �pSDI��>�ObtDќDpx�� ��2IxQA����q��-��s� �� ����� �^�OMME�h�rr/�TVpPT�P  ���qe�i����P��x ��yT�Pj� �$DUMMY9��$PS_��R�Fq�  ��:� ����!~q� XX����K�STs�ʰ�SBR��M21_�Vt�8$SV_E�Rt�O��z���CLRx�A  O�r?p? �Oր � D ?$GLOB���#LO��Յ$�o���P�!SYSADqR�!?p�pTCHM0 � ,����oW_NA��/��e�$%SR��l (:]8:m�K6 �^2m�i7m�w9m��9 ���ǳ��ǳ���ŕߝ �9ŕ���i�L�񝀤�m��_�_�_�TD�XOSCRE�ƀ�� ���STF���}��pТ6�dP] _:v AŁ� T����TYP�r�K��u�!u���O�@I�S�!��tsqUE�{t� ����H�S<���!RSM_�XuUNEXCEPWv��CpS_��{ᦵ�������÷���COUx ��� 1�O��UET�փr���PoROGM� FLn!o$CU��PO*q���c�I_�pH;� �� 8��N�_H�E
p��Q��pRY ?���,�J�*�����?�OUS>�� � @d����$BUTT��R|@���COLUM��<�u�SERVc#=��PANEv Ł� w� �PGEU�!��F��9�)$HE�LP��WRETER��)״���Q�� ����@� P�P� �IN��s�PN(ߠw v�1�����o ���LN�'� ����_��k��$H��M TEX8�#����FLAn +/RELV��D4p��������M��?,@��ӛ$����P=�USRVIEWŁ�� <d��pU�p�0NFIn i�FOsCU��i�PRILP�m+�q��TRI}P)�m�UNjp�{t� QP��XuW�ARNWud�SRT+OLS�ݕ������O|SORN��RA�Uư��T��%��V�I|�zu� =$�PATHg���CACHLOG6�O�LIMybM���x'��"�HOST6��!�r1�R�OgBOT5���IMl�	 D�C� g!��E��L���i�VCPU_�AVAILB�O�EX7�!BQNL�(��`�A�� Q��Q �\�ƀ�  QpC����@$TOOLz6�$�_JMP�� �I�u$S�S�!$��VSHI9F��|s�P�p��6�s���R���OS�URW�pRADIz��2�_�q�h�`g! �q)�LUza�$OUTPUTg_BM��IML��oR6(`)�@TILN<SCO�@Ce� ;��9��F��T�� a��o�>�3���$��w�2u�sqV�zu9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+��t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2$��2���5��`�? tpZA�BCS��  �$�2��J�
���$�$CLAS�����AB��0'@@�VIRT��O.@A�BS�$�1 <E�� < *AtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v���8��M@[�AXLրK��*B�dC  ���IqN��ā��PRE������LAR�MRECOV �<I䂥�NG�� �\K	 A  � J�\�M@PPLIMC�?<E�E��Handl�ingTool ��� 
V7.5�0P/28[�  o�H���
�w_SW�� UP*A7� ��F0ڑ���A�0�� S20��*A���:�ާ��FB �7DA5�� �#'@I�y@��None������� ��T���*A49�+xl�_��V����:g�UTOB���������HGAPO�N8@��LA��U��D� 1<EfA����������� Q 1שI Ԁ��Ԑ�:�i�n��܍�#B)B �3��\�HE�Z��r�HTTHKY ��$BI�[�m����� 	�c�-�?�Q�o�uχ� �ϫϽ��������_� )�;�M�k�q߃ߕߧ� ���������[�%�7� I�g�m������� ������W�!�3�E�c� i�{������������� ��S/A_ew �������O +=[as�� �����K//'/ 9/W/]/o/�/�/�/�/ �/�/�/G??#?5?S? Y?k?}?�?�?�?�?�? �?COOO1OOOUOgO yO�O�O�O�O�O�O?_�	__-_K_Q_��(�T�O4�s���DO_C�LEAN��e��SN�M  9� ��9oKo]ooo�o�D?SPDRYR�_%�HI��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ|��g�PLUGGҠ��Wߣ��PRC�`B�`9��o�=�OxB��oe�SEGF��K������o%o�����#�5�m���LAP �oݎ����������џ �����+�=�O�a�>��TOTAL�.����USENUʀ�׫ �X���R(�RG�_STRING �1��
��M��Sc�
��_�ITEM1 �  nc��.�@�R�d�v� ��������п������*�<�N�`�r��I/O SIGN�AL��Try�out Mode��Inp��Simulated��Out��O�VERR�` = �100�In �cycl���P�rog Abor������Stat�us�	Hear�tbeat��M?H FaulB�K�AlerUم�s߅� �ߩ߻��������� �S���Q�� f�x���������� ����,�>�P�b�t�p������,�WOR�� ����V��
.@ Rdv����� ��*<N`PO��6ц��o �����//'/ 9/K/]/o/�/�/�/�/��/�/�/�/�DEV �*0�?Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�OPALTB��A�� �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_�oo(o:o�OGRI �p��ra�OLo�o�o�o �o�o�o*<N `r������`o��RB���o�>� P�b�t���������Ώ �����(�:�L�^�xp����PREG�N ��.��������*� <�N�`�r����������̯ޯ���&�����$ARG_��D �?	���i���  w	$��	[}��]}���Ǟ�\�SB�N_CONFIG� i��������CII_SAV/E  ��۱Ҳ�\�TCELLSE�TUP i�%�HOME_IO��͈�%MOV_8�2�8�REP����V�UTOBACK�
�ƽF�RA:\�� X�Ϩ���'` ���x������ �� ��$�6�c�Z�lߙ���������������� �!凞��M�_�q�� ���2��������� %�7���[�m������ ��@�������!3E$���Jo��p�����INI�@���ε��MESSAG����q�>�ODE_D$��ĳ�O,0.��PA�US�!�i� ((Ol���� ���� /�// $/Z/H/~/l/�/�'a~kTSK  qx�����UPDT%��d0;WSM�_CF°i��еU�'1GRP 2�h�93 |�B��A|�/S�XSCRD+1;1
1; ����/�?�?�? OO$O ��߳?lO~O�O�O�O �O1O�OUO_ _2_D_�V_h_�O	_X���GR�OUN0O�SUP�_NAL�h�	ܢĠV_ED� 1�1;
 �%-B?CKEDT-�_`�!oEo$���a�o�����ߨ���e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[8�5GED4�n�#�� ~�j���ED5Z��Ǐ6� ~��8�}���ED6�����k�ڏ ~G���!�3�ED7��Z��~� ~�8V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W�Ư�
}3�����CR o�����3�տ@ϯ�����P�PNO_DE�L�_�RGE_UN�USE�_�TLAL_OUT q��c�QWD_ABO�R� �΢Q��ITR�_RTN����N'ONSe����CAM_PARA�M 1�U3
 �8
SONY �XC-56 234567890�H� � @����?���( Щ�V�|[r؀~�X�HR5k�|U�Q��ο�R57����A�ff��KOWA SC310M|[�r�̀�d @6�|V��_�Xϸ� ��V��� ���$�6���Z�l��CE_RIWA_I857ЍF�1��R|].��_LIO4W=� ���P<~�F<�GwP 1�,����_GYk*C*�  ��C1� 9J� @� G� �CL�C]� d� l� s��R� ��[�m�� v� � �� ��� C�� �"��|W��7�HEӰON�FI� ��<G_P_RI 1�+P� m®/���������'CHKPAU�S�  1E� ,�>/P/:/t/^/�/ �/�/�/�/�/�/?(?@?L?6?\?�?"O������H�1_MO�R�� �XaB�iq-���5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`��S:�(�����U�p�_)o�S  %�3Pq���R�P�_�mo8j�����Oko�o9i�(�=�(�>Okg�o�o�l�Kof�oGq:I�Z?DEF f8���)�R6pbuf.txtm�]n�@��Y��# 	`(Ж�Ao=L���zMC�21�=a� :���4��=�n׾�Cz � BHBCCPUe�B�_B�y�;��>C����CnaSWE@E?�{hD]^Dٿ�?r����D���^��G	���F��F���Cm	fF�O�OF�ΫSY���vJqG���Em�(�%.���1(��<�qѦG�x2��Ң �̢ a�D�j���E�S\��X�EQ��EJP F�E��F� G����F^F E��� FB� H,�- Ge��H3�Y����`�33� ���xV  in2xQ@��5Y���8B� A�AST<#�
� �_'�%��w�RSMOFS��،~2�yT1�0DEg �O@b 
�v(�;�"�  <�6�z�R���?�j�CC4��aSWm� W�Q�{�m�C��B-JG�Cu�@$�q���T{�FPROG C%i����c�I���� �Ɯ�f�KEY_�TBL  �vM��u� �	
��� !"#$%&�'()*+,-.�/01c�:;<=�>?@ABC�pG�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������p���͓���������������������������������耇����������������������!j�LC�K��.�j���STA�T���_AUTO�_DO���W/�INDT_ENB�b�2R��9�+�T2wߞXSTOP\߿2T{RLl�LETE�����_SCREE�N ik�csc��U��MM�ENU 1 i  <g\��L� SU+�U��p3g���� ���������2�	�� A�z�Q�c��������� ������.d; M�q����� �N%7]� m���/�� /J/!/3/�/W/i/�/ �/�/�/�/�/�/4?? ?j?A?S?y?�?�?�? �?�?�?O�?O-OfO =OOO�OsO�O�O�O�O��O_�O_P_Sy�_?MANUAL��n��DBCOU�RIG|���DBNUM�p���<���
�QPXWORK 1!R�ү�_oO.o@oRk��Q_AWAY�S^��GCP ��=��df_AL�P�db�R�Y�������X_�p �1"�� , 
�^���o xvf`%MT�I^�rl@�:s�ONTIM���&���Zv�i
õ�cMOTNEND����dRECORD �1(R�a��ua�O��q��sb�.� @�R��xZ������� ɏۏ폄���#���G� ��k�}�����<�ş4� �X���1�C���g� ֟��������ӯ�T� 	�x�-���Q�c�u��� �������>���� )Ϙ�Mϼ�F�࿕ϧ� ����:�������%�s` Pn&�]�o��ϓ�~ߌ� ��8�J�����5� � ��k����ߡ��J��� ��X��|��C�U��� �������0������	��dbTOLER7ENCqdBȺb`�L�͐PCS_C�FG )�k)wd�MC:\O L�%04d.CSVd
�`c�)sA �+CH� z�`)~����hMRC_O_UT *�[�n~SGN +�e��r��#�10-�MAY-20 1�0:46*V15-�JANj51�k? P/Vt���)~�`pa�m��PJPѬ�VERSION� SV2�.0.8.|EFLOGIC 1,�[/ 	DX�P7)��PF."PROG_�ENB�o�rj UL�Sew �T�"_WRSTJNEp�V�r�`dEMO_OPT?_SL ?	�es�
 	R575)s7)�/??*?<?|'�$TO  �-د�?&V_@pEX�Wd�u�3PAT�H ASA\p�?�?O/{ICT�a-Fo`-�gds�egM%&ASTBF_TTS�x@�Y^C��SqqF�P�MAU� t/XrMS%WR.�i�a.|
S/�Z!D_N�O0_�_T_C_x_g_�_�tSBL_FAUL"y0�[3wTDIAU �16M�ap�A�1234567G890gFP? BoTofoxo�o�o�o�o �o�o�o,>Phb�S�pP�_ ���_s�� 0`�� ���)�;�M�_�q� ��������ˏݏ��|�)UMP�!� �^�TR�B�#+�=��PMEfEI�Y_T�EMP9 È�3p@�3A v�UNI�.�(YN_BRK �2Y)EMGDI_STA�%WЕ�NC2_SCR 3��1o"�4�F� X�fv���������#��ޑ14�����)�;�����ݤ5�����x�f	u�ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/߭P�b�t� � ��xߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N���r����� ����������& 8J\n���� ����"`�F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ 4?,?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�O �O�O?�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�O�O�o�o �o
.@Rdv �������� �*�<�N�`�r����o ����̏ޏ����&� 8�J�\�n����������ȟڟ����H�ETMODE 16���� ���ƨ
R�d�v�נRR�OR_PROG �%A�%�:߽� � ��TABLE  A������#��L�RRSEV_N�UM  ��Q���K�S���_A�UTO_ENB � ��I�Ϥ_NONh� 7A�{�R�_  *������%������^�+��Ŀ8ֿ迄�HISO�͡�I�}�_ALM 1]8A� �;�����+�e�wωϛ�ȭϿ��_H���  �A���|��4�T�CP_VER �!A�!����$EX�TLOG_REQ���{�V�SIZ�_�Q�TOL  �͡Dz��A Q�_BWD����r����n�_DI�� 9��}�z�͡m���STEP����4���OP_DO����ѠFACTOR_Y_TUN�dG��EATURE �:����l��Handling�Tool ��  �- CEng�lish Dictionary���ORDEAA� Vis�� Ma�ster���96� H��nalog� I/O���H5�51��uto S�oftware �Update  ���J��matic Backup��Part&�g�round Ed�it��  8\a�pCamer�a��F��t\j6�R�ell���LO�ADR�omm��syhq��TI" ���co��
! o����pane�� �
!��tyl�e select.��H59��nD���onitor��4�8����tr��Re�liab���ad�inDiagnos"����2�2 �ual Chec�k Safety� UIF lg\�a��hanced� Rob Ser}v q ct\���lUser Fr�U��DIF��Ext. DIO ��fiA d��e�ndr Err L,@��IF�r�� � �П�90��FCTN MenuZ �v'��74� TPw In��fac�  SU (�G=�p��k Ex�cn g�3��Hi�gh-Sper S�ki+�  sO�H�9 � mmunic�!�onsg�teu�r� ����V�����conn��2���EN��Incr�stru���5�.fdKAR�EL Cmd. ML?uaA� O��Run-Ti� E�nv����K� ��+�%�s#�S/W��7�4��Licens�eT�  (Au�* ogBook(�Sy��m)��"�
MACRO�s,V/Offsme��ap��MH� ܷ���pfa5�Me�chStop Pgrot��� d�zb i�Shif��^��j545�!xr x��#��,K�b �ode Swit�ch��m\e�!o�4.�& pro��4��g��Multi-T7G���net.Po=s Regi��z��P��t Fun����3 Rz1��NCumx �����9m�|�1�  Adjuj���1 J7�7�* x����6tatuq1�EIKRDM�tot��scove�� ��@By- �}uest1�$Go�� � U5\SNPX b"���YA�"Libr���Ŀ#�� �$~@h�pd�]0�Jts in VCCM�����0��  �u!��2 RL�0�/I�08��TMILIB�M �J92�@P�Ac�c>�F�97�TP�TX�+�BRSQe9lZ0�M8 Rm���q%��692��Un�exceptr m�otnT  CV1V�P���KC������+-��~K  II�)�VSP CSXC�&.c�� e�"��{ t�@WewΌAD Q�8bvr� nmen�@�i%P� a0y�0�pf�GridAplay !� nh�@*�3R��1M-10iA(_B201 �`2V"�  F���scii��load��83� M��l����Gu{ar�d J85�0��mP'�L`���st�uaPat�&]$Cyqc���|0ori_ �x%Data'Pqu���ch�1��g`ڂ j� RLJam��5���IMI D�e-B(\A�cP" �#^0C  et�kc^0asswo\%q�)650�Ap�U�Xnt��Pve�n�CTqH�5�0�YELLOW �BO?Y��� Arc�0vis��Ch��WeldQciail4Izt�Op� X��gs�` 2@�a��poG yRjT11 NE�#HT� 3xyWb��! �pB�`gd`���p\� =P���JPN ARC�P*PR�A�� wOL�pSup̂fil�p��J�� ��7cro�670�1CX~E�d��SS�pe��tex�$ �P� S�o7 t� ssagN5 <Q�BP:� �9 "0�QrtQC��9P�l0dpn�笔��rpf�q�e�ppm�ascbin4�psyn�' pt�x]08�HELN�CL VIS P�KGS �Z@MBq &��B J8@�IPE GET_�VAR FI?S �(Uni� LU�OOL: ADD�@_29.FD�TCm���E�@DVp���`�A�ТNO WTW�TEST �� Vx�!��c�FOR �ЯECT �a!� ALSE ALA`��CPMO-130���� b D: HANG FROMg���2��R709 �DRAM AVA�ILCHECKS� 549��m�VP�CS SU֐LI/MCHK��P�0x��FF POS� F��� q8-1�2 CHARS�E}R6�OGRA ���Z@AVEH�AME���.SV��Вאn�$��9�m "y�T�RCv� SHAD~P�UPDAT k�}0��STATI�~�� MUCH ����TIMQ MO?TN-003���@OBOGUIDE DAUGH��p�b��@$tou� �@C� �0��PAT�H�_�MOVET��� R64��VM�XPACK MA�Y ASSERT�jS��CYCL`�T�A��BE CORg 71�1-�AN���RC OPTIO�NS  �`��AP�SH-1�`fix��2�SO��B��XO�����_T��	�i��0�j��du�byz p� wa��y�٠HI�������U�pb XS�PD TB/�F� /\hchΤB0����END�CE�06\�Q�p{ smay� n@�pk��L >��traff#�	�� ��~1from� sysvar scr�0R� ��d�'DJU���H�!A���/��SET E#RR�D�P7�����NDANT SC�REEN UNR?EA VM �PD�MD��PA���R�?IO JNN�0��FI��B��GRO;UNנD Y�Т�٠�h�SVIP �53 QS��DIGIT VERS���ká�NEW�� P�06�@C�1IMA�G�ͱ���8� D�I`���pSSUE��5��EPLAN {JON� DEL����157QאD��CALLI���Q��m�ޥ�IPND}�IM�G N9 PZ�1�9��MNT/��EsS ���`LocR �Hol߀=��2�PnN� PG:��=�M���can����С:� 3D mE2vi?ew d X���ea1 �0b�pof� Ǡ"HCɰ�A�NNOT ACC�ESS M cp�ie$Et.Qs a�� loMdFlex�)a:��w$qmo G�sA9�-'p~0���h0pa��eJ A�UTO-�0��!i�pu@Т<ᡠIAB�LE+� 7�a FP�LN: L�pl� m� MD<�VI��и�WIT HO�C�Jo~1Qui���"��N��USB��@�Pt & re�mov���D�vAx?is FT_7�P�GɰCP:�OS�-144 � h �s 268QՐOS�T�p  CRASoH DU��$P���WORD.$�L�OGIN�P��P:�	�0�046 is�sueE�H�: �Slow st
�c�`6����໰�IF�IMPR��S?POT:Wh4����N1STY��0VM�GR�b�N�CATZ��4oRRE�� N� 58�1��:%�'RTU!Pe -M a�SE:�@pp���A�GpL��m@acll��*0a�OCB� WA���"3 C�NT0 T9DWr}oO0alarm�ˀm0d t�M�"0��2|� o�Z@OM�E<�� ��E%  #�1-�SRE��M�s�t}0g    } 5KANJI5?no MNS@��INISITAL�IZ'� E�f�w�e��6@� dr�@ �fp "��SCI�I L�afail�s w��SYS�TE[�i��  �� Mq�1QGro8�m n�@vA�����&��n�0q��RW{RI OF Lk�>�� \ref"�
��up� de-re�la�Qd 03.��0SSchőbe�twe4�IND �ex ɰTPa�D�O� l� �ɰG�igE�soper�abil`p l,�HcB��@]�le<�Q0cflxz������OS {����v�4pfigi GLA��$�c2�7H� l�ap�0ASB� I�f��g�2 l\c��0�/�E�� EOXCE 㰁�P��H�i�� o0��Gd`�]Ц�fq�l lx9t��EFal��#�0�i�O�Y�n�CLO�S��SRNq1NT
^�F�U��FqKP�A?NIO V7/ॠ�1�{����DB ��0��ᴥ�ED��DSET|�'� �bF��NLINEb�BU�G�T���C"RLI�B��A��ABC �JARKY@��� orkey�`IL����PR��N��ITGAR� D$�R �Er *�T��a�U�0x��h�[�ZE V�� TASK p.vr�P2" .�Xf�J�srn�S谥dIcBP	c���B/��wBUS��UNN�A j0-�{��cR'�v��LOE�DIVS�CULs$cb����BW!��R~�W`P�L����IT(঱tʠ��OF��UNEXHڠ+���p�FtE���SVEMG3`NM_L 505� D*�CC_SAFE�P�*� �ꐺ� PETp��'P�`�F  !�F��IR����c i �S>� K��K�H GUNCHG���S�MECH��M$��T*�%p6u��t�PORY LEA�K�J���SPExgD��2V 74\�GRI��Q�g��C7TLN��TRe @��_�p ���EN'�IN������$���r��sT3)�i�STO�IA�s�L��͐X	����q��Y� ��T!O2�J m��0F<�K�L���DU�S��O��I3 9�J F��&���SSVGN-q1#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRK�CTR/"� �q\j�5��_�Q�S�qIN=VJ0D ZO�Pݲ ���s��г�Ui ɰ̒��a�DUAL� �J50e�x�RVO_117 AW�TH!pHr%�N�247%��52��|�&aol @���R���at�Sd�cqU���P,�LER���iԗQ0�ؖ  ST����Md�Rǰt� /\fosB�A�0Np��c����{�U��ROOP 2�b�pB��ITP4M��b� !AUt c0< � p�lete�N@�� z1^qR635 �(AccuCal�2kA���I) "P�ǰ�1a\�Ps�� ǐ� bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etacea��AT���PC�`������_p�.p�c!Ɗ��:�cir1cB���5�tl��B���:�fm+�Ί�V��b�ɦ�r�upfr�m.����ⴊ�xepd��Ί�~�pedA��D �}b�ptliabB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̈�Ϙ���c�Ӳ�5�j>�����tcȐ��	�Qr����mm 1��FT�sl^0��T�m�L��#�rm3��ub �Y�q�std}��pl;�&�ckv�=�r��vf�䊰��9�vi����ul�`�0fp��q �.f��� �daq; i Dat�a Acquisi��n�
��T`���1�89��2�2 DMCM R�RS2Z�75��~9 3 R710�o59p5\?���T "��1 (D�T� nk@���������E Ƒȵ��Ӹ�egtdmm ��ER�����gE��1�q\mo?۳�=(G����[(

�2�` !� �@JMACR�O��Skip/Offse:�a��V��4o9� &qR66!2���s�H�
 E6Bq8����9Z��43 J77� 6�J783�o ���n�"v�R5I�KCBq2 PTL�C�Zg R�3 (�s, �������03�	зJԷ�\sfmnmc "MNMC����ҹ��%mnf�FMC�"Ѻ0ª etmc�r� �8����� ,K�DV��   87?4\prdq>,�jF0���axis�HProcess� Axes e�r;ol^PRA
�Dp~� 56 J81j�[59� 56o6� ئ��0w�690 98� [!IDV�1��2q(x2��2ont�0 �
����m2���?�C��etis "�ISD��9�� FpraxRAM�P� D��defB�,�G��isbasic�HB�@޲{6�� 7�08�6��(�Ac w:������D
�/,��AMOX�� ��DvE���?;T��>Pi� RAF!M';�]�!PAM�V �W�Ee�U�Q'
bU��75�.�ceNe�� nterfac�e^�1' 5&!54x�K��b(Devam ±�/�#���/<�Ta=ne`"DNEWE����btpdnui �AI�_s2�d_r�sono���bAsf�jN��bdv_ar�Fvf�xhpz�}w��h9kH9xstc��g�AponlGzv{�ff��r���z��3{q'Td>pch'ampr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�~!�pcchmp]a�MP&B�� �mp�ev�����pc�s��YeS�� Ma�cro�OD��16 Q!)*�:$�2U"_,��<Y�(PC ��$_�;������o��J�ge�gemQ@GEMS�W�~ZG�gesndxy��OD�ndda���S��syT�Kɓ�s!u^Ҋ���n�m���L���  ���9:p�'ѳ޲��spotplusp���`-�(W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\fewatu 0FEAWD��oolo�srAn'!2 p���a�A�s3��tT.� (N. A.)��!eP!�J# (j�,��0�oBIB�oD -�.�mn��k9�"K���u[-�_���p� "�PSEqW����wop "sEЅ�&� :�J������y�|��O 8��5��Rɺ���ɰ [��X�������%�@(
ҭ�q HL�0 k�
�z�a!�B�Q�"(g�Q�����]� '�.�����&���<�!��_�#��tpJ�H�~Z ��j�����y������ �2��e������Z���� V��!%���=�]�͂���^2�@iRV� o%n�QYq͋JF0� !8ހ�`�	(^�dQueue���X\1��ʖ`�+F1tpvt�sn��N&��ftp:J0v �RDV�	f�H�J1 Q���v��en��kvstk✐mp��btkc�lrq���get����r��`�kack�XZ�sctrŬ�%�stl��~Z�np:!�`�@��q/�ڡ6!l�/HYr�mc�N+v3��_� ����.v��/\jF��� ��`Q�΋ܒ�N50 (FRA��+��͢fraparm���Ҁ�} 6�J64�3p:V�ELSE�
#�VAR $S�GSYSCFG.�$�`_UNITS 2�DG~°@�4Jg�fr��4A�@FRL -��0ͅ�3ې���L �0NE�:�=�?@�8�v�9~Qx304��;�BPRSM~QA�5�TX.$VNUM�_OL��5��DJ5�07��l� Functʂ"qwAP��琎��3 H�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TPP�R���QA�prn�aSV�ZS��AS8Dj�510U�-�`cr �`8 ��ʇ�DJR`jY�ȑH  ژQ �PJ6�a21���48AAVgM 5�Q�b0 lBު`TUP xb�J545 `b�`6�16���0VC�AM 9�CL�IO b1�59 ���`MSC8�
r�P R`\sS�TYL MNIN��`J628Q  ��`NREd�;@�`S�CH ��9pDCS�U Mete�`O�RSR Ԃ�a04� kREIOCu �a5�`542�b9vpP<�nP�a�`�R��`7�`�MA�SK Ho�.r7y �2�`OCO :��r3��p�b�p���r�0X��a�`13\m�n�a39 HRM�"�q�q��LC�HK�uOPLG \B��a03 �q.�pOHCR Ob�pCp�Posi�`fP6 {is[rJ554��N�pDSW�bM�D�p�qR�a37 }Rjr0� �1�s4 �R6�76��52�r5 �2�r�7 1� P6���R_egi�@T�u/FRDM�uSaq%��4�`930�uSN{BA�uSHLB̀�\sf"pM�NP�I�SPVC�J�520��TC�`"{MNрTMIL�{IFV�PAC W��pTPTXp6.�%�TELN N �Me�09m3�UECK�b�`UFyR�`��VCOR���VIPLpq89qSsXC�S�`VVF��J�TP �q��R6�26l�u S�`G�ސ�2IGUI\�C��PGSt�\ŀH863�S�q����ւq34sŁ68�4���a�@b>�3 �:B��1 T��96u .�+E�51 yf�q53�3�b1 ��f�b1 n�jr9 ��`VAT ߲�q7�5 s�F��`�sAW�SM��`TOP �u�ŀR52p���a8s0 
�ށXY q�澢0 ,b�`885�QXрOLp}�"p�E࠱tp�`LCM<D��ETSS����6 �V�CPE 9oZ1�VRCd3
��NLH�h��001m2Ep��3 f��p��4 /165C���6l���7PR��0�08 tB��9 -�200�`U0�pFL�1޲1 ��޲2L"����p��޲4��5� \hmp޲6 RBCF�`ళ�fsః8 �Ҋ��~�J�7� rbcfA�L�8`\PC����"�32m0�u�n�K�Rٰn�5 �5EW
n�9 �z��40 kB��3� ��6ݲ�`00iKB/��6�u��7�u���8 µ������sU�0�`�t �1 05w\rb��2 E� ��K���j���5˰���60��a�HУ`:�6�3�jAF�_���F�7 ڱ݀H�8�eHЋ��c�U0��7�p��1�u��8u��9 713������D7� �ҹ5t�97 ��8�U�1��2��1�1:���h��1np�"���8(�U1��\py�l��,࿱v ��B�8�54��1V���D�4��im��1�<��H�>br�3pr�4@pGPr�6 B���цp���1����1�`͵1{55ض157 �2��62�S����!1b��2����1Π"��2���B6`�1�<c�4 7B�5 �DR��8_�B/��1�87 uJ�8 0�6�90 rBn�1� (��202 0EW,ѱ2^��2��90�U2�p�2��2� b��4��2�a"�RB����9\�U2�`w�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`6ڰR,:7 �2��V�2��5���2^��$a^9���qr����n�5����5᥁"��8a�Ɂ}�5B���5����`UA���� ��Y86 �6 S�0���5�p�2�#�529A �2^�b1P�5~�2`���&P5��8��5��u�!ѹ5��ٵ544��5��R�ąP nB^z�c (�4������U5J�V�5��1��1^��%�����5 b21��gA���58W82� rbr��5N�E�5890tr� 1�95 �" ������c8"a��|�PL ���!J"5|6��D^!�6��B�"8�`#��+�8%�6B�AyME�"1 iC��'622�Bu�6V��dڸ 4��84�`AN�RSP�e/S� C�5� �6� ��� �\� �6� �V� 3t~��� T20CA�R��8� Hf� 1DH��� AOE� ��� ,K|�� ��0\�� �!64K���ԓrA� �1 (M-=7�!/50T�[PM��P�Th:1�C�@#Pe� �3�0� 5`M75T"� �D8pC� �0Gc� u�4��>i1-710i�1� �Skd�7j�?6�:-HS,� �RN�@�U�B�f�X�=m75!sA*A6an���!/C,B�B2.6A �0;A �CIB�A�2�QF1�UBu2�21� /70�S� �4����Aj1�3�p���r#0 B2\	m*A@C��;bi"i1�K�u"A~AAU� imm7c7��ZA@I$�@�Df�A�D5*A�EF� 0TkdR1�35Q1@�"*�@�Q�1�QC)P �1*A�5*A�EA�5B,�4>\77
B7=Q�D��2�Q$B�E7�C�D/qAHEE�W7�_|`j�z@� 2�0�Ejc7P�`�E"l7�@7�A 
1�E�V~`�W2%Q�R�9ї@0L_�#�@���"A���b��H3s=rA/2�R5nR4��74rNUQ1ZU�A�s\;m9
1M92L2�!�F!^Y�ps� 2ci��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHs�XBSt62�q`s������ ��Pxq350_*A3I)�2�d�u�0�@� '4TX�06�pa3i1A3sQ�25�c��st�r�VR1%e�q0
��j1� �O2 �A�UEiy�.� ‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ ��qA!Pvs� 5	15 aU���?PŅ���ဎ�Q9A6�zS*�7��qb5�1����Q��00P(��V7]u�ait E1���ïp?7� !?��z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ��y�00\ry�"R2�BL�tN  ��� �1DV� �2�qeR�5����_b�3�X]1m1lcBqP1�a�E�Q� 5F�䥒�!5���@M-16Q�� f���r��Q��e� ��� PN�LT�_�1��i1��9453���@�e�|�b1l >F1u*AY2�
��R�8�Q����RJ�J3�D}T� 85
Qg�/0 ��*A!P�*A�Ð𫿲��2ǿپ6t�6�=Q���Pȓ��� AQ� g�*ASt]1^u �ajrI�B����~�|0I�b��yI�\m�Qb�I�uz�A�c3Apa9q.� B6S��S��m����}�85`N�N�  �(M���f 1���6����161��55�s`�SC��U���A����5\setg06c����10�Fy�h8��a6��6��<9r�2HS ���Er���W@}�a��I�lB@���Y�ٖ�m�u� C����5�B��B��h`�F���X0���A:���C�M��AZ��@��4�6i����� e�O�-	���f1��F ��ᱦ�1F�Y	���T#6HL3��U66~`����U�dU�9D20L f0��Qv� ��fjq�� N������0v
� ��pi	�	��72lqQ�2������� \c�hngmove.�V��d���@2l_arf	�f~ ��6������9C�Z�`��~���kr41 S ���0��V��t���p���U�p7nuqQ`%�A]��V�1\�Qn�BJ�2W��EM!5���)�#:�6q4��F�e50S� \��0�=�PV���e ������E����޵�m7shqQSH"U��)��9�!A��(����� ,�K��ॲTR1�!��,�60e=�4�F�����2��	 R- ������������ ���4���LSR�)"�!lOA��Q�) ,%!� 16�
U/� �2�"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D ���5V��@2cVE֐�p��T��pt갖�1AL~E�#�F�Q��9E��#De/��RT��59 ���	�A�EiR������9\m20�2A0��+�-u�19r4�` �E1�=`O9`�1"ae��O�2��_$W.}am41�4�3�/~d1c_std��1)�!�`_T��r�_? 4\jdg�a�q �PJ%!~`-�r�+bpgB��#c300�"Y�5j�QpQb1�bq0��vB��v25�U��8����qm43� �Q <W�"PsA��e� ���t�i�P�W.� �c�FX.�e�k�E14�44�~67\j4�443sj<��r�j4up���\E19�h�PA�T�=:o �APf��coWo!\��2a��2A;_2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a:8�8J9X�l5�m1�a첚��*���(85 �&�������P6���R,52&A����q,fA9IfI50\u�z�OV
�v��}E֖aJ���Y>� 16r@�C�Y��;��1��L�� �Aq�&ŦP1��vB)�e�m�����1p�] �1DV��27��F�KAREL U�se S��FCTyN��� J97�FA+�� (�Q޵�p�%�)?�Vj9F?(�j��Rtk208 "!Km�6Q�y�j��iÄ�Pr�9�s#��v�kwrcfp�RCFt3����Q��kcctme�!ME�g����6�main�dV�� ���ru��kDº�c`���o����J�dt�rF �»�.vrT�f�����E%�!��5�.FRj73B�K����UER�HJ�O  JF�� (ڳF���F�q �Y�&T��p�F�z��19�tkvBr���V�h�!9p�E�y�<�k�������;�v���"CT ��f����)�
І�� )�V	�6���!��q FF��1q���=����ҀO�?�$"���$��j�e���TCP Au�t�r�<520 H�5�J53E193Z��9��96�!8��q9��	 �B574��52�Je�(�� Se%!Y�����u��m|a�Pqtool����������con�rel�Ftrol� Reliabl�e�RmvCU!��H5�1����� a5�51e"�CNRE¹I�c�&��i�t�l\sfutst "UTա��"X�\u��g@�i�6Q"]V0�B,Eѝ6A� �Q�)C���X��Y�f�I�1|6s@6i��T6IU��vR�d��
$e%1��2�C58�E6��8�Pv�iV4OFFH58SOeJ� mvB7M6E~O58�I�0 �E�#+@�&�F�0�� �F�P6a���)/++�|</N)0\tr1��<���P ,K�ɶ�r�maski�mskH�aA���ky'd�h	A�	�P�sDispl/ayIm�`v����?J887 ("A���+HeůצprdsP��Iϩǅ�h�0pl�E2�R2��:�Gt�@��PRD�TɈ�r�C��@Fm��D�Q�Asc	aҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@<�P�firmQ��ǀ�Pp�2�=bk�6�r�3x��6��tppl���PL���O�p<b�ac �q	��g1J�U�d�J��gait_9e���Y�&��Q���	�Sh�ap��erati�on�0��R67�451j9(`sGe�n�ms�42-f��r��p�5����2�rsg�l�E��p�G���qF�205p�5S���Ձ�r'etsap�BP�O��\s� "GCR��ö? �qngda��G��V��st2a�xU��Aa]��ba�d�_�btput�l/�&�e���tplcibB_��=�2.��8��5���cird�v��slp��x�hex���v�re?�Ɵx�k3ey�v�pm���x�us$�6�gcr���F������[�q27j�92�v�ollismqSk�9O�ݝ� (pl.���t��	p!o��29$Fo8���cg7no@�tptc;ls` CLS�o�b��\�km�ai_
�s>�v�o	�t�b����<��E�H��6�1�enu501�[m���utia|$ca�lmaUR��Cal�MateT;R51%�i=1]@-��/V� �@�Z�� �fq1�9 "K9E�L����2=m�CLMTq�S#f��et �LM3�!} �F�c�nspxQ�c���c_moq��� ��c_e�����#su��ޏ �_ �@�<5�G�join�i� j��oX���&cWv	� ���N�ve��C�c�lm�&Ao# �|$f�inde�0�STD ter �FiLANG4���R��
��n3���z0Cen���r,������J�����  ���K��Ú�=����_Ӛ��r� "F�NDR�� 3��f>��tguid�䙃0N�."��J�tq�� � ������������J����_������c��	�m�Z��\fnd�r.��n#>
B2p|��Z�CP Ma�����38A��� c��6� (���N�B������ 2�$�8�1��m_���"e x�z5�.Ӛ��c��`�bSа�efQ�p��	��RBT;�?OPTN �+# Q�*$�r*$��*$r*$ %/s#C�d/.,P�/0*>ʲDPN��$،��$*�Gr�$k �Exc�'IF�$M�ASK�%93 H�5�%H558�$5/48 H�$4-1�$���#1(�$�0 E��$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9�j0"M�49�4  ��4�4tps�h���4�P�4- DQ� �3�Q�4�R�4�p�R%0�2�r�4.b
E\����5�A�4��3ad�q\�5K979"�:E�ajO l "DAQ^E^�3i�Dq �H�4ҲO ?R�? ���q�5��T��3rAq��O�Lst�5~��7p��5��REJ#�2�@av@^Eͱ�F���4��.�5�y N� �2il(�in�4��31 J0H1�2Q4�251ݠ�4Ormal� �3)� REo�Z_�æOx����4p��^F�?onorTf ��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱH�4�REM���4yݱx"u@�RER5932f�O��47Z��5lit�y,�U��e"Di#l\�5��o ��7�987�?�25 �3hk910�3��FE��0=0P_�Hl\mhm�5��qe�=$�^��
E��u�IAymp�tm�U��BU��vste�y\�3��me�b� DvI�[�Qu�:F�Ub�`*_�
E,�su��_ Er��ox�<��4huse�E-�?�sn�������FE���,�box�����c ݌,"�������z���M��g��pdspw)�	��9���b���(��1���c ��Y�R�� �>�P����W��������'�0�ɵ�[��͂���  � ,K@�� �A�bWumpšf��B*��Box%��7Aǰ6�0�BBw���MC� (�6�,f�t I�s� ST��*��}B������w��"BBF
�>�`���)���\bbk968 a"�4�ω�bb��9va69����et�bŠ��X�����ed	�F��u�f� �sea"������'�\��,���b�ѽՑo6�H�
�x�$�f����!y���Q[�! �tperr�fd�� TPl0o� Recov,��3D��_R642 � 0��LC@}s� N@��(U�'rro���yu2r���  �
�  ����$$C�Le� ���t���������$z�?_DIGIT��������.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_� oo$j��+c:P�RODUCTM�0\PGSTKD��qV&ohozf99���D���$FE�AT_INDEX���xd���  
�`ILECOMP ;����#��`�cSETUP2 <�e��b�  N� �a�c_AP2B�CK 1=�i � �)wh0?{%&c����Q�xe %�I�m��� 8��\�n����!��� ȏW��{��"���F� Տj���w���/�ğS� ��������B�T�� x������=�үa��� ���,���P�߯t��� ���9�ο�o�ϓ� (�:�ɿ^���Ϗ� ��G���k� �ߡ�6� ��Z�l��ϐ�ߴ��� U���y����D��� h��ߌ��-���Q��� ������@�R���v� ���)�����_����� *��N��r� �7��m�&��3\�i
pP� 2#p*.VRc�*��0� /��PC/1/>FR6:/].��/+T�`�/�/�F%�/�,�`r/?�G*.F�8?	H#�&?e<�/�?;STM �2�?�.K �?�=�iPend�ant Pane	l�?;H�?@O�7.Op�?y?�O:GIF�O��O�5�OoO�O_:JPG _J_�56_�O_��_�	PANELO1.DT�_�0 �_�_�?O�_2�_So@�WAo�_o�o�Z3qo��o�W�o�o�o)�Z4 �o[�WI���
TPEINS.�XML��0\����qCusto�m Toolba�r	��PASS�WORDyF�RS:\L�� %�Passwor�d Config ���֏e�Ϗ�B0� ��T�f���������� O��s������>�͟ b��[���'���K�� 򯁯���:�L�ۯp� ����#�5�ʿY��}� �$ϳ�H�׿l�~�� ��1�����g��ϋ� � ����V���z�	�s߰� ?���c���
��.�� R�d��߈���;�M� ��q������<���`� �����%���I����� ���8����n�� �!��W�{ "�F�j|� /�Se��/� /T/�x//�/�/=/ �/a/�/?�/,?�/P? �/�/�??�?9?�?�? o?O�?(O:O�?^O�? �O�O#O�OGO�OkO}O _�O6_�O/_l_�O�_ _�_�_U_�_y_o o �_Do�_ho�_	o�o-o �oQo�o�o�o�o@ R�ov��;� _���*��N�� G������7�̏ޏm� ���&�8�Ǐ\�돀� �!���E�ڟi�ӟ� ��4�ßX�j������ ��įS��w�������B�#��$FILE�_DGBCK 1�=��/���� ( ��)
SUMMAR�Y.DGL���M�D:�����D�iag Summ�ary��Ϊ
CONSLOG��������D�ӱConsole logE��ͫ��MEMCH�ECK:�!ϯ����X�Memory �Data��ѧ��{)��HADO�W�ϣϵ�J���S�hadow Ch�angesM�'�-���)	FTP�7Ϥ�3ߨ���Z�m�ment TBD���ѧ0=4)ETHERNET��������T�ӱEthernet \��figurati�onU�ؠ��DCSVRF�߽߫������%�� verify all���'�1PY���DI�FF�����[���{%��diff]������1R�9�K���� ���X��CHGD�������c��r����2pZAS� ��GD���k���z��FY3pbI[� �/"GD���s/�����/*&UP?DATES.� �/~��FRS:\�/��-ԱUpdates List�/���PSRBWLD'.CM(?���"<?��/Y�PS_ROBOWEL��̯�?�? ��?&�O-O�?QO�? uOOnO�O:O�O^O�O _�O)_�OM___�O�_ _�_�_H_�_l_o�_ �_7o�_[o�_lo�o o �oDo�o�ozo�o3 E�oi�o��� R�v���A�� e�w����*���я`� ��������O�ޏs� �����8�͟\��� ��'���K�]�쟁�� ��4���ۯj������ 5�įY��}������ B�׿�x�Ϝ�1��� *�g�����Ϝ���P� ��t�	�ߪ�?���c� u�ߙ�(߽�L߶��� ����(�M���q� � ���6���Z������ %���I���B������2�����h����$�FILE_� PR�� ��������MDONLY 1=.~�� 
 ��� q���������� ~%�I�m �2��h�� !/�./W/�{/
/�/ �/@/�/d/�/?�//? �/S?e?�/�??�?<? �?�?r?O�?+O=O�? aO�?�O�O&O�OJO�O �O�O_�O9_�OF_o_~
VISBCKL|6[*.VDv_|�_.PFR:\�_��^.PVisi�on VD file�_�O4oFo\_jo T_�oo�o�oSo�owo �oB�of�o �+������ �+�P��t������ 9�Ώ]�򏁏��(��� L�^�������5��� ܟk� ���$�6�şZ���~�����
MR_GRP 1>.�L��C4  ;B���	 W������*u����RHB ���2 ��� �?�� ���B��� ��Z�l���C���D������Ŀ��J�!�LL#��J���'F�5US���Qw^���ֿ� G�%�Fb���E��y.���9:�~�@]����A&�}A���-f�?�2�A��]r��E�?� F@ �������ھ��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<�,6\b��B��Y%���A��o=�@�eߋ�^�A��߲�v���r����� �
�C�.�@�y�d�� ��������������?�Z�lϖ�BH��� ��R�@(���E�������
0�P=?��P�V'��ܿ�� �B���/ ��@'�33:��.�g^&�@UUU�U���q	>u.�?!rX��	�-�=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!��7�:����D��@ D�� CYϥ��C������ ��0.��P/����/N� �/r��/���/�?? ;?&?_?J?\?�?�?�? �?�?�?O�?O7O"O [OFOOjO�O�O�O�O X�ߵ��O$_�OH_3_ l_W_�_{_�_�_�_�_ �_o�_2ooVohoSo �owo�o�i��o�o�o ��);�o_J� j������� %��5�[�F��j��� ��Ǐ���֏�!�� E�0�i�{�B/��f/�/ �/�/���/��/A�\� e�P���t�������� ί��+��O�:�s� ^�p�����Ϳ���ܿ � ��OH��o�
ϓ� ~ϷϢ���������� 5� �Y�D�}�hߍ߳� ���������o�1�C� U�y��߉����� ��������-��Q�<� u�`������������� ��;&_J\ ���������� ڟ�F�j4��� ������!// 1/W/B/{/f/�/�/�/ �/�/�/�/??A?,? e?,φ?P�q?�?�?�? �?O�?+OOOO:OLO �OpO�O�O�O�O�O�O _'__K_�o_�_�_ �_l��_0_�_�_�_#o 
oGo.okoVoho�o�o �o�o�o�o�oC .gR�v��� ��	���<�`� *<��`����� ޏ��)��M�8�q�\� ������˟���ڟ� ��7�"�[�F�X���|� ��|?֯�?�����3� �W�B�{�f�����ÿ ���������A�,� e�P�uϛ�b_������ �_��߀�=�(�a�s� Zߗ�~߻ߦ������� � �9�$�]�H��l� ������������#� �G�Y� �B������� z�������
ԏ:�C .gRd���� ��	�?*c N�r����� /̯&/�M/�q/\/ �/�/�/�/�/�/�/? �/7?"?4?m?X?�?|? �?�?�?�?��O!O3O ��WOiO�?�OxO�O�O �O�O�O_�O/__S_ >_P_�_t_�_�_�_�_ �_�_o+ooOo:oso ^o�o�op��o��  ��$��o�o� ~������� 5� �Y�D�}�h����� ��׏����
�C� .�/v�<���8����� �П����?�*�c� N���r��������̯ ��)��?9�_�q��� JO�����ݿȿ�� %�7��[�F��jϣ� ���ϲ�������!�� E�0�i�T�yߟߊ��� ���߮o�o��o>� t�>��b������ �����+��O�:�L� ��p������������� 'K6oZ� Z�|�~����� 5 YDi�z� �����/
// U/@/y/@��/�/�/�/ ���/^/???Q?8? u?\?�?�?�?�?�?�? �?OO;O&O8OqO\O �O�O�O�O�O�O�O_��O7_��$FNO ���VQ��
F�0fQ kP FLA�G8�(LRRM_�CHKTYP  �WP��^P��WP�{QOM�P_MsIN�P����P��  XNPSS�B_CFG ?�VU ���_���S ooIUT�P_DEF_OW�  ��R&hI�RCOM�P8o�$�GENOVRD_�DO�V�6�flT[HR�V d�edkdo_ENBWo k`�RAVC_GRP� 1@�WCa X "_�o_1U< y�r����� 	��-��=�c�J��� n��������ȏ�� ��;�"�_�F�X���ib�ROU�`FVX�P��&�<b&�8�?��埘��������  D�?�јs���@@g�B��7�p�)�ԙ���`S+MT�cG�mM����� �LQHOSTC��R1H���P�\�at�SM��f��\���	12�7.0��1��  e��ٿ����� ǿ@�R�d�vϙ�0�*��	anonymous����������֣([�� � � ����r����ߨߺ��� ��-���&�8�[�I� �π������ 1�C��W�y���`�r� �����ߺ������� %�c�u�J\n�� �������M�" 4FX��i��� ���7//0/B/ T/���m/��/ �/�/??,?�/P?b? t?�?�/�?��?�?�? OOe/w/�/�/�?�O �/�O�O�O�O�O=?_ $_6_H_kOY_�?�_�_ �_�_�_'O9OKO]O__ Do�Ohozo�o�o�o�O �o�o�o
?o}_R dv���_�_oo !�Uo*�<�N�`�r� �o������̏ޏ�?�Q&�8�J�\���>�E�NT 1I�� sP!􏪟  ����՟ğ������� A��M�(�v���^��� ��㯦��ʯ+�� � a�$���H���l�Ϳ�� ���ƿ'��K��o� 2�hϥϔ��ό��ϰ� ������F�k�.ߏ� R߳�v��ߚ��߾����1���U��y�<�QUICC0��b�t����1�����%����2&���u�!ROUTERv�R�d����!PCJOG�����!192�.168.0.1�0��w�NAME �!��!ROB�OTp�S_CF�G 1H�� ��Auto�-started^�tFTP�� ����� 2 D��hz���� U��
//./�v� ��/���/�/�/ �/�/�!?3?E?W?i? �/?�?�?�?�?�?�? ���AO�?eO�/�O �O�O�O�?�O�O__ +_NO�OJ_s_�_�_�_ �_
OO.OoB_'ovO Ko]ooo�oP_>o�o�o �o�oo�o5GY k}�_�_�_�� 8o��1�C�U�$y� �������ӏf���	� �-�?�����Ə ���ϟ����� ;�M�_�q���.�(��� ˯ݯ��P�b�t��� ��m���������ǿٿ �����!�3�E�h�� {ύϟϱ����$�6� H�J�/�~�S�e�w߉� ��jϿ��������*߀��=�O�a�s��YT_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��.FFF9E�3�?�FRS:DEFAULT�<�FANUC �Web Server�:
�����<�kO}O�O�O�O�O��W�R_CONFIGw O�� �?���IDL_CPU�_PC@�B���7P�BHUMI�N(\��<TGNR_�IO������PN�PT_SIM_D�OmVw[TPMO_DNTOLmV �]_PRTY�X7RTOLNK 1P����_o!o3oEoWo|io�RMASTElP���R�O_CFG��o�iUO��o�bC�YCLE�o�d@_?ASG 1Q����
 ko,>Pb t�������p��sk�bNUM�����K@�`IPCH��o��`RTRY_�CN@oR��bSC�RN����Q��� �b�`�bR���Տ���$J23_D_SP_EN	�����OBPROC��U�iJOGP1�SY@��8��?�!�T�!�?*�P�OSRE�zVKANJI_�`��o_��$ ��T�L�6͕����CL_LGP<�_����EYLOGGI�N�`��L�ANGUAGE YYF7RD w����LG��U�?⧕��x� �����Z=P��'0��$� NMC:\RSCH\00\���LN_DISP V��
���������OC�R.RDzVTA�{�OGBOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ��
�3�8��r��ۯ_MOx�_D�=R^��PL_NA_ME !6��p��!Defau�lt Perso�nality (�from FD)� �RR2eq 1�j)TUX)TX9��q��X dϏ8� J�\�n���������ȏ ڏ����"�4�F�X� j�|������2'�П �����*�<�N�`�r��<��������ү �����,�>�P�b�: �Rdr 1o�y �{\�, �3����� @D� M ��?�����?�<���A'�6�����;�	lʲ	 ��x�J����� �< �"��� �(pK���K ��K=*��J���J���JV���Z��ƌ��rτ́p@j��@T;f����f��ұ]�l��Ik��p������������b��3���o�  �
`�>�����bϸ�z��;꜐r�Jm��
� B�H�˱]Ӂt��q�	� p� W P�pQ�p��p|  Ъ�g����c�	'� � ���I� � � ����:����
�È=����"�s��	�ВI  �n @B� cΤ�\��ۤ��tq��y߁rN���  '������@2�@�����/��C��C�C�@ �C������
��A��  W @<�P�R�%
h�B�b�A��j������������Dz ۩��߹�����j���( �� -��C���'�7L�����q�Y������ �?�ff ���gy �����q+q��
�>+�  PƱj�( ����7	���^|�?����xZ��p<
6b<���;܍�<����<� <�&Jσ�AI�ɳ+�|���?fff?I��?&�k�@�.���J<?�` �q�.�˴fɺ�/ ��5/����j/U/�/ y/�/�/�/�/�/?�/0?q��F�?l? ?�?/�?+)�?�?ؿE�� E�I�G+� F��?)O �?9O_OJO�OnO�Of�BL޳B�?_h�.� �O�O��%_�OL_�?m_ �?�__�_�_�_�_�
��h�Îg>���_Co�_goRodo��o�GA�ds�q�C��o�o�o|���ؠ$]Hq���D���pC���pCHmZZ7t���6q�q���ܶN'�3A�A��AR1AO��^?�$�?��K�0±
=ç�>����3�W�
=�#�W��eۣצ�@�����{����<�����(�B�u���=B0������	L���H�F�G����G��H�U�`E���C�+����I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3�l� W���{��������՟ ���2��V�A�z��� w�����ԯ������ ��R�=�v�a����� �������߿��<� '�`�Kτ�oρϺϥ� �������&��J�\� G߀�kߤߏ��߳��� ����"��F�1�j�U� ��y���������� ��0��T�?�Q�����(�1��3/E�y����5����<��q3�8�����q4Mgs&�IB+2D�a���{�^^	�@�����uP2	P7Q4_A��M00bt��R��`����/   �/�b/P/�/t/�/  *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?��?�?O 2 F;�$�vGb�/�Aa��@�a�`�qC��C�@�o�O2���OF�� DzH@�� F�P D���O�O�ys<O!_3_E_�W_i_s?���@U@pZ.t22�!2~
  p_�_�_�_	oo-o?o Qocouo�o�o�o�o��Q ��+��1���$MSKCF�MAP  �5?� �6�Q��Q"~�cONREL7  
q3��bEXCFENB�?w
s1uXqFNC�_QtJOGOVLKIM?wdIpMrd�bWKEY?w�u�bWRUN�|�u�bSFSPDTY�xavJu3sSIGN?>QtT1MOT�Nq��b_CE_GRoP 1p�5s\r���j�����T�� ⏙������<��`� �U���M���̟��� ���&�ݟJ��C��� 7�������گ��������4�V�`TCOM_CFG 1q}��Vp�����
P�_/ARC_\r
jyUAP_CPL���ntNOCHECK� ?{  	r��1�C�U�g� yϋϝϯ����������	��({NO_WA�IT_L�	uM�NMTX�r{�[m�o_ERRY�2sy3� &��������r�c� ��T_�MO��t��, ��$�k�3�PAR�AM��u{���V[��!�u?�� =�9@345678901��&���E�W� 3�c�����{������� ����=��UM_RSPAC�E �Vv��$ODRDSP���jx�OFFSET_C�ARTܿ�DIS���PEN_FI�LE� �q��c֮�O�PTION_IO���PWORK kv_�ms � P(�R�Q
�j.j�	 ��Hj&6$�� RG_DSBL'  �5Js�\���RIENTTO>p9!C��PqfA�� UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	�lmb�`�x7J�`������a�< ���`� ��b, H(���H3k7HS�M5G�22G�?��Gp
��
��!��'|, CR�>�>q�GsuaT��3���  �4spBpyr  ]o��*SB_����=j]��t�q� ��rna �,��~�6  ��UPQ�|N��M�,k�!�	'�� � ��I�� �  ��%�=��ͭ����ba	���I  �n @��~����p����� �N	 W�  '!o�:q:�pC	 C�@@sBq��|��� m�
�T!�h@ߐ�n��$��Z�B	 �A����p� �-�qbz �P��t�_�������( �� -��恊�n�ڥD[A]Ѻ�b4�'!��~(p �?�ff� ��
����OZ�R���8��z���>΁  Pia��(�ವ@����ک�a�c�dF#?˙���x����<
�6b<߈;����<�ê<�? <�&�o&ς)�A�lcΐI�*�?offf?�?&c�ޒ�@�.uJ<?�`��Yђ ^�nd��]e��[g��G� �d<����1��U�@� y�dߝ߯ߚ����߼� 	���-������&��~"�E�� E��?G+� Fþ��� ��������&��J�(5��bB��AT�8� ђ��0�6���>���J� n�7��[m��0��h��1��>�M�I
�@��A�[���C-�)��?Ƀ��� /�Y���Jp��vav`CH�/������}!@�I�Y�'�3A��A�AR1A�O�^?�$�?�����±
=�ç>����3�W
=�#�����+e��ܒ������{����<���.(�B��u��=B0�������	��*H�F�G����G��H��U`E���C��+�-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�? O�?3OOWOBOTO�O xO�O�O�O�O�O�O_ /__S_>_w_b_�_�_ �_�_�_�_�_oo=o (oaoLo�o�o�o�o�o �o�o�o'$] H�l����� ��#��G�2�k�V� ��z���ŏ���ԏ� ��1��U�g�R���v� ����ӟ�������-�:�(���������a����xQ�c�,!3�8�}�<��,!4Mgs�����ɢIB+կ篴a?���{����A�/�e�S���w��P!�P�������7�`�ӯ�ϑ�R9��Kτ�oχϓϥ�  ���χ����)�� M����������{߉�����ߒߤ�������  )�G�q��_���2 wF�$�&Gb����n�[ZjM!C��s�@j/�A�S���F�� Dz���� F�P D��W����)������������x?��ͫ@@
9�E��E��E��
 v����� ��*<N`ܷ*P ���˨��1��$PARA�M_MENU ?�-�� � DEF�PULSEl	�WAITTMOU�T�RCV� �SHELL_�WRK.$CUR�_STYL��,OPT�/PT�B./("C�R_DECSN���,y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?��USE_PROG %�%�?�?�3CCR�����7�_HOST !F�!�44O�:T̰�?PCO)ARC�O�;_TIME�XB��  �GDEB�UGV@��3GINP_FLMSK�O��IT`��O�EPGA�P �L��#[CH��O�HTYPE����?�?�_�_�_�_ �_oo'o9obo]ooo �o�o�o�o�o�o�o�o :5GY�}� ���������1�Z��EWORD �?	7]	RS�`�	PNS��$��JOE!>�T�Es@WVTRACE�CTL 1x-��� ��3 ��Ӱ��Ɇ_DT Qy-��~�D � ��oӱ4� P :�L :�GP:�D :�T@ :�8�8�	8�U
8�8�8�8�E8�8�X@:�8�U8�8�8�8��:�8�8�x�:�A8�P�:�d :�8�A8���:�
�:�!8�E"8�#8���:�%8�U&8�'8�(8�)8�Q*8���:�,8�-8�U.8�/8�08�18� ,���ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�X�(�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_d��_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п�_� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$)��$PGTRACELEN  #!�  ���" �8&_UP �z���g!�o S!h 8!_C�FG {g%�Q#"!x!�$J �" �|"DEFSPD �|�,!!J ��8 IN TRL �}�-" 8�(I�PE_CONFI�� ~g%��g!�$�$�"8 LI�D�#�-74GR�P 1�7Q!��#!A ���&�ff"!A+33D��� D]� C�À A@+6�!��" d�$�9�9*1*0� 	 +9�-+6��? ´	C�?�;B @3AO�?OIO3OmO�"!>�T?�
�5�O�O�N�O =?��=#�
�O_ �O_J_5_n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_ Roxoco�o�o�o�o�o �o�o>)bM���;
V7.1�0beta1�$�  A�E>�rӻ�A " �p�?!G��q>�嚻r��0�q��޻qBQ��qA\��p�q�4�q�p�"�BȔ2�D�V�h�w�!�p�?�?)2{ȏ w�׏���4��1� j�U���y�����֟�� ����0��T�?�x� c�������ү����!o �,�ۯP�;�M���q� ����ο���ݿ�(π�L�7�p�+9��sF@ �ɣͷϥ�g% ������+�!6I�[� �������ߵߠ����� ����!��E�0�B�{� f����������� ��A�,�e�P���t� ����������� =(aL^��� ����'9$ ]�Ϛ��ϖ����� ��/<�5/`�r߄� �ߏ/>�/�/�/�/�/ ?�/1??U?@?R?�? v?�?�?�?�?�?�?O -OOQO<OuO`O�O�O �O�O���O_�O)__ M_8_q_\_n_�_�_�_ �_�_�_o�_7oIot ���o�o���o�o �o(/!L/^/p/�/{ *o������� ��A�,�e�P�b��� �������Ώ��+� =�(�a�L���p����� �Oߟ񟠟� �9�$� ]�H���l�~�����ۯ Ư���#�No`oro�o n��o�o�o�oԿ�� �8J\ng���� vϯϚ�������	��� -��Q�<�u�`�r߫� ���ߺ�������;� M�8�q�\�������� z������%��I�4� m�X���|��������� ��:�L�^���Z�� ���������$� 6�H�Swb� ������// =/(/a/L/�/p/�/�/ �/�/�/?�/'??K? ]?H?�?��?�?f?�? �?�?O�?5O OYODO }OhO�O�O�O�O�O�O &8J4_F_��� �_�_��_�_"4 -o�O*ocoNo�oro�o �o�o�o�o�o) M8q\���� �����7�"�[� m��?����R�Ǐ��� ֏�!��E�0�i�T� ��x��������_$_ V_ �2�l_~_�_������R�$PLID_�KNOW_M  ��T�|����SV ��U�͠�U ��
��.�ǟR�=�O������mӣM_GROP 1��!`0u���T@ٰo�ҵ�
���Pзj��` ���!�J�_�W�i�{� �ϟϱ����������V��MR�����T��s�w� s��ߠ޴� �߅��ߩ߻�����A� ��'������ ��������=��� #���������}�������S��ST��1 1Ն�U# ���0�_ A .��,> Pb������ ��3(iL^�p�����2r*���<-/�3/)/;/M/4 f/x/�/�/5�/�/�/�/6??(?:?�7S?e?w?�?8�?�?�?�?MAD  d#`�PARNUM  �w�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a��OT_CMP_0��B@�P@'˥T�ER_CHK'U���˪?R$_6[RS8l�¯��_MOA@�_�U_�_RE_RES_G ��>�o o8o+o\oOo�oso�o �o�o�o�o�o�o�W �\�_%�Ue B af�S� ����S 0����SR0�� #��S�0>�]�b��S�0�}������RV 1�x����rB@c]��}t�(@c\��}��D@c[�$����RTHR_IN�Rl�DA��˥d,�M�ASS9� ZM�M�N8�k�MON_QUEUE ���X˦��x� RDNP�UbQN{�P[��ENqD���_ڙEXE韌ڕ�@BE�ʟ��O�PTIOǗ�[��P�ROGRAM %��%��ۏ�O��?TASK_IAD0�OCFG ���xtO��ŠDATA��]�Ϋ@��27� >�P�b�t���,����� ɿۿ�����#�5�G�^��INFOUӌ�������ϭϿ����� ����+�=�O�a�s� �ߗߩ߻��������4^�jč� yġ~?PDIT �ί|c���WERFL
���
RGADJ ��n�A����?�����@���IORI�TY{�QV���MPGDSPH�����Uz�y���OTOEy��1�R� (!�AF4�E�P]����!tcph����!ud��!�icm��ݏ6�XYm_ȡ�R��ۡ)� *+/ ۠�W:F�j ������%@7[B�*��OPORT#�BC۠�����_CAR�TREP
�R� S�KSTAz��ZSS�AV���n�	2500H863��P�r�$!�R����q�n�}/�/�'^� URGE�B��6rYWF� DO{�r�UVWV��$�A�WR�UP_DELAY� �R��$R_HOTk��%O]?�$�R_NORMAL�k�L?�?p6SEMI�?�?�?3AQSKI�P!�n�l#x 	1/+O+ OROdO vO9Hn��O�G�O�O�O �O�O_�O_D_V_h_ ._�_z_�_�_�_�_�_ 
o�_.o@oRoovodo �o�o�o�o�o�o�o *<Lr`����n��$RCVT�M�����pDC�R!�LЈqC�q�C�2AC�ĳu?�A�>�R�<|�{4M��l�� ���´�ʿ�������[�|���4Oi��O <
6�b<߈;܍��>u.�?!<�&{�b�ˏ ݏ��8�����,�>� P�b�t���������Ο ���ݟ��:�%�7� p�S������ʯܯ�  ��$�6�H�Z�l�~� ������ƿ���տ� ��2�D�'�h�zϽ��� ����������
��.� @�R�d�Oψߚ߅߾� ����������<�N� ��r��������� ����&�8�#�\�G� ����}����������� S�4FXj|� �������� 0T?x�u� ���'//,/>/ P/b/t/�/�/�/�/�/ �/�?�/(??L?7? p?�?e?�?�?��?�?  OO$O6OHOZOlO~O �O�O�?�?�O�O�O�O  __D_V_9_z_�_�? �_�_�_�_�_
oo.o�@oRodovo�X�qGN_ATC 1��� AT&�FV0E0�k�ATDP/6/9�/2/9�hAT�A�n,AT�%G1%B960��i+++�o,��aH,�qIO_TYPE  �u��sn_�oREFP�OS1 1�P{O x�o�Xh_ �d_�����K� 6�o�
���.���R�����{{2 1�P{ ���؏V�ԏz����q3 1��$�6�p���ٟ���S4 1�����˟���n���>%�S5 1�<�N��`�����<���S6 1�ѯ���/������ѿO�S7 1� f�x���ĿB�-�f��S8 1������Y�������y�SMA�SK 1�P  q
9�G��XNOM����a~߈ӁqMO�TE  h�~t��_?CFG �������рrPL_RAN�G�ћQ��POWE/R ��e���SM_DRYPR/G %i�%��J���TART ��
�X�UME_PR�O'�9��~t_EX�EC_ENB  y�e��GSPD��p����c��TDB����RM��MT_�!�T���`OB�OT_NAME �i���iOB�_ORD_NUM� ?
�\q�H863  ��T��������bP�C_TIMEOU�T�� x�`S23�2��1��k L�TEACH ?PENDAN ��ƅ�}���`M�aintenance Cons�R�}�m
"{�dKC�L/Cg��Z ���n� No Use}�	��*�NPO��х����(CH_Lf�������	�~mMAVAIL���{��ՙ�SPA�CE1 2��| d��(>��&����p��M,8�?�ep/eT/�/ �/�/�/�W//,/>/ �/b/�/v?�?Z?�/�? �9�e�a�=??,?>? �?b?�?vO�OZO�?�OP�O�Os�2�/ O*O<O�O`O�O�_�_@u_�_�_�_�_[3_ #_5_G_Y_o}_�_�o��o�o�o�o[4 .o@oRodovo$�o�o ����"�	�7�[5K]o��A�� ��	�̏�?�&�T�[6h�z�������^� ԏ���&��;�\�C�q�[7��������͟ {���"�C��X�y�`���[8����Ưد ꯘ��0�?�`�#�u���}ϫ�[G �Ni� �ϋ
G� ����$�6�H� Z�l�~ߐ��8 ǳ�� ���߈��d(�� �M�_�q����� �������?���2�%� 7�e�w����������� ���������!�RE� W�����������?Q `�� @0��� �rz	�V_� ����
/L/^/|/ 2/d/�/�/�/�/�/�/ ?�/�/�/*?l?~?�? R?�?�?�?�?�?�?�?�2O�?
��O[_MODE  ��^�IS ���vO,*ϲ�O-_���	M_v_#dCWOR�K_AD�Ml[�P%aR  ���ϰ�P{_�P_INT�VAL�@����JR_OPTION�V� �EBpVAT_GRP 2���w�(y_Ho �e_vo�o�oYo �o�o�o�o�o*< �bOoNDpw�� ����	���?� Q�c�u�����/���Ϗ Ꮳ����)�;���_� q���������O�ɟ� ��՟7�I�[�m�/� ������ǯٯ믁�� !�3���C�i�{���O� ��ÿտ���ϡ�/� A�S�e�'ωϛϭ�o� ��������+�=��� a�s߅�Gߕ߻����� ����'�9�K�]��� �����y�����������5�G�Y��E�$�SCAN_TIM�AYuew�R ��(�#((�<}0.aaP%aP
Tq>��Q��o�����O+O2/��:	d/JaR��WY��^���^R^	�r  P��w� �  8�P��	�D�� GYk}���������Qp/@/R//)P�;�o\T��Qp�g-�t�_D�iKT��[  � lv%������/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OWW�#�O�O �O�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_olO~Od+ No`oro�o�o�o�o�o �o�o&8J\ n������u�  0�"0g�/�-� ?�Q�c�u��������� Ϗ����)�;�M� _�q�����$o��˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�����Do�� ������ҿ����� ,�>�P�b�tφϘϪπ����������w
�  58�J�\�n߀ߒ� �կ���������	�� -�?�Q�c�u������ ��-���� � �2�D�V�h�z�����������������;�& ��%�	123456{78�" 	��/� `r�������� (:L^p���� ���� //$/6/ H/Z/l/~/��/�/�/ �/�/�/? ?2?D?V? h?�/�?�?�?�?�?�? �?
OO.O@Oo?dOvO �O�O�O�O�O�O�O_ _*_YON_`_r_�_�_ �_�_�_�_�_ooC_ 8oJo\ono�o�o�o�o �o�o�oo"4F Xj|���������	��s3��E�W�{�Cz  �Bp��   ���2���z�$SC�R_GRP 1��(�U8(�\x�^ @�  �	!�	 ׃���"�$�  ��-��+��R�w�7���D~������#����O����M-10iA 8909905 Ŗ5 ?M61C >4���Jׁ
� � ��0�����#�1�	"�z�������¯Ҭ ���c� ��O�8�J�������!�����ֿ��B�y���������9A��$�  @��<�D �R�?��d���Hy��u�O���F@ F�`�§�ʿ�϶��� ����%��I�4�m��<�l߃ߕߧ߹�B���\����1��U� @�R��v������ �����;���*<�=�
F���?�d�<�>gm���@�:�n�� B���З�Й���EL_DE�FAULT  ~����B��MIPOWE?RFL  �$�1 WFDO� $��ERVENT 1������"�pL!DU�M_EIP��8���j!AF_IN�E �=�!FT$���!��4� ��[!RPC_MAIN\�>�J�nVIS�w=���!TMP�PU��	d��?/!
PMON_�PROXY@/�e ./�/"Y/�fz/�/�!RDM_SR�V�/�	g�/#?!�R C?�h?o?!%
pM�/�i^?�?�!RLSYNC̼?8�8�?O!gROS�.L�4�? SO"wO�#DOVO�O�O �O�O�O_�O1_�OU_ _._@_�_d_v_�_�_ �_�_o�_?oocoi�ICE_KL ?�%y (%S?VCPRG1ho8��e���o�m3�o�o�`4 �`5(-�`6PU�`7x}�`H���l9��{�d :?��a�o��a�oE� �a�om��a���aB ���aj叟a���a �5��a�]��a��� �a3����a[�՟�a�� ���a��%��aӏM��a ��u��a#����aK�ů �as���a��mob�` �o�`8�}�w������� ɿ���ؿ���5�G� 2�k�VϏ�zϳϞ��� �������1��U�@� y�dߝ߯ߚ��߾��� ����?�*�Q�u�`� ����������� �;�&�_�J���n������������sj_D�EV y	��MC:P�_]OUT"�,REC 1��Z� d   	 	�������
 ��PJ�%6 (�&�[w��,�*  VT - �- �A�- c|�P��� ��//B/0/f/x/ Z/�/�/�/�/�/�/�/ ?�/?P?>?t?b?�? �?�?�?�?�?�?OO OLO:OpO�OdO�O�O �O�O�O�O�O$__H_ 6_X_~_l_�_�_�_�_ �_�_�_ ooDo2oTo zo\o�o�o�o�o�o�o �o.R@vd ����},�� ��4�"�X�F�|��� p�����֏ď���� 0��@�f�T���x��� ��ҟ�Ɵ���,�� <�b�P���h�z����� �ί��(�:��^� L�n�p�������ܿ� п� �6�$�Z�H�j� ��rϴϢ�������� ��2�D�&�h�Vߌ�z� �ߞ�����������
�@�.�d�R��ZjV� 1�w P�m���	x  P� ���
TY�PEVFZN_�CFG ���d7�G�RP 1�A�c� ,B� A� D�;� B��� � B4RB{21HELL:�i�(
� X�|���%RSR�� ��E0iT�x ������/�Sew������%w������#�������2#�d�����HK 1��� �k/f/x/�/�/�/ �/�/�/�/??C?>?�P?b?�?�?�?�?��OMM ����?���FTOV_ENB� ���+�HOW_R�EG_UIO��I_MWAITB�.JKOUT;F��LIwTIM;E���O�VAL[OMC_UN�ITC�F+�MON�_ALIAS ?�e�9 ( he ��_&_8_J_\_��_ �_�_�_�_j_�_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]n��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� ���������ӟ~��� 	��-�?��c�u��� ����V�ϯ����� �;�M�_�q������ ��˿ݿ����%�7� I���m�ϑϣϵ�`� ������ߺ�3�E�W� i�{�&ߟ߱������� ����/�A�S���w� ����X������� ���=�O�a�s���0� ������������' 9K]���� b���#�G Yk}�:��� ���/1/C/U/ / f/�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_O
O�O�O�O �O�OvO�O__%_7_��C�$SMON_�DEFPRO ����`Q� *SY�STEM*  d�=OURECAL�L ?}`Y (� �}4xcop�y fr:\*.�* virt:\tmpback�Q�=>192.16�8.4�P46:6976 �R�_�_�_�K}5�Ua�_�_�V��_goyo�o}9�Ts�:orderfil.dat.l@oVo��o�o}0�Rmdb:+o�o�Q�obt �c�_2o?U�� 
�o��Sod�v�����
xyzrate 61 +�=�O�����������2848 ��ҏc�u� ���o�o56�ٟ��� "��5�џb�t���r�6����emp:�2392 W����:��.��*.d��Ư Яa�s����� +�=� O�����)�Ҳ�� ҿc�uχϚ���5�ͧ �������"���̨�� b�t߆ߙ����Q�U� ����
������T��� g�y��ϰ�9�T��� ��	�߷�@���c�u� ����-�?������� ����N�_q��� ��:L���&��p5372?��b t����4�5�� ��"��5�b/t/��/������p4016 W/�/�/�/��/ �)�/`?r?�?���;? M?�?�?O'�4�? �?cOuO�O��5/�' �O�O�O/"/�O�(�O b_t_�_����IDV_��_�_o�_�_6  �_goyo�o�O�O9_T_ �o�o	_�o@_�oc u��_-o?o�_�� �o��No_�q��� �o�o1�oݏ���&��J[�m������$SNPX_AS�G 1�������� P� 0 '%�R[1]@1.1,����?���%֟� �&�	��\�?�f��� u��������ϯ��"� �F�)�;�|�_����� ��ֿ��˿���B� %�f�I�[Ϝ�Ϧ��� ��������,��6�b� E߆�i�{߼ߟ����� ������L�/�V�� e���������� ��6��+�l�O�v��� ������������2 V9K�o�� �����&R 5vYk���� �/��<//F/r/ U/�/y/�/�/�/�/? �/&?	??\???f?�? u?�?�?�?�?�?�?"O OFO)O;O|O_O�O�O �O�O�O�O_�O_B_ %_f_I_[_�__�_�_ �_�_�_�_,oo6obo Eo�oio{o�o�o�o�o �o�oL/V� e������� �6��+�l�O�v��������PARAM ������ W�	��P�����OFT_KB_CFG  ������PIN_SI/M  ���C��U�g�����RVQS�TP_DSB,��򂣟����SR ��/�� & M�ULTIROBO�TTASK������TOP_ON_ERR  ����PTN �/�@�A�	�RING_PR�M� ��VDT_GRP 1�ˉ�  	������ ������Я����� *�Q�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߣߠ߲������� ����0�B�i�f�x� ������������� /�,�>�P�b�t����� ����������( :L^p���� ��� $6H Z�~����� ��/ /G/D/V/h/ z/�/�/�/�/�/�/? 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�__\_��VPRG_�COUNT��8@���RENBU��U�M�S��__UPD� 1�/�8  
s_�oo*oSoNo `oro�o�o�o�o�o�o �o+&8Jsn �������� �"�K�F�X�j����� ����ۏ֏���#�� 0�B�k�f�x������� ��ҟ������C�>� P�b���������ӯί������UYSDOEBUG�P�P�)��d�YH�SP_PA�SS�UB?Z�L�OG ��U��S)�#�0�  ���Q)�
MC:�\��6���_MPC ���U���Qñ8�� �Q�SAV ������ǲ&��ηSV;�TEM_TIME 1��[� (m�=&�:�:�}YT1SVGU�NS�P�U'�U����ASK_OPT�ION�P�U�Q�Q���BCCFG ��[u� n�A�a�`a�gZo��߃� ���߹�������:� %�^�p�[����� ���� �����6�!�Z� E�~�i���������&�������&8�� nY�}�?��� � ��(L: p^������ �/ /6/$/F/l/Z/ �/~/�/�/�/�/�/�/ �/2?8 F?X?v?�? �??�?�?�?�?�?O *O<O
O`ONO�OrO�O �O�O�O�O_�O&__ J_8_n_\_~_�_�_�_ �_�_�_o�_ o"o4o joXo�oD?�o�o�o�o �oxo.TBx ��j����� ���,�b�P���t� ����Ώ��ޏ��(� �L�:�p�^������� ʟ��o��6�H� Z�؟~�l�������د ���ʯ ��D�2�h� V�x�z���¿���Կ 
���.��>�d�Rψ� vϬϚ��Ͼ������� *��N��f�xߖߨ� ��8���������8� J�\�*��n����� ��������"��F�4� j�X���|��������� ����0@BT �x�d���� �>,Ntb� �����/�(/ /8/:/L/�/p/�/�/ �/�/�/�/�/$??H? 6?l?Z?�?~?�?�?�? �?�?O�&O8OVOhO zO�?�O�O�O�O�O�O 
__�O@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<o^o�oro�o �o�o�o�o�o  J8n$O���� �X���4�"�X��B�v��$TBCS�G_GRP 2��B�� � �v� 
 ?�  ������׏�� �����1��U�g�z����ƈ�d, ����?v�	 HC{��d�>����~e�CL  B����Пܘ������\)��Y  A��ܟ$�B�g�B�Bl��i�X�ɼ���X��  D	J���r������C����үܬ���D�@v�=�W�j�}� H�Z���ſ���������v�	V�3.00��	mw61c�	*X�0P�u�g�p�>���v�(:�� ��p͟�w  O����p������z�JCFG [�B��� ��V��������=��=�c�q�K� qߗ߂߻ߦ������ ��'��$�]�H��l� ������������#� �G�2�k�V���z��� �����������p *<N���l�� �����#5G Y}h���� v�b��>�// /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?d?R? t?v?�?�?�?�?�?O �?*OO:O`ONO�OrO �O�O��O�O�O_&_ _J_8_n_\_�_�_�_ �_�_�_�_�_�_oFo 4ojo|o�o�oZo�o�o �o�o�o�oB0f T�x����� ��,��P�>�`�b� t�����Ώ������ �&�L��Od�v���2� ����ȟʟܟ� �6� $�Z�l�~���N����� دƯ�� �2��B� h�V���z�����Կ¿ ����.��R�@�v� dϚψϪ��Ͼ����� ��<�*�L�N�`ߖ� �ߺߨ����ߚ��� ����\�J��n��� ��������"���2� X�F�|�j��������� ������.TB xf������ �>,bP� t�����/� (//8/:/L/�/�ߚ/ �/�/h/�/�/�/$?? H?6?l?Z?�?�?�?�? �?�?�?O�?ODOVO hO"O4O�O�O�O�O�O �O
_�O_@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<oro`o�o �o�o�o�o�o�o& �/>P�/��� ������4�F� X��(���|�����֏ ����Ə0��@�B� T���x�����ҟ���� ��,��P�>�t�b� ������������� �:�(�^�L�n����� ��2d�����̿� $�Z�H�~�lϢϐ��� �����Ϻ� ��0�2� D�zߌߞ߰�j����� �����
�,�.�@�v� d����������� ��<�*�`�N���r� ������������& J\�t��B ������F 4j|��^��p��/�  2 �6# 6&J/6"��$TBJOP_G�RP 2����  ?i�X,i#�p,� ��x�J� �6$�  �_< �� �6$� @2 �"	 ߐC�� �&b � Cق'�!�!>�c��
559>�0�+1�33=�{CL� fff?+0?�ffB� J1�%�Y?d7�.��/>��2\)?0�5����;��hC=Y� �  @� �!?B�  A�P?�?��3EC�  Dp�!�,�0*BOߦ?��3JB��
:���Bl�0��0�$�1��?O6!Aə�A�ДC�1D�G6��=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH��1ts�A@333@?1� C�� �@�_�_&_8_>��D��UV_0�LP�Q30<'{�zR� @�0�V �P!o3o�_<oRifoPo ^o�o�o�oRo�o�o�o �oM(�ol�pP~��p4�6&�q�5	V3.00��#m61c�$�*(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�N�aF���F�^�lF���F�:�
F�)F���3G�G���G��G,I�R�CH`�C��dTDU�?D���D��DE(�!/E\�E���E�h�E��ME��sF�`F+'\FD���F`=F}�'�F��F��[
F���F���M;S@;Q�*�|8�`rz@/&�
8�6&<��1�w��^$ESTPARS�  *({ _#HR���ABLE 1̒p+Z�6#|�Q� (� 1�|�|�|�5'T=!|�	|�
|�|�T˕6!|�|�|����RDI��z!�ʟܟ� ��$���O ������¯ԯ�����	S��x# V���˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �U-����ĜP�9�K� ]�o��-�?�Q�c�u����6�NUM  V�z!� > � Ȑ����_CFGG �����!@b �IMEBF_TT�����x#��a�VER腣b�w�a�R 1=�p+
 (3�6"	1 ��  6!���� ������ �9�$�:�H� Z�l�~����������� ����^$��_���@x�
b MI_CWHANm� x� k�DBGLV;0o��x�a!n ETHER_AD ?�� �y�$"�\&n oROUT��!p*�!*�SNM�ASK�x#�255.h�fx^$�OOLOFS_D�I��[ՠ	ORQCTRL �p+ ;/���/+/=/O/ a/s/�/�/�/�/�/���/�/�/!?��PE_�DETAI��P�ON_SVOFF��33P_MON ��H�v�2-9ST�RTCHK ����42VTCOMPATa8�24:0�FPROG %��%MULTI?ROBOTTO!O<06�PLAY��L:_INST_MPe GL7YDUS���?�2LCK�LPKQ?UICKMEt �O��2SCRE�@>�
tps��2 �A�@�I��@_Y����9�	SR_GRP� 1�� ���\�l_zZg_�_ �_�_�_�_�^�^�o j�Q'ODo/ohoSe� �oo�o�o�o�o�o�o !WE{i�������	1?234567���!���X�E1�V[
� �}ipnl�/a�gen.htmno��������ȏ~��Panel _setup̌}�?���0�B�T�f�  ��񏞟��ԟ��� o����@�R�d�v��� ���#�Я����� *���ϯůr������� ��̿C��g��&�8� J�\�n�����϶��� ������uϣϙ�F�X� j�|ߎߠ����;��߀����0�B��*NU�ALRMb@G ?�� [���� �������� ��%�C��I�z�m�������v�S�EV  �����t�ECFG �Ձ=]/BaA$ �  B�/D
  ��/C�Wi{�� ����� PRց; �To\�o�I�6?K0(% ����0����� //;/&/L/q/\/�/0�/�/l�D �Q��/I_�@HIST� 1ׁ9  �(  ��(/�SOFTPART�/GENLINK�?current�=menupag�e,153,1 �Ec0p?�?�?�?/C�s� >?P=962n?��?
OO.O�?�?�136c?|O�O�O�OAOSO �?�O__0_�O�O_L u_�_�_�_:_�/�_�_ oo)o;o�__oqo�o �o�o�oHo�o�o%7I~��a81�ou ������o�� �)�;�M��q����� ����ˏZ�l���%� 7�I�[��������� ǟٟh����!�3�E� W����������ïկ �v���/�A�S�e� Pb������ѿ��� ���+�=�O�a�s�� �ϩϻ�������ߒ� '�9�K�]�o߁�ߥ� ���������ߎ�#�5� G�Y�k�}������ ���������1�C�U� g�y���v��������� ��	�?Qcu ��(���� )�M_q�� �6���//%/ �I/[/m//�/�/�/ D/�/�/�/?!?3?�/ W?i?{?�?�?�?���� �?�?OO/OAOD?eO wO�O�O�O�ONO`O�O __+_=_O_�Os_�_ �_�_�_�_\_�_oo 'o9oKo�_�_�o�o�o �o�o�ojo�o#5 GY�o}�������?��$UI_�PANEDATA 1������  	�}�0�B�T�f�x��� )����mt�ۏ ����#�5���Y�@� }���v�����ן���� ���1��U�g�N���.��� �1��Ï ȯگ����"�u�F� ��X�|�������Ŀֿ =������0�T�;� x�_ϜϮϕ��Ϲ������,ߟ�M��j� o߁ߓߥ߷������ `��#�5�G�Y�k��� ������������� ��C�*�g�y�`��� ������F�X�	- ?Qc����߫� ���~;" _F��|��� ��/�7/I/0/m/ �����/�/�/�/�/�/ P/!?3?�W?i?{?�? �?�??�?�?�?O�? /OOSOeOLO�OpO�O �O�O�O�O_z/�/J? O_a_s_�_�_�_�O�_ @?�_oo'o9oKo�_ oo�oho�o�o�o�o�o �o�o#
GY@} d��&_8_��� �1�C��g��_���� ����ӏ���^��� ?�&�c�u�\������� ϟ���ڟ�)��M� ����������˯ݯ 0�����7�I�[�m� ���������ٿ�ҿ ���3�E�,�i�Pύπ�φ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#������� � �$�6��Z�A�~�e� w����������� 2��V�h�O�����v��p��$UI_PA�NELINK 1��v�  ��  ���}1234567890����	- ?G ���o��� ��a��#5�G�	����p&���  R���� �Z��$/6/H/Z/ l/~//�/�/�/�/�/ �/�/
?2?D?V?h?z? ?$?�?�?�?�?�?
O �?.O@OROdOvO�O O �O�O�O�O�O_�O�O�<_N_`_r_�_�_�0,���_�X�_�_�_ o 2ooVohoKo�ooo�o �o�o�o�o�o�� ,>r}������ ������/�A� S�e�w��������я ���tv�z���� =�O�a�s�������0S ��ӟ���	��-��� Q�c�u�������:�ϯ ����)���M�_� q���������H�ݿ� ��%�7�ƿ[�m�� �ϣϵ�D�������� !�3�Eߴ_i�{�
�� �����߸������/� �S�e�H���~�� R~'�'�a��:�L� ^�p������������� �� ��6HZl ~���#�5���  2D��hz� ����c�
// ./@/R/�v/�/�/�/ �/�/_/�/??*?<? N?`?�/�?�?�?�?�? �?m?OO&O8OJO\O �?�O�O�O�O�O�O�O [�_��4_F_)_j_|_ __�_�_�_�_�_�_o �_0ooTofo��o�� �o��o�o�o, >1bt���� K����(�:�� ��{O������ʏ܏ �uO�$�6�H�Z�l� ��������Ɵ؟��� �� �2�D�V�h�z�	� ����¯ԯ������ .�@�R�d�v������ ��п���ϕ�*�<� N�`�rτ��O�Ϻ�Io ���������8�J�-� n߀�cߤ߇����߽� ���o1�oX��o|� ������������ �0�B�T�f������ ��������S�e�w�, >Pbt��'� ����:L ^p��#��� � //$/�H/Z/l/ ~/�/�/1/�/�/�/�/ ? ?�/D?V?h?z?�? �?�???�?�?�?
OO .O��ROdO�߈OkO�O �O�O�O�O�O_�O<_ N_1_r_�_g_�_7O�M�m�$UI_�QUICKMEN�  ���_AobREST�ORE 1��  �A|��Rto�o�im�o �o�o�o�o:L ^p�%���� ��o����Z�l� ~�����E�Ə؏��� � �ÏD�V�h�z��� 7�������/���
�� .�@��d�v������� O�Я�����ßͯ 7�I���m�������̿ ޿����&�8�J�� nπϒϤ϶�a����� ��Y�"�4�F�X�j�� �ߠ߲������ߋ����0�B�T�gSCR�E`?#m�u1sco`u2���3��4��5��6ʏ�7��8��bUS#ERq�v��Tp���Sks����4��5��6��7��8��`N�DO_CFG m�#k  n` `PDATE ����None�bSEUFRAM/E  �TA�n��RTOL_ABRqTy�l��ENB��~��GRP 1�ci�/aCz  A� ����Q�� $6BHRd��`U������MSK  h�����Nv�%�U��%���bVIS�CAND_MAXλI��FA?IL_IMG� �P�ݗP#��IMR_EGNUM�
,�[SIZ�n`��A�,VONTM�OU��@����2��a��a�����FR�:\ � �MC:\�\L�OG�B@F� �!�'/!+/O/�Uz MCV��8#UD1r&EX�{+�S�PPO6�4_��0'fnm6PO��LIb��*�#V���,fy@�'�/� =	�(wSZV�.����'�WAI�/STAOT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_J�MPERR 1��#k
  �2345678901dF �ψO{O�O�O�O�O�O _�O*__N_A_S_�_<
� MLOWc>
 ��_TI�=�'�MPHASE'  ��F��P�SHIFT�1 9�]@<�\�Do �U#oIo�oYoko�o�o �o�o�o�o�o6 lCU�y��� �� ��	�V�-�e�2����	VSF�T1�2	VMN�� �5�1G� ����%A�  B8*̀̀�@ pكӁb˂�у��z�ME@Ľ?�{��!c>&%��aM1��k�0��{ �$`0TDINGEND��\�O� �z����S��w��P���ϜREL�E�Q��Y���\�_ACTIV��:�R�A ��e����e�:�RD� ���Y?BOX �9�دV�6��02����190.0.��83��2�54��QF�	 ��X�j��1�?robot���   p��<���5pc��̿ �����7�����-�f�ZABC�����, ]@U��2ʿ�eϢω� �ϭϿ����� ��߀V�=�z�a�s߰�E�Z��1�Ѧ