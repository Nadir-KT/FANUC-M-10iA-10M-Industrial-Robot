��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1�~FPCUREQ1� � $SO{FT; T_ID��TOTAL_EQf� $� � NO��PS_SPI_I�NDE��$�X��SCREEN_�NAME ^�SIGN���� PK_FIL~	$THKYM�PANE�  	$DUMMY )� u3|4|G�RG_STR1� � $TIT�P$I��1��{�����5��6�7�8�9�0��z���T��1�1�1 '�1
'2"GSBN�_CFG1  �8 $CNV_�JNT_* |$�DATA_CMN�T�!$FLAG�S�*CHECK��!�AT_CEL�LSETUP � P $HO_ME_IO,G�}%�#MACRO�"�REPR�(-DR�UN� D|3S�M5H UTOBA�CKU0 � ?$ENAB��!oEVIC�TI� � D� DX�!2ST� ?0B�#$�INTERVAL�!2DISP_UNsIT!20_DOn6�ERR�9FR_F�!2IN,GRE5S�!0Q_;3!4C_WA�471�8G�W+0�$Y $D�B� 6COMW�!2MO� H.	� \rVE�1$qF�RA{$O��UDcB]CTMP1_5FtE2}G1_�3�B~�2���AX�D�#
 d �$CARD_EX�IST4$FS?SB_TYP!A?HKBD_SNB�1�AGN Gn �$SLOT_NUyM�APREV4DEBU� g1G ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP��U0LETE_OK��BUS�P_CR��A$;4AV� 0LACIw1�R�@�k �1$@MEN�@$D�V�Q`PvVAh{QL� OU&R ,A�0�!� =B� LM_O�
e=R�"CAM_;1� xr$A�TTR4�@� AN�NN@5IMG_H�EIGH�AXcWI7DTH4VT� �U�U0F_ASPE�C�A$M�0EX�P�.@AX�f�C�F�D X $�GR� � S�!.@B�PNFLI�`�d� �UIRE 3T!GI�TCH+C�`N� S&�d_LZ`AC�"�`SEDp�dL� J�4S�0� <za�!p;�G0 � 
$WARNM�0f�!p�@� -s�pNST� �CORN�"a1FL{TR{uTRAT� �T}p  $ACCa1�p��|{�r�ORI�P�C�kRTf0_S~B\qHG,]I1 [ T�`4�"3I�pTYD�@*2 3`#@� �!,�B*HDDcJ* C�d�2_�3_�4_�5�_�6_�7_�8_�9~4DB:�CO�$ <� �o�o�hK3� 1#`O_Mc@AC/ t � E#63NGPvABA� �c�1�Q8��`,��@nr1�� d�P�0e�]p,� cvnpUP&P�b26���p�"J�p_)R�rPBC��J�rĘߜJV�@U� B��s}��g1�"YtP_*0O�FS&R @� RcO_K8T��aIT�3�T�NOM_�0�1�p�34 >��D Ԑ� Ќ@��hPV��mE!X�p� �0g0ۤ�p��r
$TF�2C$7MD3i�TO�3�0yU� F� ��)Hw2tC1(�Ez�g0#E{"F�"F�40�CP@�a2 �@�$�PPU�3Nc)ύRևAX�!�DU��AI�3B�UF�F=�@1 �|pp���pPITV� PP�M�M��y��F�SIMQ�SI�"ܢVAڤT��=�w T�`(zM��P�B�qFACTb�@EW�P1��BTv?�MC�5 �$*1JB`p脎*1DEC��F����=�� �H0CHNS_EMP1�G$G��8��@_4��3�p|@P��3�TC c�(r/�0-sx��ܐ�� MBi��!����JR|� i�SEGFR���Iv �aR�TpN�C��PVF4>�bx &��f{u Jc!�Ja��� !28�ץ8�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb��Ӏq�۽�н����Lp�3�B���CRC�e�3CCp����c� �mcҞb�1J�cѿ�.�T���D$ICb�Cq��5r�ե��@v�'���E�V���zF��_��FR,pN��ܫ�?�84�0A�! �r�� �h�Ϩ��p�2�͕a��� �د�R�Dx Ϗ��o"2�7�!ARV�O`C�$LG�pV�B�1�P��@�t�aA�0'�|�+01Ro�� MEp`"1� CRA 3 A�ZV�g6p�O �FCCb�`�`F�`K������ADI��a� A�bA'�.p��p�`��c�`S4PƑ�a�AMIP��-`Y�3P�M��]pUR��QUA1  ]$@TITO1/S�@S�!����"0�DBOPXWO��B0!5�O$SK���2@�DBq�!"�"�PR�� 
� =���΁!# S q1$�2�$z���L�)$��/���� %�/�$Cr�!&?�$ENE�q�.'*?�Ú RE|�p2(H ���O�0#$L|3$�$�#�B[�;���FO�_D��ROS�r�#������3RIoGGER�6PApS|����ETURN�2n�cMR_8�TUw���0EWM���M�GN�P���BLA�H�<E���P��&$P� �'P@�Q3�CkD{��DQ���4��11��FGO_AWAY�BMO�ѱQ#!�DCS_�o)  �PIS�  I gb {s�C��A��[ �B$�S��AbP�@�EW-�TNTVճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_S}V�bEXCLU�:�nONL2��S1Y�*a&�OT�a'�HI_V�4��B���_ *P0� 9�9_z��p ���A;SG�� +nrr� @6Acc*b��G�#@E��V.iHb?fANNU�N$0.$fdID�U�2�SC@�`�i�a���j�fp�z��@I$2,�O�$FibW$}�O�T9@�1 $DUMMYT��da��d�n�� � �E- ` ͑HE4(sg��*b�SAB��SUFFmIW��@CA=��c5�g6�a�DwMSW�E. 8Q��KEYI5���TM`�10s�qA�vIN��p�ї!��/ D��oHOST_P!�r T��ta��tn��tsp�p�EMӰV��� SB�Lc ULI�0 � 8	=ȳ�r�D�Tk0�!1 � �$S��ESAMPL���j�۰f璱f���I��0��[ $SUB �k�#0�C��T�r#a�SAVʅ��c����C��P�fP$n0E��w YN_B#2� 0Q�DI{dlpO�(��9#$�R_�I�� �ENC�2_S� 3  5�C߰�f�- �SpU����!4�"g�޲r�1T���5X� j`ȷg��0�0K�4�<AaŔAVER�qĕ�9g�DSP�v��PC��r"��(���ƓoVALUߗHE��ԕM+�IPճ��OkPP ��TH���֤��P�S� �۰F��df�J� ��p��C1+6 H�bLL_DUs�~a3@{�0�3:���OTX"����s�r�0NOAUkTO�!7�p$)�H$�*��c4�(�Cy�%8�C, �"�&��L�� 8H *8�LH <6����c "�`, `Ĭ�kª�q���q��sq��~q��7*��8��9��0����U1��1̺1ٺ1�U1�1 �1�1ʥ2(�2����2̺2�ٺ2�2�2 �2��2�3(�3��3T��̺3ٺ3�3�U3 �3�3�4(�(���?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?g �@P?9��5�9�E�@A��a��A� ;p$T�P�$VARI�:�Z���UP2�P< ���TDe����K`Q���a��BAC�"= T�p��e$�)_,�bn�kp+ IF�IG�kp�H  ��P���@`�!>�t ;E��sC�ST�D� D���c�<� 	C��{� �_���l���R  �����FORCEUP�?b��FLUS�`H��N>�F ���RD_CM�@E������ p��@vMP��REMr F�Q��1k@���7�Q
K4	NJ�5EF1Fۓ:�@IN2Q��sOVO�OVA�	�TROV���DT<Հ�DTMX�  ��@�
ے_PH",p��CL��_TpEȓ@�pK	_(�Y_T���v(��@A;QD� ������!0tLܑ0RQ���_�ad����M�7�CL�d�ρRIV'�{��E�ARۑIOHPCȸ@����B�B��CM�9@���R �GC3LF�e!DYk(Ml�ap#5TuDG���� �%��FSSD �s? P�a�!�1����P_�!�(�!1R��E�3�!3�+5�&O�GRA��7�@��i;�PW��ONn��EBUG_SD2H��P{�_E A�`ꁣ��TER�M`5Bi5P��ORI#e0C�9S�M_�P��e0D�9T�A�9E�9UP\�F�� -�A{�A�dPw3S@B$SEG��:� EL{UUSE.�@NFIJ�B$��;1젎4�4C$UFlP=�$,�|QR@"��_G90Tk�D��~SNST�PATx����APTHJ��E�p%B`�'EC���AR$P�I�aSHFTy�A�A�H_SHORР꣦6% �0$�7PE��E�GOVR=��aPI�@��U�b �QAYLOW���IE"�r�A8��?���ERV��XQ �Y��mG>@�BN��U\��R2!P.uA�SYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC����EP;�uP;�6WOR�>@M`�!�GRSM5T6�G3�GR��13�aPAL@���`�q�u_H � ���'TOCA�`P	P�`$OP����pѡ�`0O��R%E�`R4C�AO�p��Be�`R�Eu�h|�A��e$PWR�3IMu�RR_�cN�\�q=B I&2H���p_ADDR��H_LENG�B�q�qT�q$�R��S�JڢSS��SKN��u\�0�u̳�uٳSE�A��jrS��MN�!K������b����O�LX��p����`ACRO3pJ�@��X��+��Q��6�OUP3�b_�IX��a�a1��}򚃳���(�� H��D��ٰ��氋�VIO2S�D������	�7�L $xd��`Y!_OFFr^�PRM_��"�_HTTP_+�H:�wM (|pOBJ]"l�p��$��LE~C�d���N � \��֑AB_�Tq�b��S�`H�LVh��KR"uHITC�OU��BG�LO�q���h�����`���`SS� ���HQW�#A:�Oڠ<`�INCPU2VISIOW�͑��n��t�o��to�ٲ �IO�LN��P 8��R���p$SLob� PUT_n�$�p��P& ¢��Y F�_AS�"Q��$AL������Q  U�0�	P4A��^���ZPH�Y��-��u���U9OI �#R `�K�����$�u�"pP pk���$��������UJ5�S-���NE�6WJOGKG̲DI�S���Kp���#T� (�uAVF�+`�C�TR�C
�FLAG�2�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w�  m�_�{0a�^��cg��� 4�����Ǝ���{0��� SCH_���a7��N�d�VW���E �"����4��UM�A�r�`LJ�@�DAUfՃEAU�p��d|�r�GqH�b����BOO��WL ?�6 I�T��y0�REC���SCR ܓ�Dx
�\���MARGm� !��զ ��d%�����	S����W���U� ��JGM[�MNCH|J���FNKEY\��K��PRG��UF���7P��FWD��H]L��STP��V��=@��А�RS��HO`����C9T��b ��7�[�UL���6�(R�D� ����Gt��@P�O��������MD�F�OCU��RGEX.��TUI��I��4�@�L�����P����`��P��NE��CANA��Bj�oVAILI�CL !~�UDCS_HII4���s�O�(!�S���S��a���BUFF�!X�?PTH$m���vP`�ěԃ�AtrY��?P��j�3��`OSU1Z2Z3Z�|�� Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�C���K�&&8���![ LQ��+00� 	P���`#qdt
�U�dw�<���_ \ �?�4Г�\��Ѩ#��MC4�] ��C�LDPL��UTRQ�LI��dڰ�)�$F�LG&�� 1�#�D���'B�LD�%�$�%ORGڰ5�2�PV� �VY8�s�T�r �#}d^ ���$6��$�%�S�`T� �B0�4>�6RCLMC�4]?0o?�9세�MI�p}dg_ d=њRQ�=�DSTB�p�c ;F�HHAX�R� JHdLEXCE�Sra�BM!p�a`���/B�T�F��`a�p=F_A7Ji��K�bOtH�0K�db \�Q���v$MBC�L�I|�)SREQUI�R�R�a.\o�AXDESBUZ�ALt M���c�b�{P����2FANDRѧ`�`d;Ҙ2�ȺSDC��N�I�Nl�K�x`��X� N�&��aZ���UPS�T� ezrLO�C�RIrp�EX�<fA�p�9AX�0OwDAQ��f XY�3OND�rMF,� �f�s"��}%�e/� �� �FX3@IGG>�� g ��t"���ܓs#N�s$R�a%��iL��hL�v�@��DATA#?pE��%�tR��Y�Nh t $MD`qI}�)nv� ytq�yt�HP`�Pxu��(�zsANSW)�yt@��yu�D+�)Yr���0o�i[ �@CUw�V�p� 09AARR2��j� Du�{Q��7Bd$OCALIA@��G�:�2��RIN��"�=<��INTE��C�k�r^�آ�]���_N�qlk���9�D����Bm��DIVFD�H�@���qnI$�V,��S�$���$Z�X�o�*�����oH �$�BELT�u!ACCEL�.�~�=��IRC�� ���D�T<�8�$PS�@�"L���r��#^�S�xEы T�PATH3����I���3x�p�A_@W��ڐ���2nC���4�_MG�$D�D��T���$FW��Rp9��I�4��D}E7�PPABN��ROTSPEE�[g�� J��[�C@�4���$USE_d+�VPi��SYY����1 �aYN!@A��ǦOFF�qǡM�OU��NG���O9L����INC�tMa�6��HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]�ౌB��VE��#�y�2�3_UP񕋳LOWL���p� B���Du�9B#P`�x ����BCv�r�MOSI���BMOU��@�7P�ERCH  ȳOV��â
ǝ���� D�ScF�@MP����B� Vݡ�@y�j�LU0k��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A���x�����N`�F�RT1I�A$��MOUІЀHB�BS0�p7D5����ë�Z�DUM2�ԓS_BCKLSH_Cx�k���� ϣ���=���ޡ �	ACLAL"q��1М�@��CHK� �S�RTY��^�%�E1Qq_�޴_UM��@�C#��SCL�0�r�LMT_J1_L��9@H�qU�EO�p�b�_�e�k�e�SPC��u���N�PC�N�Hz \P�2�C�0~"XT��CN_:�N9��I�SF!�?�V���U� /���x�T���CB!�SH�:��E�E1TрT����y���T��P�A ��_P��_ � =������!�����J6 L�@��OG|�G�TORQU��ONֹ��E�R��H�LE�g_W2���_郠����I�IJ�I��Ff`xJ�1X�~1�VC3�0BD:B�1�@SB�JRKF9�0D�BL_SM��2M��P_DL2GR�V����fH�_��d���COS���LNH� �������!*,��aZ���fMY��_(�TH��)T�HET0��NK2a3���"��CB�&CB�CAA�B�"�0�!��!�&SB� 2N�%GTS�Ar�CI Ma�����,4#97#$DU���H\1�  �:Bk62�:AQ(rSf'$NE�D�`I��HB+5��$̀�!A�%��5�7���LPH�E�2���2SC% C%�2-&FC0JM&̀EV�8V�8߀LVJUV!KV/KV=KVKKVYKVgIH�8FRPM��#X!KH/KH=KUHKKHYKHgIO�<�O�8O�YNOJO�!KO/KO=KOKKO
YKOM&F�2�!+i%�0d�7SPBALA�NCE_o![cLE60H_�%SPc� &��b&�b&PFUL�C�h�b�g�b%p�1=k%�UTO_���T1T2�i/�2N ��"�{�t#�Ѱ`�0(�*�.�T��OÀ<�>v INSEG"�ͱ�REV4vͰl�DI�F�ŕ�1lzw��1m��OBpq�я?��MI{���nLCHgWARY�_�AB��~!�$MECH�!�o ��q�AX��P�����7Ђ�`n 
p�d(�U�ROB���CRr�H���k(��MSK_f`�p� P �`_��R /�k�z�����1S�~��|�z�{���z��qIN�Uq�MTCOM�_C� �q  ����pO�$NO�REn����pЂ7r 8p GRe�u�SD�0AB�$?XYZ_DA�1a���DEBUUq�������s z`$��COD�� L���p��$BUFIwNDX|�  <��MORm�t $فUA��֐����y��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p} =�C�}pt�@b�D��FRIrӚ�T��RO@ \�Ex}'���OPWOY�q�v0Y�SYS�BU/@v�$SOP�ġd���ϪUΫ}pPgRUN����PA���D���rɡL�_OUbo顢q�$)�/IMAG��w��0�P_qIM��L�IN�v�K�RGOVR!Dt��X�(�P*�J�|��0L_�`]��0�RB1�0��ML��ED}��p ��%N�PMֲ��Uc�w��SL�`q�w x �$OVSL4vS;DI��DEX�� ��#���-�V} *�N4�\#�B�2�G�B�2_�M�x� �q�>E� x Hw��p^��ATUSW����C�0o�s���BTMT�ǌ�I�k�4��x�԰q�y Dw�E&���@E�r��7�8�жЗ�EXE�����������f q�z �@w���UP'��$�pQ�XN�����x����� �PG΅�{ h $SUB����0_���!�_MPWAIv�P7�&��LOR�٠F\p˕�$RCVFAI�L_C��٠BWD�΁�v�DEFSP>!p | Lw����Я�\���UNI+�����H�R�+�}�_L\pP����P��p�}H�> �*�j��(�s`~�N�`KET�B�%�J�PE Ѓ~z��J0SIZE�����X�'���S�OR~��FORMAT�``��c ��WrEM�t��%�UX��G���PLI��p� � $ˀP_SWqI�pq�J_PL��?AL_ ����ХA��B��� C��Dn�$E��.��C_�U�� �� � ���*�J�3K0����TIA4��5��6��MOM���������ˀB��AD����������PU� NR�������G��m��� A$PI�6q��	 �����K4�)6��U��w`��SPEEDgPG������ ��Ի�4T�� �p @��SAMr`���\�]��MOV _�_$�npt5��5���1���2���������'�S�Hp�IN�'�@�+�����4($4+T+GAM�MWf�1'�$GE�T`�p���Da���
�
pLIBR>�II.2�$HI=�_g�t�$�2�&E;��(A�.� �&LW�-6<�)56��&]��v�p��V��$PDCK��D�q��_?����� q�&���7��4���9�+� �$IM_SR�pD�s�rF�L�r�rLE���Om0H]��0�	-�pq���PJqUR_S�CRN�FA���S_?SAVE_D��dE@�NOa�CAA�b� d@�$q�Z�Iǡs	�I � �J�K� ����H� L��>�"hq��� ���ɢ�� bW^U�S�A�S��M4� ��a��)q`��3�WW� I@v�_�q�.MUAo��� � $PY�+�$W�P�vNG�{��P:��RA��RH��RO�PL�����qP� ��s'�X;�OI��&�Zxe ���m�� p��ˀ�3s�O�O��O�O�O�aa�_т� |��q�d@��.v��.v��d@��[wFv��E����%s�t;B�w�t|�tP���PMA��QUa ��Q�8��1٠QTH�H{OLG�QHYS��3ES��qUE�pZB���Oτ�  ـP�ܐ(�A����v�!�t�O`�q��u�"���8FA��IROG�����Q2���o�"��p�^�INFOҁ�׃hV����R�H�OI���� (�0SLEQ ������Y�3����Á��P0Ow0��5�!E0NU���AUT�A�COPAY�=�/�'��@Mg��N��=�}1������ ���RG��Á���X_�P�$;ख�`
��W��P��@��������EXT_CY�C bHᝡRpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�H�SdB����2�$��F�p���GPLeAdA
�TAR �Б@���P�2��裔d� ,�0FL�`�o@YN��K�Mz��Ck��PWR+��9ᘐ��DELA4}�dY�pAD�a� �QSKIP4�� �A�$�OB`NeT�} ��P_$� M�ƷF@\bIpݷ�ݷ �ݷd����빸��@Š�Ҡ�ߠ�9���J2R� ��� m4V�EX� TQQ� ����TQ������ ���`�#�RDC�V� )�`��X)�R�p������r��m$RGE7AR_� IOBT�2�FLG��fipER��DTC���Ԍ���2�TH2NS}� S1���G T\0' ���u�M\Ѫ`qI�d��REF��1Á� l�h��E�NAB��cTPE �04�]����Y�]��� �Qn#��*��"�����
��2�Қ�߼�����(����3�қ'�9�K�]�o���4�Ҝ�������������5�ҝ!�3�E�W�i�{�
�6�Ҟ��������(�����7�ҟ-�?Qcu�8�Ҡ��������SWMSKÁ�l��aڝ�EkA��MO[TE6�����@0�݂TQ�IO}5�)IS�tR�W@��� �pJ����p�����E�"$DS?B_SIGN�1UQ��x�C\��S23�2���R�iDEVICEUS�XRSR�PARIT��4!O�PBIT�QI�O?WCONTR+�TQX��?SRCU� MpS�UXTASK�3Nx�p�0p$TATU�PK�S�0������p_XPC)�$F�REEFROMS8	pna�GET�0���UPD�A�2E#P|� :��� !$USAN�na&����ERI�0�Rp�RYq5*"_j@�P8m1�!�6WRK9K�D���6��QFRIgEND�Q�RUFg��҃�0TOOL�6M�Y�t$LENG�TH_VT\�FI!R�pC�@ˀE> +IOUFIN-RM���RGI�1ÐAIT�I�$GXñ3IvFG2v7G1���p3�BơGPR�p�1F�O_0n 0��!RE��p�53҅U�TC��3A�A��F �G(��":���e1n!��J�8�%����%]��%�� 74�OX O0�L��T�3H&��8���%b4J53GE�W�0�WsR�TD����T��M�����Q�T]�$V C2����1�а91�8��02�;2k3�;3 �:ifa�9-i�aQ���NS��ZR$V��2BVBwEV�	V�B;�����&�S�`��F�"�kX�@�2a�PS�E���$r1C��_$Aܠ6wPR��7vMU�cS�t '��529�G� 0G�aV`��p�d`���50�@��-��
25S�� �"�aRW����B�&�MN�AX�!�A:@�LAh��rTHIC¤1I���X�d1TF�Ej��q�uIF_C	H�3�qI܇7�Q�pG1RxV���]��:��u�_JF~�PR|ԀƱ�RVAT��� ��`���0R�榀DOfE��COU�Ա��AXI���O�FFSE׆TRIGNS���c����h������H�Y��IG#MA0PA�pJ�E��ORG_UNEV��J� �S������d �$CА��J�GROU����TqOށ�!��DSP���JOGӐ�#��_Pӱ�"O�q����@�&7KEP�IR��ܔ2�@M}R��AP�Q^��Eh0��K�SYS��q"K�PG2�BRAK�B��߄�pY�0=�d����`AD_������BSOC���N���DUMMY14�p@SV�PDE_�OP�#SFSPD�_OVR-���C���ˢΓOR٧3N�]0ڦF�ڦ��OV���SF��p���F�+�r!���CC��1q"L�CHDL��REC�OVʤc0��Wq@M������RO�#��Ȑ9_+��� @0�e@�VER�$OF�Se@CV/ �2WD��}��Z2���T�R�!���E_F�DO�MB_CM4���B��BL�bܒ#��adtVQR�$0pd���G$�7�AM5�`�� eŤ��_M;��"'����8$CA�'�E�8�8$HB�K(1���IO<�8����QPPA�������
��Ŋ����DVC_DBhC;��#"<Ѝ�r!S�1[ڤ�S�y3[֪�ATIOq 1q� ʡU�3���CABŐ�2�CvP���9P^�B���_� �S�UBCPU�ƐS �P �M�)0NS�c�M�"r�$HW_AC��U��S@��SA�A~�pl$UNITm�l_�AT���e�Ɛ�CYCLq�NEC�A���FLTR_2_FIO�7(��)&�B�LPқ/�.�_S[CT�CF_`�Fb�l���|�FS(!E�e�CHA�1��4�D°"3�RSD��$"}�����_Tb�PROX����� EMi_��ra�8!�a !�̹a��DIR0�RAOILACI�)RMr�CLO��C���Qq���#q�դ�PR=�S��AC/�c 	���FUNCq�0rRINP�Q�0��2�!3RAC �B ��[8���[WARn���#BL�Aq�A�����DAk�\���LD0���Q��q2eq�TI"r8��K�hPRIA�!r"AF��Pz!=�;���?,`�RK���MǀI�!�DF_@B�%1�n�LM�FAq@H�RDY�4_�P@R�S�A�0� �MUL�SE@���a ���ưt��m�m$�1$�1$1�o����� x*�EG00����!cAR���Ӧ�09�2�,%� 7�AXE��RKOB��WpA��_l-���SY[�W!‎&S&�'WRU�/-1��@��STR������Eb� 	�%��J��A�B� ���&9�����O�To0 	$��A�RY�s#2��Ԓ�	�ёFI@��$LGINK|�qC1�aI_�#���%kqj2XYZ��t;rq�3�RC1j2^8'0B���'�4����+ �3FI���7�q����'���_Jˑ���O3�QO�P_�$;5���AT�BA�QBC��&�D�Uβ�&6��TURN߁"r�E11:�p��9GFL�`_���* �@�5�*7��Ʊ 1��� KŐM��&8����"r��ORQ ��a�(@#p=�j��g�#qXU�����mTOVEtQ:�M��i�� �U��U��VW�Z�A �Wb��T{�, ��@;� uQ���P\�i��UuQ�W`e�e�SERʑ
e	��E� O���UdAas��4S�/7����AX��B�'q ��E1�e��i��irp �jJ@�j�@�j�@�jP �j@ �j�!�f��i� �i��i��i��i� y�y�'y�7yTq�HyDEBU8�$ 32���qͲf2G �+ AB����رnSVS�7� 
#�d�� L�#�L��1W��1W�JA W��AW��AW�QW�@!�E@?D2�3LAB��29U4�Aӏ��C 7 o�ERf�5�� � $�@_ A6��!�PO��à��0#�
�_MRA�t�� d � T��ٔERR����;STY&���I��V�0��cz�TOQ�d�PL�[ �d�"��	��C�! � pp`T8)0���_V1Vr�a(Ӕ����2ٛ2�E�ĺ��@�H�E���$QW�����V!��$�P��o�cI��a�Σ	 HELL_�CFG!� }5��B_BASq��SR3��� �a#Sb���1�%���2��3��4��5*��6��7��8����RO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CYO. U�OUG�P~ �����m�������TPհ_KAR�l�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h��]��l0SEM�4�(�Ml4�6�TYN�SO���DIZ�~�A������m_TM�MAN�RQ��k0E�����$KEYSWIT�CH���m���HE���BEAT��EF- LE~�����U���F!Ĳ���B�O_H�OM=OGREFUPPR&��y!� [��C��O��-ECO�C��Ԯ0_IOCMxWD
�a�'(k��� � Dh1���	UX���M�βgPgC�FORC�����O}M.  � @�T5(�U�#P, 1�֔, 3��45 �SNPX_ASt�w� 0��ADD�о�$SIZ���$VAR���TI�P/�.��A�ҹ�M�ǐ��/�1�+ U"S��U!Cz���FRI	F��J�S���5Ԓ��NF�Ѝ� � mxp`SI��TE�C\���CSGL��TQ2��@&����� ��S'TMT��,�P �&�BWuP��SHOW�4���SV�$��� �Q�A00 �@Ma}���� ��ਅ�&���5��6��7*��8��9��A��O ����Ѕ�Ӂ���0��F ��� G��0G���0 G���@G��PG��U1	1	1	1+	U18	1E	2��2��U2��2��2��2��U2��2��2��2��U2	2	2	2+	U28	2E	3��3��U3��3��3��3��U3��3��3��3��U3	3	3	3+	U38	3E	4�4��U4��4��4��4��U4��4��4��4��U4	4	4	4+	U48	4E	5�5��U5��5��5��5��U5��5��5��5��U5	5	5	5+	U58	5E	6�6��U6��6��6��6��U6��6��6��6��U6	6	6	6+	U68	6E	7�7��U7��7��7��7��U7��7��7��7��U7	7	7	7+	e78	7E��VP���UPDs�  ��`NЦ�5�YSL}Ot�� � L�`��d���A�aTA�80d��|�ALU:ed��~�CUѰjgF!aIgD_L�ÑeHI�j�I��$FILE_����d��$2�fS�A>�� hO��`E_BLCK��b$�>�hD_CPUyM�@yA��c�o�d��Y��ޅ�R �Đ
P�W��!� oqLA®�S=�ts�q~tRUN�qst�q~t���p�qst�q~t �T���ACCs��Xw -$�qLEN;� �tH��ph�_�I��ǀLOW_AXI�SF1�q�d2*�MZ���ă��W�Im�ւ�a�R�TOR��pg�Dx�Y���LACEk��ւ�pV�ւ~�_MA�2�v�������TCV��؁��T��ي���@��t�V����V�Jj�R�MA�i�J��m�u�)b����q2j�#аU�{�t�K�JK��V�K;���H���3��J�0����JJ��JJ��AAL��ڐ��ڐ�Ԗ4Օ5���N1����ʋƀW�LP�_�(�g�,��pr��{ `�`GROUw`���B��NFLI�C��f�REQUI;RE3�EBU��qB���w�2����p��x�q5�p�� \��/APPR��C}�Y��
ްEN٨CLO7��S_M��H����u�
�qu�� ���MC�����9�_MG��C�Co��`M��в�N�BRKL�N�OL|�N�[�R��_CLINђ�|�=�J����Pܔ�����������������6ɵ�̲�8k�D�����# ��
��q)��7�PATH3�L�BàL��H�wࡠ�J�CN�CA�Ғ�ڢB�IN�rUCV�4a��-C!�UM��Y,����aE�p����ʴ�~��PAYLOA���J2L`R_AN�q�Lpp���$��M�R_F2LSHR��N�LOԡ�R����`ׯ�ACRL_@G�ŒЛ� ��Hj`�߂$HM���FL�EXܣ�qJ�u� :�����׀�������1�F1�V�j�@�R�d�v�������E����ȏڏ ����"�4�q���6� M���~��U�g�y����T��o�X��H��� ���藕?�����ǟ ِݕ�ԕ����%��7��P��J�� � �V�h�z���`AT؃採@�EL�� �S��J|�Ŝ�JE�y�CTR��~�TN��FQ��HAND_VB-���v`�7� $��F2M�����ebSW�q�'��?� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)F�QAW�Z`i�Aw�A��PX X�'pi�Dw�D��ePf�G�p�)STk�h�!x��!N��DY�p נM�9$`%Ц�H�� H�c�׎���0� ��Pѵڵ�������t��J��� ����1��R�6��QAS�YMvř���v��pJ���cі�_SH>� �ǺĤ�ED����������J�İ%��C�I\Dِ�_VI�!X|�2PV_UNIX�FThP�J��_R�5_R c�cTz�pT�V��@��� İ�߷��U ��������Hqpˢ���aEN�3�DI����O4d �`J��� x g"IJAA �az�aabp�coc�`a��pdq�a� ��OMME��� �b�RqAT(`PT�@� S��a7�;�Ƞ�@�h�a��iT�@<� $�DUMMY9Q�o$PS_��RFC�vE`$v � 8���Pa� XƠ����STE���SB}RY�M21_VF�8$SV_ERF�qO��LsdsCLRJtEA��Odb`O�p� � D $�GLOBj�_LO ���u�q�cAp�r�@awSYS�qADR`�`�`TCH  �� ,��ɩb�W_NA���7�Ac��TSR���l ���
*?�& Q�0"?�;'?�I)?�Y) ��X���h���x����� �)��Ռ�Ӷ�;��Í�v�?��O�O�O�D�XOSCRE栘p�����ST��s}Hy`���Ea/_H�A�q� TơgpTYP�b���G�a�G���Od0ISb_䓀d�UEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI@m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1 �ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���>�VSHIF��Nc�P�`ג�E�ȐyR����OSUR��=Wk`RADILѮ��_�a��:�9a��`a��r��LULQ$O�UTPUT_BM����IM�AB �@��rTILSC	O��C7��� ����&��3��A����q���m�I�2 G���q�y@Md�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM���F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? �4�ZABC%��  $�"R���
E`�$$CLA}S������!�E`4�� � VIRT8]��/ 0ABS�����1 5�� <  �!F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o �$6HZi{0-�A�XL�p��"�63  �{tIN��qztGPRE�����v�p��uLARMRECOV 9�rwt�NG�� .;	 A   �.�0�PPLIC��?�5�p�H�andlingT�ool o� 
�V7.50P/2�3-�  �Pfv��
��_SWt�w UP�!� x�#F0��t���A� v� 864��� �it�y� r�2 7wDA5�� �� ?Qf@ϐo��Noneisͅ�˰ ��T��~�!LAex>�E_l�V�uT��s9�UTO�"�Њt�y��?HGAPON
0g��1��Uh�D 1581����̟�ޟry����Q 1���p�,�蘦����;�@��q_��"{�" �c��.�H���D�HTTHKYX��"� -�?�Q���ɯۯ5��� �#�A�G�Y�k�}��� ����ſ׿1����� =�C�U�g�yϋϝϯ� ����-���	��9�?� Q�c�u߇ߙ߽߫��� )�����5�;�M�_� q�������%��� ��1�7�I�[�m�� ��������!���� -3EWi{�� ����)/ ASew���� /��/%/+/=/O/ a/s/�/�/�/�/?�/ �/?!?'?9?K?]?o? �?�?�?�?O�?�?�?0O#O]���TO�E��W�DO_CLEA�N��7��CNM  � �__�/_A_S_�DSPDgRYR�O��HIc��M@�O�_�_�_�_o o+o=oOoaoso�o�o0���pB��v �u����aX�t������9�PLUGG���G��U�WPRCvPB�@��_�orOr_7�/SEGF}�K[mw xq�O�O�����?rqLAP�_�~q� [�m��������Ǐُ�����!�3�x�TO�TAL�f yx�USWENU�p�� �H����B��RG_STRING 1u��
�Mn�S�5�
ȑ_ITE;M1Җ  n5��  ��$�6�H�Z�l�~� ������Ưد����� �2�D�I/O SIGNAL̕�Tryout� ModeӕI�np��Simul�atedבOu�t��OVER�R�P = 100�֒In cyc�l��בProg� Abor��ב~��StatusՓ�	Heartbe�atїMH F�aul��Aler'�W�E�W�i�{ύ���ϱ�������  �CΛ�A����8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|���WOR{pΛ��(� ������ ��$�6�H� Z�l�~���������������� 2PO ̛�X ��A{�� �����/ ASew�����SDEV[�o �#/5/G/Y/k/}/�/ �/�/�/�/�/�/??�1?C?U?g?y?PALTݠ1��z?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O_�?GRI�`ΛDQ �?_l_~_�_�_�_�_ �_�_�_o o2oDoVo�hozo�o�o�o2_l�R ��a\_�o"4F Xj|����� ����0�B�T��oPREG�>�� f� ��Ə؏���� �2� D�V�h�z��������ԟ���Z��$AR�G_��D ?	����;���  	$�Z�	[O�]O���Z�p�.�SBN_C�ONFIG �;�������CI�I_SAVE  �Z�����.�TC�ELLSETUP� ;�%HO�ME_IOZ�Z�%MOV_��
��REP�lU�(�UT�OBACKܠ���FRA:\z� \�z�Ǡ'`�z���ǡi�WINI�0z����n�MESSAG༠�ǡC���ODEC_D������%�O��4�n�PAUSX!��;� ((O >��ϞˈϾϬ����� �����*�`�N߄��rߨ߶�g�l TSK�  wͥ�_�q�UgPDT+��d!�~A�WSM_CF���;���'�-�G�RP 2:�?� �N�BŰA��%�XS�CRD1�1
7� �ĥĢ������ ����*�������r� ����������7���[� &8J\n��|*�t�GROUN�|UϩUP_NA��:�	t��_E�D�17�
 ��%-BCKED�T-�2�'K�`����-t�z��q�q�z���2 t1�����q�kp�(/��ED3/ ��/�.a/�/;/M/ED4�/t/)?�/.p?p?�/�/ED5`? ?�?<?.�?O�?�?ED6O�?qO�?.pMO�O'O9OED7�O `O_�O.�O\_�O�O�ED8L_,�_�^�-�_ oo_�_ED!9�_�_]o�_	-9o�oo%oCR_  9]�oF�o�k� � ?NO_DEL���GE_UNUSE���LAL_OU�T ����W?D_ABORﰨ~���pITR_RT�N��|NONS�k���˥CAM�_PARAM 1�;�!�
 8
�SONY XC-�56 23456�7890 �~��@���?��( А\�
����{����^�HR5pq�̹��ŏR57ڏ��Aff��K�OWA SC31�0M
�x�̆�d @<�
��� e�^��П\�����*�<��`�r�g�CE�_RIA_I�j!�=�F��}�vz� ��_LIU�Y]�����<���FB�GP 1��Ǯ�M�_�q��0�C*  ����CU1��9��@��G��Z�CR�C]��d��l��s��R�����U[Դm��v����}����� C���ő(�����=�HE�`ONFIǰ�B��G_PRI 1�{V���ߖϨϺ�����������CHK�PAUS�� 1K� ,!uD�V�@� z�dߞ߈ߚ��߾��� ���.��R�<�b���O��������_MOR�� =�^Biq-���� 	 �����*�@�N�`�������$?��q?;�;����)K��9�P���ça�-:���	�

��M���pU��ð��<��,~��D�B���튒)
m�c:cpmidb1g�f�:�0���+¥�p�/�_  �(��(���� �s>��pY�pZU��?􌐨�Ug�/���p�W�f�M/w�O/�
DE�F l��s)��< buf.txAts/�t/��ާ��)�	`�����=L����*MC��1�����?43��1���t�īCz  �BHH�CPUeB��_B�y;���>C���C�nY
K�E?{�hD]^Dْ�?r���1D���^�=G	��F���F��C�m	fF�O�F'�ΫY	���&w�K1���s���).�pT���BDw��M@x8��1Ҩ��̨�g@D�p@�0E�Y�1X�EQ��EJP F�E��F� G���=F^F E��� FB� H,�- Ge��H3�Y��:�  >�?33 ���~�  n8�~@��5�Y�E>�ðA��Y<7#�
"Q ����+_�'RSMOFSb�p�.8��)T1���DE ��F �
Q��;�(P  QB_<_��R����,	op6C4P�Y
s@E ]AQ�2s@C�0)B3�MaC{@@*cw���UT�pFPROG %�z�o�oig�I�q���v��ldKEY_TBL  �&�S�#� �	
��� !"#$�%&'()*+,�-./01i�:;�<=>?@ABC�� GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����vq���͓��������������������������������������������������?�������p`�LCK�l4�p`�`S�TAT ��S_AU_TO_DO����5�INDT_EN�B!���R�Q?�1�Ty2}�^�STOPb����TRLr`LET�E��Ċ_SCR�EEN �Z_kcsc��U���MMENU 1 ~�Y  <�l �oR�Y1�[���v�m� ��̟�����ٟ�8� �!�G���W�i����� ���ïկ��4��� j�A�S���w������ ��ѿ����T�+�=� cϜ�sυ��ϩϻ�� �����P�'�9߆�]� o߼ߓߥ�������� :��#�p�G�Y��� ���������$���� 3�l�C�U���y����� ������ ��	VY)��_MANUAL���t�DBCO[�R�IGڇ
�DBNUIM� ��B1 e
��PXWORK 1!�[�_U/4�FX�_AWAYz�i�GCP  b9=�Pj_AL� #��j�Y��܅ `�_�  1"�[ , 
�od�&/�~&lMZ�IdPx@|P@#ONTIMه�� d�`&�
��e�MOTNEN�D�o�RECOR/D 1(�[g2�/{�O��!�/ky "?4?F?X?�(`?�?�/ �??�?�?�?�?�?)O �?MO�?qO�O�O�OBO �O:O�O^O_%_7_I_ �Om_�O�_ _�_�_�_ �_Z_o~_3o�_Woio {o�o�_�o o�oDo�o /�oS�oL�o ����@��� +�yV,�c�u���� ����Ϗ>�P����� ;�&���q���򏧟�� P�ȟ�^������I� [����� ���$�6��������jTOL�ERENCwB����L�͖ CS_CFG )��/'dMC:\�U�L%04d.C�SV�� c��/#A� ��CH��z� �//.ɿ��(S�RC_OUT *����SGN �+��"��#�1�7-FEB-20� 18:5701�5-JANp�0:�51+ P/�Vt�ɞ�/.��f��pa�m��P�JPѲ��VERSION Y��V2.0.8�4,EFLOGIC� 1,� 	�:ޠ=�ޠL��PROG_ENB�\�"p�ULSk' �����_WRSTJ�NK ��"fEMO�_OPT_SL �?	�#
 	R575/#=������0�B����TO�  �ݵϗ��V�_F EX�d�%���PATH AY�A\�����5+�ICT�Fu-��j�#e�gS�,�STBF_TTS�(�	d���l#t!w�� MAU��\z�^"MSWX�.���4,#�Y�/�
! J�6%ZI~�m��$SBL_F�AUL(�0�9'TDIA[�1<�� ����1234567890
��P��HZl~ �������/� /2/D/V/h/�� P� ѩ�yƽ/ ��6�/�/�/??/? A?S?e?w?�?�?�?�?��?�?�?�,/�UMP����� �ATRp���1OC@PMEl�~OOY_TEMP?�È�3F���G�|D�UNI��.�YN_?BRK 2_�/��EMGDI_ST�A��]��ENC2_�SCR 3�K 7(_:_L_^_l&_�_��_�_�_)��C�A14 _�/oo/oAoԢ�B:�T5�K�ϋo ~ol�{_�o�o�o '9K]o��� ������#�5� �/V�h�z��л`~��� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� ��x���������ү� ����,�>�P�b�t� ��������ο��� �(�f�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������:� �2�D� V�h�z�������� ����
��.�@�R�d� v�������������� *<N`r� ������ &8J\n��� �������/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?��?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_�_NoETMODE� 16�5�Q+ �d�X
X_j_�|Q�PRROR_P�ROG %GZ%��@��_  �UTA�BLE  G[�?oo)oRjRRS�EV_NUM  y�`WP�QQ�Y`�Q_AUTO_?ENB  �eOS��T_NOna 7�G[�QXb  *U��`��`��`��`�d`+�`�o�o�o�dH�ISUc�aOP�k_A�LM 18G[ e�A��l�P+�o�k}�����o_\Nb�`  G[�a��R
�:PTCP_V_ER !GZ!�_��$EXTLOGo_REQv�i�\�SIZe�W�TOoL  �aDzr��A W�_BW�D�p��xf́t�_D�I�� 9�5��d�T�asRֆSTE�P��:P�OP_�DOv�f�PFA�CTORY_TU�NwdM�EATU�RE :�5̀�rQHand�lingTool� �� \sfm�English� Diction�ary��rodu�AA Vis��� Master�����
EN̐n�alog I/O�����g.fd̐u�to Softw�are Upda�te  F OR��matic B�ackup��H5�96,�gro�und Edit�ޒ  1 H5Camera�F��OPLGX�e�ll𜩐II) nX�ommՐshw�n��com��co����\tp���pa�ne��  opl���tyle se�lect��al �C��nJ�Ցoniwtor��RDE���tr��Reli�ab𠧒6U�Diagnos(�푥��5528�u��h�eck Safe�ty UIF��E�nhanced �Rob Serv>%�q ) "S�r�User Fr[������a��xt. oDIO �fiG�s sŢ��endx��Err�LF� p$Ȑĳr됮� �����  !��FCTN_ Menu`�v-��ݡ���TP In�ېfac�  E�R JGC�p�בk Exct�gޠ�H558��ig�h-Spex�Sk�i1�  2
P���?���mmunic'�ons��&�l��ur�ې��ST xǠ��conn���2��TXPL��n{cr�stru�����"FATK�AREL Cmd�. LE�uaG�5�45\��Run-�Ti��Env��dG
!���ؠ++��s)�S/W��[��License�Z��� 4T�0�ogBook(Syڐ�m)��H54O�M�ACROs,\�/�Offse��Lo�a�MH������r�, k�MechS�top Prot����� lic/�M=iвShif����ɒMixx��)����xStS�Mode Switch��7 R5W�Mo�:�=.�� 74 ����g��K�2h�ul�ti-T=�M���L�N (Pos�Regiڑ�������d�ݐt Fun��ǩ�.�����Nu�m~����� lne���ᝰ Adju�p�����  - =W��tatuw᧒}T�RDMz��ot��scove
 U�9���3����uest 49�2�*�o�����62~;�SNPX b Ҟ��8 J7`���Lgibr��J�48��D�ӗ� �Ԅ�
�6O��� Parts in VCCMt�32���	�{Ѥ�J�990��/I� �2 P��TMILKIB��H���P��AccD�L�
T�E$TX�ۨ�ap�1S�Te����pkCey��wգ�d���Unexce{ptx�motnZ�0�������є��� O���� 90�J�єSP CSX�C<�f��Ҟ� P�y�We}���PRI��>vr�t�me�n�� ��iP�ɰa�����vGr{id�play�İv��0�)�H1�M�-10iA(B2�01 �2\� 0�\k/�Ascii��l�Т�ɐ/�Coyl��ԑGuar�� 
�� /P-�ޠ"�K��st{Patt ��!S�Cyc�҂�orie��I�F8�ata- qu�Ґ�� ƶ��mH5�74��RL��am����Pb�HMI �De3�(b����P�CϺ�Passw�o+!��"PE? S1p$�[���tp��� �ven��Tw�N�p��YELLOW sBOE	k$Arc��'vis��3*�n0�WeldW�cia�l�7�V#t�Opd����1y� 2F�=a�portN�(�p�T1�T� �� f��xy]�&TX��tw�igj�1� b�� ct\�JPN� ARCPSU cPR��oݲOL� wSup�2fil� p&PAɰאcro�� "PM(����O$�SS� eвtexF�� r���=�t�OssagT��P���P@�Ȱ�锱�r�tW��H'>r�dp9n��n1
t�!� z ��ascbin4psyn���+Aj�M HEL��NCL VIS� PKGS PL;OA`�MB �,��4VW�RIPE� GET_VAR� FIE 3\t���FL[�OOL:� ADD R72�9.FD \j8�'�CsQ�QE��DV�vQ�sQNO WT�WTE��}PD  �^��biRFOR ��ECTn�`���ALSE ALA�fPCPMO-130  M" #h��D: HANG �FROMmP�AQf�r��R709 D�RAM AVAILCHECKSO!���sQVPCS S�U�@LIMCHK� Q +P~dFF P�OS��F�Q R5�938-12� CHARY�0�P?ROGRA W��SAVEN`AME.�P.SV��7��$�En*��p?FU�{�T�RC|� SHAD�V0UPDAT K�CJўRSTATI��`�P MUCH �y�1��IMQ MOTN-003���}�ROBOGUI�DE DAUGHp�a���*�tou�����I� Šhd�AT�H�PepMOVET��ǔVMXPAC�K MAY AS�SERT�D��YC�LfqTA�rBE ?COR vr*Q3r�AN�pRC OP�TIONSJ1vr�̐PSH-171ZZ@x�tcǠSU1��1Hp^9R!�Q�`_TP�P��'�j�d{t�by app w�a 5I�~d�PHI����p�aTEL�MXSPD TB5b�Lu 1��UB6@�qEmNJ`CE2�61���p��s	�may 1n�0� R6{�R�} �Rtraff)��� 40*�p��f�r��sysvar scr J7��cj`DJU��bH� V��Q/�PSET� ERR`J` 6�8��PNDANT� SCREEN UNREA��'�J`MD�pPA���pR`�IO 1���PFI��pB�pGROUN�PD��G��R�P�QnRSVIP !p�a�P�DIGIT VE�RS�r}BLo�UE�Wϕ P06  �!��MAGp�ab�ZV�DI�`� S�SUE�ܰ�EP�LAN JOT` 'DEL�pݡ#Z�@=D͐CALLOb�Q� ph��R�QIP�ND��IMG�R�719��MNT/��PES �pVL�c��Hol�0Cq���t�PG:�`C�M�c�anΠ��pg.v~�S: 3D mK�view d�` L�p��ea7У�b� �of �Py���AN�NOT ACCE�SS M��Ɓ*�tn4s a��lok�^�Flex/:�Rmw!mo?�PA?��-�����`n�pa �SNBPJ AUTO-�06f����T|B��PIABLE1q� 636��PLN�: RG$�pl;pNnWFMDB�VI��>�tWIT 9x�0@o��Qui#0�ҺP�N RRS?pUS�B�� t & r/emov�@ )�_�v�&AxEPFT_=�� 7<`�pP:�O�S-144 ��h� s�g��@OST�� � CRASH� DU 9��k$P�pW� .$��_LOGIN��8&��J��6b046 i�ssue 6 J�g��: Slow� �st��c (�Hos`�c���`I�L`IMPRWtSPOT:Wh:0�T��STYW ./�VM�GR�h�T0CAT.��hos��E�q�T�� �O�S:+p�RTU' k�-S� ,����E:��pv@�2��� t\hߐ��m� ��all��0� 9 $�H� WA͐���3 CNT0 T��� WroU�al�arm���0s�d �� �0SE1���r R{�OMEBp���K�7 55��REàSE�st��g   �  �KANJI��no���INISITALIZ-p��dn1weρ<��d�r�� lx`�SC�II L�fai/ls w�� ��`�YSTEa���o��PNv� IIH���1W��Gro>Pm ol\wpSh@�P��Ϡ?n cflxL@А�WRI �OF Lhq��p?�F�up��de-rela�_d "APo SY��ch�Abetwe>:0IND t0$FgbDO���r� `��GigE�#op�erabilf  �PAbHi�H`��c�l�ead�\etfp�Ps�r�OS 0�30�&: fig��GLA )P ��i��}7Np tpswx�-B��If�g�������5aE�a EX�CE#dU�_�tPCL{OS��"rob�+NTdpFaU�c�!����PNIO V750�Q1��QaN��DB ��P M��+P�QED�DET���-� \rk��O�NLINEhSBU�GIQ ߔĠi`Z�I�B�S apABC? JARKYFq�9 ���0MIL�`� �R�pNД �p0G+AR��D*pR��PN�"! jK�0cT�P�Hl#n�a�ZE }V�� TASK�$VP2(�4`
�!�$��P�`WIBPK0�5�!FȐB/��B�USY RUNN��� "�򁐈��R�-p�LO�N�DI�VY�CUL��f3sfoaBW�p����30	V��ˠIyT`�a505.�@{OF�UNEX�P�1b�af�@�E��S�VEMG� NML�q� D0pCC_SGAFEX 0c�08"q]D �PET�`N@N�#J87����RsP��A'�M�K�`K��H GUNCH�G۔MECH�pM�c� T�  y, �g@�$ ORY L�EAKA�;�ޢS�PEm�Ja��V�tG�RIܱ�@�CTLN�TRk�FpepnR�j50�EN-`#IN�����p �`�Ǒk!��T3/dqo��STO�0A�#�L��p �0�@�Q�АY0�&�;pb1TO8pP�s���FB�@Yp`�`DU��aO�supk��t4 � P�F� Bn�f�Q�PSVGN-q1��V�SRSR)J�UP�a2�Q�#D��q l O��QBRKCTR5Ұ�|"�-�r�<pc�j!IN=VP�D ZO� ���T`h#�Q�cHset�,|D��"DUAL�� w�2*BRVO1/17 A]�TNѫt8�+bTa2473��q.?��sAUz�i�B��complete���604.� �-�`hanc�U�� F��e8�� 	 ��npJtPd!q��`���� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP���R(}\xPe� aʰI���E��1��p�� j  �� xSt�'^t �A�AxP�q\ 5 sig��a��"AC;a��
�b�CexPb_p��.p�c]l<bHbcb_c�irc~h<n�`tl 1�~`xP`o�dxP�b]o2�� �cb�c�ixP>�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`>�cptlibxzxP�lcr�xrxP\�b�lsazEdxP_fm �}gcxP�x���o|sp��o�mc(��ob_jDzop�u6�wf���t��wms�1q��s1ld�)��jmc�o\��n��nuhЕ��|st�e��>�pl�qp�iwcck���uvf0uxߒ��lvisn��CgaculwQ
E� F  ! Fc.sfd�Qv�� qw����Data Ac_quisi��nF�<|1�RR631`��T}R�QDMCM ��2�P75H�1�P5k83xP1��71��k59`�5�P57<P xP�Q����(���Q̖�o pxP!da�q\�oA��@��y ge/�etdms�?"DMER"؟,�GpgdD���.�m��8�-��qaq.<᡾FxPmo��h���f{��u�`13��MACR�Os, Sksaf�f�@z����03�SR��Q(��Q6��1�Q9�ӡ�R�ZSh��PxPJW643�@7ؠ6�P,�@�PRS�@���e x�Q�UС PIK�Q52 PTLC�W���xP3 (��p/O��!�Pn �xP�5��03\sfm�nmc "MNM�Cq�<��Q��\$AcX�FM���ci,Ҥ��X����cdpq+�
�s�k�SK�xP�SH560,P��,�y��refp "RE�Fp�d�A�jxP	�o�f�OFc�<gy�to�TO_����ٺ���+je�u��caxis2�xPE��\�e�q"ISDT�c��]�prax ���MN��u�b�isde܃h�\�w�xP�! isbasi5c��B� P]��QoAxes�R6��8����.�(Ba�Q�ess��xP����2�D�@�z�atis ���(�{�����~��m��FMc�u�{�<
ѩ�MNIS��ݝ ����x����ٺ���x� j75��De�vic�� Interfac�RȔQJ754��� xP�Ne`��xP�ϐ`2�б����dn� �"DNE���
t�pdnui5UI��ݝ	bd�bP>�q_rsofOb~
dv_aro��u�����stchkc��z	 �(�}onl��G!ffL+H�J(��"l"�/�n�b��z�h�amp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!�2��xpc_2pcc{hm��CHMP_�|8бpevws��2�쳌pcsF��#C� SenxPacrao�U·�-�R6�P�d�xPk�����p��g8T�L��1d M�2`���8�1c4ԡ�3 qem��GEM,\i(�>�Dgesnd�5��`�H{�}Ha�@sy����c�Isu�xD��Fmd��I��7�4���u����AccuCal �P�4� ��ɢ7ޠBU0��6+6f�6��C99\aFF q�S(�U��2�
X�p�!Bdf��cb_�SaUL��  �� ?�ܖt�o��otplus\tsrnغ�qb��Wp��t���1��T�ool (N. �A.)�[K�7�Z�(P�m����bfc�ls� k94�"Kp4p��qtpap�� "PS9H�stpswo��p�L7��t\�q����D�yt 5�4�q��w�q��� ��M�uk��rkey�����s��}t�sfoeatu6�EA��� cf)t\Xq�����̜d�h5���LR0C0�md�!�587���aR�(����2V���8c?u3l\�pa�3}H�&r-�Xu���t,�� �q "�q�Ot� �~,���{�/��1c�}����y�p�r��5� ��S�XAg�-�y���W�j874�- i�RVis���Queu�� Ƒ�-�6H�1���(����u����tӑ����
�tp�vtsn "VTCSN�3C�+�� v\p�RDV����*�pr�dq\�Q�&�vs�tk=P������n�m&_�դ�clrq8ν���get�TX��Bd���aoQϿ�0qstr�D[� ��at�p'Z����npv��@�enlIP0��`D!x�'�|���sc ����tvo/��2�q���vb����q ���!���h]��(�� Control^�PRAX�P5��g556�A@59�P[56.@56@5A��J69$@982� J552 IDVR7�hqA���16��H���La�� ���Xe�frlpa�rm.f�FRL��am��C9�@(F�����w6{���A<��QJ643�� �50�0LSE
�_pVAR $SG�SYSC��RS_?UNITS �P�2��4tA�TX.$V�NUM_OLD �5�1�xP{�50�+�"�` Funct���5tA� }��`#@��`3�a0�cڂ��9���@H5נ� �P���(�A����۶�}����ֻ}��bP�Rb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`��2�1���96����@�%C�� Aف��J�bIncr�	����\����1o5qni4�MNINp	xP�`���!��Hour�  � �2�21 ��AAVM���0y ��TUP ��J545 ���6162�V�CAM  (��CLIO ���R6�N2�MS�C "P ��STYL�C�2�8~ 13\�NRE "FHRM �SCH^�DC�SU%ORSR �{b�04 �oEIOC�1 j o542 � os| ~� egist������7�1��MASK�93�4"7 ��OCO) ��"3�8��12���� 0 HB���� 4�"39N� �Re�� �LCH=K
%OPLG%��3"%MHCR.%M�C  ; 4? ��6 6dPI�54�s� �DSW%MD� pQ�K!637�0�0p"��1�Р"4 �6~<27 CTN K V� 5 ���"7���<25�%/�T�%FRDM� �Sg!���930 FB( NB�A�P� ( HLB o Men�SM$@<jB( PVC ��s20v��2HTC�~CTMIL��~\@PAC 16U��hAJ`SAI \@EL�N��<29s�U�ECK �b�@FR3M �b�OR����IPL��Rk0CS�XC ���VVF�naTg@HTTP ��!26 ��G��@obIGUI�"%IPGS�r� H863 qb�!�07rΈ!34 �r�84 \so`! Qx`CC�3 Fb�21�!9s6 rb!51 ����!53R% 1!s(3!��~�.p"9js �VATFUJ775�"��pLR6^RP�W;SMjUCTO�@xT158 F!80���1�XY ta3!770� ��885�UO	L  GTSo
�{` �LCM �r| TS�S�EfP6 W�\@C�PE `��0VR�� l�QNL"��@001 imrb�c3 =�b�0���0�`�6 w�b-P- Ru-�b8n@5EW�b9 �Ґa� ���b�`�ׁ�b2 2000$��`3��`4*5�`A5!�c�#$�`7.%~�`8 h605? ;U0�@B6E"aRpm7� !Pr8 t��a@�tr2 iB�/�1vp3�vp5 �Ȃtr9Σ�a4@-�p�r3 F��r5`&�re`u��r7 ��r8�U�p9 \h�738�a�R2DK7"�1f��2&�y7� �3 7iCЊ�4>w5Ip�Or6�0 C�L�1bEN�4 I�pyL�uP��@LN�-PJ8�N�8Ne�N�9 H�r`�E"�b7]�|���8�В����9 2��a`0�qЂ5�%U097 0��@1�0����1 (�q�3 5R���0���mpU��0�0�7*�H@x(q�\P"RB6�q124�b;��@���f@06� x�3 p�B/x�u ��x�6 /H606�a1� ����7 6 ���<p�b155 ����}7jUU162 ��3 g��4*�6?5 2e "_��PF�4U1`���B1��z�`0'�174 �q���P�E186 R� ��P�7 ��P�8�&�3 (�90 B/�s191����@�202��6 30���A�RU2� d���2 b2h`��4Ģ᪂2�4���19�v Q�2��u2d�TRpt2� ��H�a2hPd�$�5���!U2�pD�p
�2�p��@5�0H-@��8 @�9��TX@�� �e5�`rb26Af�2^R�a�2 Kp��1y�b5Hp�`

�5�0@�gqGA��F�a52ѐ�Ḳ6�K60ہ5� ׁ2��i8�E��9�EU5@�ٰ\�q5hQ`S�2
ޖ5�p\w�۲�pJh �-P��5�p1\t�ZH�4��PCH�7j��phiw�@��P�x�~�559 ldu�  P�D���Q�@�������� �`.��P>��8��581�"�q58�!AM۲T�A iC�a589��@�x�����5 �a��12@׀0.�1���,�2��8��,�!P\h8��Lp� ��,�7��6�08�40\� ANRS 0C}A��p��{��ran��FRA ��Д�е���A% ���ѹ�Ҍ�����( ����Ќ���З��� ������ь����$�!G��1��ը���������� xS�`q�  �����`�64��M��iC/50T-H������*��)p46��� C���N����m75s�֐� Sp��b4�6��v����ГM-71?�7�З�����42������C��-��а�70�r�E��/h����O$���rD���c7c7C@�q��Ѕ���L���/��2\imm7c7�g������`���(��e����� "�������a r�L�c�T,�Ѿ�"��,�� ��x�Ex�m77t����k���a5�����)�iC��-HS-� B
_�@>���+�Т�7U��]���Mh7�s�7������-9~?�/260L_� �����Q������4��]�9pA/@���q�S�х鼔��h621��c��92������.�)92c0�g$�@ �����)$��5$����pylH"O"
�21p���t?�350� ���p��$�
��� �350!���0���9�U/0\m9��M9A3��4%� s��3M$��X%yu���"him98 J3����� i d�"m4~�103p�� ����h794̂�&R���H�0����\���g� 5AU��՜��0���*2@��00��#06�`�АՃ�է!07{r ��������kЙ @����EP�#�� ����?��#!�;&�07\;!�B1P��߀A��/ЁCBׂ2��!�:/��?�ҽCD2C5L����0�"l�2BL
#��B��\20�2_�r�re ���X��1��N����A$@��z��`C�p0U��`��04��DyA�\�`fQ����sU���\�5  ���� p�^t��<$85���+�P=�ab1l��1LT��lA8�!uDnE\(�20T��J�1 e�bH85���b����5[�16Bs��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3� � ��b�s��-`�_�Wa8�_����6I	$2�X5�1�U85��R�p6S����/�/+q��!�q��`�6o��58m[o)�m6sW��Q��?��set06�p ��3%H�5��10�p$����g/�JrH~��  ��A�856����F�� ���p/2��h�܅�✐)�5��̑v0��(��m6��Y�!H�ѝ̑m�6�Ҝ���a6�DM����-S�+��H2������ ��� �r̑��✐0��l���p1���Fx���2�\t6h T6H����Ҝ�'V l���ᜐ�V7ᜐP/����;3A7��@p~S��������4�`@圐�V���!3��2�PM[��%ܖO�7chn��vel5�p���Vq���_arp#���̑�.���2l_�hemq$�.�'�6415���5���?�� ��F�����5g�L�ј[���1��𙋹y1����M7NU�@�М��eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h����� �u���㜐��`ZS�!ܑ4���M-����S�$̑�ք �� �0��<�����07shJ�H�v�À�sF ��S*󜐳���̑�� �vl�3�A�T�#��`QȚ�Te��q�pr��,��T@75j�5�dd� ̑1�(UL�&�(�,����0�\�?���̑�a��? xSt���a��e�w�2��(�	�2�C��A/���\�+px�����21 (ܱ�CL S����B�̺��7F���?�<�lơ1L����c� ��b�u9�0����e/q���O���9�K��r9 (��,�Rs�ז�x5�G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O����1!41w���2<T@� _std��G��y� �ң�H� jdgm����w0\� �1 L���	�P�~�W*�b��t 5������%3�,���E{�������L��5\L��3�L�|#~���~!���4�#��O����h�L6A������2璥���44������[6\j4s��·���#��ol�E"w�8Pk�����?0 xj�H1�1Rr�>��6]�2a�2Aw�P ��2��|41�8��ˡ���{� �%�A<���  +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R� �ˑb�W���Fs��� �)�ѐ�!���a�1��ڛ�5��16�16�C��C����0\imBQ��d����b���\B5�-���DiL ���O�_�<ѠPEtL�E�RH�ZǠPgω�am1l��u���̑��b�<����<�$�T �̑�F����Ȋ�D�pb��X"�ᒢ��pw� ���^t���9�0\� j971\kckrcfJ��F�s�����c��e "CTME�r������!�a�`main.p[��g�`run}�_vc�#0�w�1O�ܕ_u����bctm�e��Ӧ�`ܑ�j7�35�- KAREL Use {�	U���J��1��
�p� Ȗ�9�B@���L�9��7j[�a�tk208 "KP��Kя��\��9���a��̹����cKRiC�a�o ��kc�q J�&s�����Grſ� fsD��:y��s��A1X3\j|хrdtB�,� ��`.v�q�� ��sǑIf�Wfj52��TKQuto S�et��J� H5nK536(�932�Z��91�58(�9�BA�1(�74O,A$�?(TCP Ak��В/�)Y� �\t�pqtool.v��v���! co�nre;a#�Control Re��ble��CNRE (�T�<�4�2���D�)����S�552��q(g�� (򭂯4X�cO�ux�\sfuts�UTS`�i�栜����t�棂��? 68�T�!�SA OO+D6���������,!��6c+� ig.t�t6i��I0�TW8 ���la��vo58�o�bFå򬡯i�Xh��!Xk�0Y!�8\m6e�!6EC���v��6���������<16�A���A�6s����U�g�TX|ώ���r1�qR��˔Z4�T�����,#�eZp)g����<O NO0���uJ��tCR;�x�F�a� xSt�f���prdsuchk �1��2&&?���	t��*D%$�r(��@���娟:r��'�s�q8O��<scrc�C�<\At�trldJ"�o�\�V����Pa�ylo�nfir1m�l�!�87��7� �A�3ad�! ��?ވI�?plQ��3���3"�q��x p�l�`���d7��l�calC�uDu���;���mov�����i'nitX�:s8O�p�a�r4 ��r67A4�|�e GenerGatiڲ���7g2�q$��g R� (#Sh��c ,|�bE��$Ԓ\�:�"��4��4�4�. sg��5�F$d6�"e�!p "SH�AP�TQ ngcr pGC�a(�&"<� ��"GDA¶��r6�"aW�/�$�dataX:s�"t�pad��[q�%tput;a__O7;a�o8(�1�yl+s�r�?�:H�#�?�5x�?�:c O��:y O�:�IO�s`O%g�qǒ�?�@08\��"o�j92;!�P�pl.Colli=s�QSkip#��@ 5��@J��D��@\ވP�C@X�7��7��|s2��ptclsF�LS�DU�k?�\_ ets�`�< \�Q��@���`dc�KqQ�FC;��J,�n��` (��4eN����T�{��� 'j(�c�q���/IӸaxȁ��̠H������зa�e\mc�clmt "CL�M�/��� mate�\��lmpALM0�?>p7qmc?����2vm�q��%�3s���_sv90�_x_m#su�2L^v_� K�o�{in�8(3r<�c_logr�N�rtrcW� �v_3�~yc��d��<�te��derv$cCe� Fiρ�R��Q�?�l�enter߄|��d(Sd��1�TX�+�fK�r�a99sQ9x+�5�r\tq\�� "FNDR����STDn$�LANG�Pgui��D⠓�S����Ơ�sp�!ğ֙uf �ҝ�s����$�����e+�=����������ࠓ���w�H�r\f�n_�ϣ��$`x�tc�pma��- TC�P�����R638� R�Ҡ��38
��M7p,���Ӡ�$Ӏ��8p0Р�VS,�>�tk��99�a��B3�� �PզԠ��D�2�����UI��t���hqB���8��������p���rqe�ȿ��exe@ 4φ�B���e38�ԡG��rmpWXφ�var@�φ�3N������vx�!ҡ��q��RBT $cO�PTN ask �E0��1�R MA�S0�H593/�9�6 H50�i�48
0�5�H0��m�Q�QK��7�0�g�Pl��h0ԧ�2�ORD�P��@"��t\mas��0�a��"�ԧ�����k�գR�����¹`m��b��7�.f���u�d��r��splayD�E���1>w�UPDT Ub���887 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q `�䗣�#��К�`2�� vlv��Ù�`$�>�b���! S���Easy/К�U�til��룙�51G1 J�����R7 Θ�Nor֠��inGc),<6Q�� �`�c��"4�[���98Q6FVRx So����q�nd6����P�� 4�a\ (��
  ����D���d��K�bdZ����men7���- Me`tyFњ�Fb¨0�TUa�57	7?i3R��\��5�u?��!� n����f������l\mh�Ц�űE|Ghmn�	��<\HO���e�1�� l!D��y��Ù�\|�p����B���Ћmh�@��:.aG! ���/�t�55�6�!X�l�.us��Y/k)�ensubL���eK�h�� �B\1;5�g?y?�?�?D��?*r�m�p�?Ktbox  O2K|?�G��C?A%�ds���?1ӛ#�  �TR��/��P�4B�`��U�P�V�P"�Q�P0@�U�PO��P�"�T3�U@�P�f�Pk"�2}�4�T@�P�f�P2�"�Q5�S��Q���R?Ă�Q3t.��P׀al��P+O�P517��IN�0a��Q(}g��PESTf3ua�PB�l��ig�h�6�aq��P? � xS��`�  n�0mbum�pP�Q969g�6!9�Qq��P0�baAp|�@Q� BOX��,>vche�s�>v�etu㒣=wffse�3���]�;u0`aW��:zol�sm�<ub�a-��]D�K�ibQ�c����Q<twaǂ� tp�Q҄Tar�or Recov�b�O�P�642 ����a�q��a⁠Q3Erǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>�pjot��PXc���C�1�adb -�ail��nag���b�QR629�a�Q��b��P  �
�  �P��$$C�L[q ���t������$�PS_DIGIT�.��"�!� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv��������*璬1:PRODUCT�Q0\PGSTK�bqV,n�99��\���$FE�AT_INDEX���~��� 搠ILECO_MP ;��)���"��SETU�P2 <�~��  N !��_AP2BCK� 1=�  #�)}6/E+%,/i/��W/�/~+/�/ O/�/s/�/?�/>?�/ b?t??�?'?�?�?]? �?�?O(O�?LO�?pO �?}O�O5O�OYO�O _ �O$_�OH_Z_�O~__ �_�_C_�_g_�_�_	o 2o�_Vo�_zo�oo�o ?o�o�ouo
�o.@ �od�o���M �q���<��`� r����%���̏[��� ����!�J�ُn��� ����3�ȟW������ "���F�X��|���� /���֯e������0� ��T��x������=� ҿ�s�ϗ�,ϻ�9��b�� P/ 2>) *.VRiϳ�!�*�������ߌ��PC�7�!�OFR6:"�c������T��߽�Lը���ܮx���*.F��>� �	N�,�k���ߏ��STM @�����Qа���!��iPendant Panel���H��F���4�������GIF��������u����JPG &P��<�����	PANEL1.DT��������2�Y�G��
3w�� ���//�
4�a/��O///�/�
T�PEINS.XM)L�/���\�/�/��!Custom Toolbar?��PASSWO�RD/�FRS�:\R?? %P�assword ?Config�?� �?k?�?OH�6O�?ZO lO�?�OO�O�OUO�O yO_�O�OD_�Oh_�O a_�_-_�_Q_�_�_�_ o�_@oRo�_voo�o )o;o�o_o�o�o�o* �oN�or��7 ��m��&��� \�����y���E�ڏ i������4�ÏX�j� �������A�S��w� ����B�џf����� ��+���O������� ��>�ͯ߯t����'� ��ο]�򿁿�(Ϸ� L�ۿpς�Ϧ�5��� Y�k� ߏ�$߳��Z� ��~�ߢߴ�C���g� ����2���V����� ����?����u�
� ��.�@���d������ )���M���q����� <��5r�%� �[�&�J �n��3�W ���"/�F/X/� |//�/�/A/�/e/�/ �/�/0?�/T?�/M?�? ?�?=?�?�?s?O�? ,O>O�?bO�?�OO'O �OKO�OoO�O_�O:_ �O^_p_�O�_#_�_�_ Y_�_}_o�_�_Ho)f��$FILE_D�GBCK 1=���5`��� ( �)
�SUMMARY.�DGRo�\MD:�o�o
`Dia�g Summar�y�o�Z
CONSLOG�o�o�a
J��aConsol�e logK�[��`MEMCHEC�K@'�o�^qM�emory Da�ta��W�)}�qHADOW���P��sSha�dow Chan�gesS�-c-�?�)	FTP=���9����w`qmme?nt TBD׏�W�0<�)ETHERNET̏�^�q��Z��aEthe�rnet bpfi�guration�[��P��DCSVR�Fˏ��Ïܟ�q%��� verif�y allߟ-c1�PY���DIFF�ԟ��̟a��p%��diffc���q¡�1X�?�Q�� �����X��CHGD��¯ԯi��p!x��� ���2`�G�Y�� ��� ��GD��ʿܿq��p8���Ϥ�FY3h�O�a��� ��(σGD������y��p��ϡ�0�UPDA�TES.�Ц��[�FRS:\������aUpdates� List���kP�SRBWLD.C	M.��\��B��_p�PS_ROBOWEL���_����o�� ,o!�3���W���{�
� t���@���d����� /��Se���� �N�r� = �a�r�&�J ���/�9/K/� o/��/"/�/�/X/�/ |/�/#?�/G?�/k?}? ?�?0?�?�?f?�?�? O�?OUO�?yOO�O �O>O�ObO�O	_�O-_ �OQ_c_�O�__�_:_ �_�_p_o�_o;o�_ _o�_�o�o$o�oHo�o �o~o�o7�o0m �o� ��V�z �!��E��i�{�
� ��.�ÏR�������� ��.�S��w������ <�џ`������+��� O�ޟH������8����߯n����$FI�LE_��PR����������� �MDON�LY 1=4�� 
 ���w�į ��诨�ѿ������� +Ϻ�O�޿sυ�ϩ� 8�����n�ߒ�'߶� 4�]��ρ�ߥ߷�F� ��j�����5���Y� k��ߏ���B����� x����1�C���g��� ����,���P����������?��Lu�VISBCKR�<�a�*.VD|�4 �FR:\���4 Vision� VD file � :LbpZ� #��Y�}/$/ �H/�l/�/�/1/ �/�/�/�/�/ ?�/1? V?�/z?	?�?�???�? c?�?�?�?.O�?ROdO O�OO�O;O�O�OqO _�O*_<_�O`_�O�_�_%_�_�MR_G�RP 1>4��L�UC4  B��P	 ]�ol`��*u����RHB ��2� ��� ��� ���He�Y�Q`o rkbIh�oJd�o�Sc��o�oLP�L�c`�J�gwF��5U�aS?��o�o E�]��F�nEwB��.��99��ߓ>�E}A%�'Az�/lq?�R4Az��xq�0~�� F@ �r�d�a}J��N�Jk�H9��Hu��F!��/IP�s}?�`��.9�<9���896C'�6<,6\b�1�,.�g�R���^x�PA�����|�ݏ x���%��I�4�F� �j�����ǟ���֟���!��E�`r�UBH�P �~��������W
6�P=��PQ��˯�o�o�B��P5���@�3�3@���4�m�,�@�UUU��U�~w�>u.�?!x��^��ֿ���3��=�[z�=�̽=�V6<�=�=�=$q��~���@8�i7�G��8�D�8@9!�7���@Ϣ���cD�@ D�� CϫoV��C��P��P'� 6��_V� m�o��To�� xo�ߜo������A� ,�e�P�b����� ��������=�(�a� L���p���������^� ������*��N9r ]������� �8#\nY� }�������/ ԭ//A/�e/P/�/p/ �/�/�/�/�/?�/+? ?;?a?L?�?p?�?�? �?�?�?�?�?'OOKO 6OoO�OHߢOl��ߐ� ���O�� _��G_bOk_ V_�_z_�_�_�_�_�_ o�_1ooUo@oyodo vo�o�o�o�o�o�o Nu�� �������;� &�_�J���n������� ݏȏ��%�7�I�[� "/�描�����ٟ�� �����3��W�B�{� f�������կ����� ��A�,�e�P�b��� �����O�O�O��O �OL�_p�:_������ ���������'��7� ]�H߁�lߥߐ��ߴ� ������#��G�2�k� 2��Vw�������� ���1��U�@�R��� v������������� -Q�u��� r��6��) M4q\n��� ���/�#/I/4/ m/X/�/|/�/�/�/�/ �/?ֿ�B?�f?0� BϜ?f��?���/�?�? �?/OOSO>OwObO�O �O�O�O�O�O�O__ =_(_a_L_^_�_�_�_ ���_��o�_o9o$o ]oHo�olo�o�o�o�o �o�o�o#G2k V{�h���� ���C�.�g�y�`� ���������Џ�� �?�*�c�N���r��� �����̟��)�� M�_�&?H?���?���? �?�?����?@�I�4� m�X�j�����ǿ��� ֿ����E�0�i�T� ��xϱϜ�������� �_,��_S���w�b߇� �ߘ��߼������� =�(�:�s�^���� �������'�9� � ]�o����~������� ������5 YD V�z����� �1U@yd ��v�����/Я */��
/�u/��/�/ �/�/�/�/�/??;? &?_?J?�?n?�?�?�? �?�?O�?%OOIO4O "�|OBO�O>O�O�O�O �O�O!__E_0_i_T_ �_x_�_�_�_�_�_o �_/o��?oeowo�oP� �oo�o�o�o�o+ =$aL�p�� �����'��K� 6�o�Z������ɏ�� 폴� ��D�/ / z�D/��h/ş���ԟ ���1��U�@�R��� v�����ӯ������ -��Q�<�u�`���`O �O�O���޿��;� &�_�J�oϕπϹϤ� �������%��"�[� F��Fo�ߵ����ߠo ��d�!���W�>�{� b������������ ��A�,�>�w�b��� �������������=��$FNO ����\��
F0�l q  FLAG�>�(RRM_C�HKTYP  r] ��d �] ���OM� _MI�N� 	���� ��  XT SSB_CFG ?\ �����OTP�_DEF_OW � 	��,IR�COM� >�$G�ENOVRD_D�O��<�lTH�R� d�dq_�ENB] qR�AVC_GRP s1@�I X( / %/7//[/B// �/x/�/�/�/�/�/? �/3??C?i?P?�?t? �?�?�?�?�?OOO�AO(OeOLO^O�OoR�OU�F\� ��,�B,�8�?���O�O�O	_|_���  DE_��Hy_�\@@m_B��=�vR/��I�O�SMT�G�SUoo|&oRHOSTC�s1H�I� ���zMSM�l[�bo�	127�.0�`1�o  e�o�o�o#z�o�FXj|�l60s	�anonymou�s������Qao�&�&��o �x��o������ҏ� 3��,�>�a�O�� ��������Ο�U%�7� I��]����f�x��� �����ү����+� i�{�P�b�t������ ������S�(�:� L�^ϭ�oϔϦϸ��� ���=��$�6�H�Z� ����Ϳs�������� ��� �2���V�h�z� ��߰���������
� �k�}ߏߡߣ���� ����������C�* <Nq�_���� ��-�?�Q�c�eJ ��n����� ��/"/E�X/j/ |/�/�/�%'/ ?[0?B?T?f?x?� �?�?�?�?�??E/W/�,O>OPObO�KDaEN�T 1I�K P�!�?�O  �P �O�O�O�O�O#_�OG_ 
_S_._|_�_d_�_�_ �_�_o�_1o�_ogo *o�oNo�oro�o�o�o 	�o-�oQu8 n������� �#��L�q�4���X� ��|�ݏ���ď֏7����[���B�QUICC0��h�z�۟���1ܟ��ʟ+���2�,���{�!ROUTER|�X�j�˯!PCJOG̯���!192.�168.0.10���}GNAME �!�J!ROBO�T�vNS_CFG� 1H�I ��Auto-started�$/FTP�/���/ �?޿#?��&�8�J� �?nπϒϤ�ǿ��[� �����"�4ߵ&���� ������濜������� ���'�9�K�]�o�� �����������/ �/�/G���k��ߏ��� ����������1 T���Py���� �"�4�	H-|�Q cu�VD��� �/�;/M/_/q/ �/����/
/�/> ?%?7?I?[?*/?�? �?�?�/�?l?�?O!O 3OEO�/�/�/�/�?�O  ?�O�O�O__�?A_ S_e_w_�O4_._�_�_ �_�_oVOhOzO�O�_ so�O�o�o�o�o�o�_ '9Kno�o� ����o*o<oNo P5��oY�k�}����� pŏ׏����0����C�U�g�y���_�T_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
 �.�FFF9E3����FRS:D�EFAULT��FANUC W�eb Server�
������q��������������WR�_CONFIG ;O�� ����IDL_CPU_kPC"��B���= �BH#MIN�.�BGNR_I�O��� ���% NP�T_SIM_DO�s}TPMOD�NTOLs �_�PRTY�=!O�LNK 1P�� �'9K]o>�MASTEr ��|���O_CFG�ƟUO����CY�CLE���_A�SG 1Q���
 q2/D/V/h/z/ �/�/�/�/�/�/�/
?�?y"NUM�x��Q�IPCH���£RTRY_C�N"�u���SCRQN������ ���R����?���$J23_DS/P_EN����~�0OBPROC�3ܷ�JOGV�1S�_�@��8�?р';ZO'??0CPO�SREO�KANJI_�Ϡu�A#��3T ���E�O�ECL_LM B2e?�@�EYLOGGINʭ������LA�NGUAGE ,_�=� }Q���LG�2U�����J �x�����PC �� �'0������MC:\RS�CH\00\˝L�N_DISP �V�������TOYC�4Dz\A�S�OGBOOK W+��o���o�o���Xi�o�o�o�o�o�~}	x(y��	�ne�i�ekElG_BUFF 1X�	��}2����Ӣ ������'�T� K�]�����������ɏ ۏ���#�P��Ëq�DCS Zxm =���%|d1h`�ฟʟܟ�g�IO ;1[+ �?'����'�7�I�[�o�� ������ǯٯ���� !�3�G�W�i�{�����б�ÿ׿�El TM  ��d��#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g��yߋߝ߈t�SEVt�0m�TYP΁� ��$�}�AR�S"�(_�s�2FL 31\��0�������������5�T�P<P���DmNGNAM�4�U�f�7UPS`GI�5�A��5s�_LOAD�@G %j%@_MOV�u�����MAXUALRM B7�P8��y���3�0Q]&q��Ca]s�@3�~�� 8@=@^+� طv	���V0+�P�A5d�1r���U�� ����E(i Ty������ �/ /A/,/Q/w/b/ �/~/�/�/�/�/�/? ?)?O?:?s?V?�?�? �?�?�?�?�?O'OO KO.OoOZOlO�O�O�O �O�O�O�O#__G_2_ D_}_`_�_�_�_�_�_ �_�_o
ooUo8oyo do�o�o�o�o�o�o�o��o-��D_LDX�DISA^�� �M�EMO_APX�E� ?��
  �0y�����������ISC 1_�� �O�� ��W�i�����Ə�� ���}��ߏD�/�h� z�a����������� ���@���O�a�5� �����������u�� ׯ<�'�`�r�Y���� ��y�޿�ۿ���8� ��G�Y�-ϒ�}϶ϝ� ����m�����4��X��j�#�_MSTR �`��}�SCD 1as}�R���N��� �����8�#�5�n�Y� ��}���������� ��4��X�C�|�g��� ������������	 B-Rxc��� ����>) bM�q���� �/�(//L/7/p/ [/m/�/�/�/�/�/�/ ?�/"?H?3?l?W?�?�{?�?�?�?n�MKC_FG b���?~��LTARM_�2�cRuB ��3WpTNBpMETsPUOp�2�����NDSP_CMN�TnE@F�E�� 	d���N�2A�O�D��EPOSCF�G��NPSTOL 1�e-�4@�<#�
;Q�1;UK_YW7_Y_ [_m_�_�_�_�_�_�_ o�_oQo3oEo�oio�{o�o�a�ASING_CHK  �M^AqODAQ2CfO��7J�eDEV }	Rz	MC:'|�HSIZEn@�����eTASK %�<z%$123456789 ��u�gTRIG 1g�� l<u%���3`���>svvYPaq���kEM_INF� 1h9G �`)AT&�FV0E0(���)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏP� �t�������]�ί�� ���(�۟�^�� #�5�����k�ܿ� � ��ů6��Z�A�~ϐ� C���g�y�������� 2�i�C�h�ό�G߰� �ߩ��ߙϫ������ ��d�v�)ߚ��߾�y� ��������<�N�� r�%�7�I�[������ 9�&��J[��g��>ONITO�R�@G ?;{  � 	EXEC�1�3�2�3�4��5��p�7�8
�9�3�n�R� R�RRR R(R4R@RL�R2Y2e2q2�}2�2�2�2��2�2�3Y3�e3��aR_GRP_SV 1it���q(�a>�0��Z���h�1�ȇ$���'x~q_DCd~�1P�L_NAME �!<u� �!D�efault P�ersonali�ty (from� FD) �4RR�2k! 1j)TE�X)TH��!�AX d�?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�Ox2-?�O�O�O__@0_B_T_f_x_�b<�O �_�_�_�_�_�_o o�2oDoVoho&xRj" �1o�)&0\�b,� �9��b�a �@D�  �a?�ľc�a?�`�a�aA'�6�ew;�	�l�b	 ��xJp���`�`	p �<w �(p� �.r�� K�K ���K=*�J����J���JV�`�kq`q�P�x��|5p@j�@T;;f�r�f�q�a�crs�I�����p���p�r�p�h}�3��´  ��>��ph��`z���Ζ"�Jm�q�  H�N��ac���dw���  �  �P� Q� �� | � а�m�Əi}	�'� � ��I� �  {����:�È�?È=���(�ts��a	���I  �n @H�i~�ab�Ӌ�b�w��uryN0��  'Ж��q�p@2��@�c���r�q5�C�p}C0C�@ C�����`
�AT1]w@B�V~X�%
nwB0h�A��p��ӊ�p@����aDz ���֏���Я	�pv��( �� -��I��-�=�L�A�a�we_q�`��p �?�ff ���m��� ����Ƽuq@ݿ뺝>1�  P�apv( �`ţ� �=�qst^��?���`x`��5p<
6b<���;܍�<����<� <�&P�ό�AO��c1�|�ƍ�?fff?O��?&��qt@�.��J<?�` ��wi4����dly�e� �g;ߪ�t��p�[ߔ� ߸ߣ����� ����6�wh�F0%�r� !��߷�1ى�����E�� E�O�G+� F�!���/� ��?�e�P���t���lyBL�cB��Enw4� ������+��R��s ����������h�Ô�>���I�mXj����A�y�weC��������ؠ#/*/c/N/wi������v/C�`� CHs/`
=$�p�<!�!���ܼ�'�3A�A��AR1AO��^?�$�?���5p±
=ç�>����3�W�
=�#�]�;e��?�����{�����<��>(�B�u���=B0��?����	R��z�H�F�G����G��H�U`�E���C�+���}I#�I���HD�F���E��RC�j�=�>
I���@H�!H�(� E<YD0 w/O*OONO9OrO]O �O�O�O�O�O�O�O_ �O8_#_\_G_�_�_}_ �_�_�_�_�_�_"oo oXoCo|ogo�o�o�o �o�o�o�o	B- fQ�u���� ���,��P�b�M� ��q�����Ώ���ݏ �(��L�7�p�[��� ���ʟ���ٟ����6�!�Z�E�W���#1(�$1��9�K���<ĥ%����Ư!3�8���!�4Mgs��,�I�B+8�J��a���{�d�d������ȿ���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ��ϰ�������  %��  ��h�Vߌ�z߰�&ڀg�/9�$������� 7����A�S�e�w�  ��������������2 F��$�&Gb��������!C���@����8�����F�� DzN�� F?�P D�������)#B�'9K]�o#?���@@*v
��8�8��u8�.
 v ���!3EW i{����:�� ��ۨ�1���$MSKCFM�AP  ��� ����(.�ONREL  �!9��EXCFENBE'q
#7%^!FNCe/�W$JOGOVLI�ME'dO S"d�K�EYE'�%�R�UN�,�%�S?FSPDTY0g&<P%9#SIGNE/W$�T1MOT�/T!��_CE_GRP� 1p��#\ x��?p��?�?�?�? �?O�?OBO�?fOO [O�OSO�O�O�O�O�O _,_�OP__I_�_=_ �_�_�_�_�_oo�_�:o�TCOM_�CFG 1q	-оvo�o�o
Va_A�RC_b"�p)U?AP_CPL�ot$�NOCHECK {?	+ � x�%7I[m ���������!�.+NO_WAI�T_L 7%S2NT�^ar	+�s�_7ERR_12s	)9�� ,ȍޏ��x����&��dT_M�O��t��, v�*oq�9�PARAuM��u	+��`a�ß'g{�� =?��345678901��,��K�]�9� i�������ɯۯ��&g������C��cU�M_RSPACE�/�|����$OD�RDSP�c#6p(O�FFSET_CAsRT�o��DISƿ���PEN_FIL�E尨!�ai��`OPTION_IO�/���PWORK 5ve7s# ��Vŀؤ��p�4�p�	C ���p��<����RG_DSBL  ��P#��ϸ�RIENTTOD ?�C�� !l��UT_SIM_D�$�"���V��LCT w}�h�i���a[�1�_PEXE�j�RATvШ&p%�� ��2^3j)TE�X)TH�)�X d3������� %�7�I�[�m���� �����������!�3�E���2��u����������������c�< d�ASew��� �����Ǎ�^0�OUa0o(�꘯(����u2�, ���O H �@D�  [?��aG?��cc�D�][�Z�;�	l�s��xJ��������< ���� ��ڐH(���H3k7HSM�5G�22G���Gp
͜�'fc�/-,ڐCR�	>�D!�M#{Z/���3�����4 y H "�c/u/�/0�B_����j�c��t�!�/ �/�"t32����/�6  ��P�%�Q%��%�|T���S62�q?'e	'� �� �2I� �  ��+==��ͳ?�;	�h�	�0�I  �n @�2�.��ODv;��ٟ?&gN�]O  ''�uD@!� C�C�@F#H!�/t�O�O sb
��*�@�@��@�e0@B�QA�0Yv:G �13Uwz$o�V_�/z_e_�_�_	���( �� -�2�1�1ta�Ua�"c���:A-���. ? �?�ff���[o"o�_U�`oX�0A�8���o�j>�1  	Po�V(���eF0�f��Y���L�?�嚫�xb0@<
6�b<߈;܍��<�ê<� <�&�,/a�A�;r�@Ov0P?f7ff?�0?&ip�T�@�.{r�J<?�`�u#	�Bdq t�Yc�a�Mw� Bo��7�"�[�F�� j�������ُ�� ��3����,���(��E�� E��3G+� F��a��ҟ �����,��P�;���B�pAZ�>��B ��6�<OίD���P�� t�=���a�s�����6j��h��7o��>��S��O����όFϑ�A�a�_��C�3Ϙ�/�%?��?�A��������#	Ę�a�P �N||CH����Ŀ������@I��_�'�3A��A�AR1AO��^?�$�?������±
=���>����3�?W
=�#� U���e���B��@���{����<������(�B�u���=B0������	�b��H�F�G����G��H�U�`E���C�+���I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻���������  �9�$�]�H�Z���~� ������������#5  YD}h��� ����
C. gR������ �	/�-//*/c/N/ �/r/�/�/�/�/�/? �/)??M?8?q?\?�? �?�?�?�?�?�?O�? 7O"O[OmOXO�O|O�O �O�O�O�O�O�O3_Q�(������b�y�gUU��W_<i_2�3�8��_�_2�4Mgs�_�_�R�IB+�_�_�a���{�miGo@5okoYo�o}l��P'r	P�nܡݯ�o=_�o0�_�[R?Q`�u���  �p���o��/��S� �z
uүܠ�������ڱ�����������  /�M�w�e�𛟉����l2 F;�$��Gb��t�a�a�`�p�S�C�y��@p�5�G�Y�۠F�� Dz�� F�P D��]����پ��ʯܯ�� ��~�?���@U@�?�K�K�꺡K���
  �|�������Ŀֿ� ����0�B�T�fϽ��V� ���{��1���$PARAM�_MENU ?�3�� � DEFP�ULSEr�	W�AITTMOUT���RCV�� �SHELL_W�RK.$CUR_oSTYL��	��OPT��PTB�4�.�C�R_DECSN���e��ߑ� ������������!�3�\�W�i�{���U�SE_PROG �%��%�����C�CR���e����_HOST !��#!��:���T�`��V��/�X����_�TIME��^�� � ��GDEBU�G\�˴�GINP?_FLMSK����qTfp����PGA e ����)CH��^��TYPE�����������  -?hcu� ������// @/;/M/_/�/�/�/�/ �/�/�/�/??%?7?�`?��WORD ?}	=	RSfu_	PNSU��2JOK�DRTE�y�]TRACEC�TL 1x3��� �` �&�`�`�>�6D/T Qy3�%@�0�D � � #T�2@�8B%�6D&6D'6D(6D)�6D*6D`8B,6D-�6D.6D/6D06D1<6A�c�a8@!U��BR��HI�8BTF�8B6D6D	6DU
6D6D6D6DE6D6D^�8B6DU6D6D6D6DT�8B6D6D6DA6DV�8Bj�8B6DA6DҀ8B�8B!6D"6D5OGOYOkO}O�O*�O�D�D�C�P M �R�O�O�O__/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׈.A�Ev��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p���Er� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������� �*��$PGTR�ACELEN  �)�  ���(��>�_U�P z���2m�u�Y�n�>�_CFG {m�#W�(�~���P���� ��DEFSP/D |���aP���>�IN��TR�L }��(�8���IPE_CON�FI��~m��mњ��Ԛ�>�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�8��1��� ´�����B�9����O��9�s�(�>�T?��
5�������� �=��=#�
 ����P;t_�������� G Dz (�
 H�X~i��� ���/�/D///�h/S/�/��
V7�.10beta1���  A��E�"ӻ�A �(�� ?!G��!>����"����!{���!BQ��!�A\� �!���!2p
����Ț/8?J?\?�n?};� ���/� �/�?}/�?�?OO:O %O7OpO[O�OO�O�O �O�O�O_�O6_!_Z_ E_~_i_�_�_�_�_�_ �_'o2o�_VoAoSo �owo�o�o�o�o�o�o .R=v1�/�#F@ �y�}� �{m��y=��1�'� O�a��?�?�?������ ߏʏ��'��K�6� H���l�����ɟ��� ؟�#��G�2�k�V� ��z��������o� �ίC�.�g�R�d��� �������п	���-� ?�*�cώ���Ϯ� �����B�;�f� x�������DϹ��߶� �������7�"�[�F� X��|��������� ��!�3��W�B�{�f� �������� ����� /S>wbt� �����= OzόϾψ����� �� /.�'/R�d�v� �߁/0�/�/�/�/�/ �/�/#??G?2?k?V? h?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O���O�O�O__ ?_*_c_N_�_r_�_�_ �_�_�_o�_)oTf x�to���/�o />/P/b/t/m o�|����� ��3��W�B�{�f� x�����Տ������ �A�S�>�w�b����O ��џ������+�� O�:�s�^�������ͯ ���ܯ�@oRodo�o `��o�o�o��ƿ�o� ��*<N�Y��}� hϡό��ϰ������� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�c�N�ﲟ��� l��������;�&� _�J���n��������� ��,�>�P�:L�� ���������� (�:�3��0iT� x�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?a?s?��?�?X?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O *\&_8_r����_�_��$PLI�D_KNOW_M�  ��� Q�TSV ���P��?o"o4o�OXo�CoUo�o R�SM_?GRP 1��Z'U0{`�@�`uf
�e�`
�5� �gpk 'Pe] o�������X���SMR�c��m1T�EyQ}? yR�� ��������폯���ӏ �G�!��-������� ����韫���ϟ�C� ��)������������寧���QST�a1W 1��)���P;0� A 4��E 2�D�V�h�������߿ ¿Կ���9��.�o� R�d�vψ��ϬϾ�����2�0� Q�	<3��3�/�A�S߂�4l�~ߐߢ��5 ���������6
��.�@��7Y�k�}���8��������M_AD  )���PARNUM  !�}o+��WSCHE� S�
��pf���S��UPDf��x��_CM�P_�`H�� �'��UER_CHK-���ZE*<�RSr��_�Q_MO�G���_�X�_R/ES_G��!��� D�>1bU� y�����/�	/����+/� k�H/g/l/��Ї/�/ �/�	��/�/�/�X� ?$?)?���D?c?h?�����?�?�?�V �1��U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_�INRr�J�b�Ud�2FMASS?O Z�SGMN>OqCMON�_QUEUE a��U�V P~P X�N$ UhN�FV�@�END�A��IEX1E�O�E��BE�@�O>�COPTIO�G���@PROGRAM7 %�J%�@�?����BTASK_I�G�6^OCFG ኤOz��_�PDATuA�c��[@Ц2=�DoVohozo�j2o �o�o�o�o�o)x;M jINFO[��m��D��� �����1�C�U� g�y���������ӏ����	�dwpt�l �)�QE DIT ��_i��^WERF�LX	C�RGADoJ �tZA���¿�?נʕFA��IOORITY�GW���MPDSPNQ�����U�GD��OTO�E@1�X� (/!AF:@E� c�~Ч!tcpn�>��!ud����!icm���?<��XY_�Q�X�=��Q)� *�1�5��P��]�@�L� ��p��������ʿ� �+�=�$�a�Hυϗ�=*��PORT)QH���P�E��_C?ARTREPPX�>�SKSTA�H�
�SSAV�@�tZ	�2500H86A3���_x�
�'��X�@�swPtS��x�ߧ���URGE�@�B��x	WF��DO�F"[W\��������WRUP_DEL�AY �X���RO_HOTqX	B%��c���R_NORM�ALq^R��v�SE�MI�����9�QS�KIP'��tUr�x 	7�1�1�� X�j�|�?�tU������ ��������$J \n4����� ���4FX |j������ �/0/B//R/x/f/�/�/�/tU�$RCgVTM$��D�� �DCR'������!Bz8aB����C	0>?D���<?�7�l�2:��x�Ŝ����ӷG��:��o?�� <
6b�<߈;܍��>u.�?!<�&�?h?�?�? �@>��?O O2ODOVO hOzO�O�O�O�O�O�? �O�O__@_+_=_v_ Y_�_�_�?�_�_�_o o*o<oNo`oro�o�o �o�_�o�o�o�o�o 8J-n��_�� �����"�4�F� X�j�U������ď�� �ӏ���B�T�� x���������ҟ��� ��,�>�)�b�M��� ���������ïկ� Y�:�L�^�p������� ��ʿܿ� ����6� !�Z�E�~ϐ�{ϴϗ� ����-�� �2�D�V� h�zߌߞ߰������� ��
���.��R�=�v� ��k��������� �*�<�N�`�r����� �����������& J\?���� ����"4F�Xj|��!GN_�ATC 1�	;� AT&F�V0E0�A�TDP/6/9/�2/9�ATA��,AT%G1%B960�_+++�,��H/,�!IO_T?YPE  �%�#�t�REFPO�S1 1�V+ 'x�u/�n�/ j�/
=�/�/�/Q?<? u??�?4?�?X?�?�?^�+2 1�V+�/��?�?\O�?�O�?�!3 1�O*O<OvO�O��O_�OS4 1� �O�O�O_�_t_�_+_S5 1�B_T_f_�_o	oBo�_S6 1��_�_�_5o�o�o|�oUoS7 1�lo�~o�o�oH3l�oS8 1�%_����SMAS�K 1�V/  
8?�M��XNOS/�r�������!MOT�E  n��$��_CFG ����q����"PL_RANG������POWER� �����S�M_DRYPRG %o�%�P��TART ���^�UME_PRO�-�?����$_EXE�C_ENB  <���GSPD��Ր8ݘ��TDB��
�sRM�
�MT_'��T����OBO�T_NAME �o����OB_�ORD_NUM �?�b!H863  ��կ���PC�_TIMEOUT��� x�S232�Ă1�� L�TEACH PENDAN��w���-��Ma�intenanc?e Cons����s�"���KCLC/Cm��

���t��ҿ No U�se-��Ϝ�0�N�PO�򁋁z��.�CH_L��3����q	��s�?MAVAIL����糅��SPAC�E1 2��, j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��� ���ߚ� �2�D��� hߊ�|��`������ ����� �2�D�� h��|���`�������(��y���2���� 0�B���f�����{ ���3) ;M_����@��/� /44 FXj|*/���/��/�/?(??=?5 Q/c/u/�/�/G?�/�/ �?O�?$OEO,OZO6n?�?�?�?�?dO�? �?_,_�OA_b_I_w_7�O�O�O�O�O�_ �O_(oIoo^oofo�o8�_�_�_�_�_ �oo6oEf){�x��G �o�� ���
M� ���*�<�N�`� r�������w���o�収���d.��%� S�e�w����������� Ǐَ���Θ8�+�=� k�}�������ůׯ͟ ����%�'�X�K�]� ��������ӿ�������#�E�W� `� @�������x�����\�e����� ������R�d߂�8� j߬߾߈ߒߤ���� ������0�r���X� ������������8�����
�ύ�_M?ODE  �{��/S ��{|�2ς0�����3�	�S|)CWORK�_AD��:��^+R  �{�`�� �� _INTV�AL���d���R_�OPTION� ���H VAT_�GRP 2��u;p(N�k|��_� ����/0/B/�� h�u/T� }/�/�/�/ �/�/�/?!?�/E?W? i?{?�?�?5?�?�?�? �?�?O/OAOOeOwO �O�O�O�OUO�O�O_ _�O=_O_a_s_5_�_ �_�_�_�_�_�_o'o 9o�_Iooo�o�oUo�o �o�o�o�o�o5G Yk-���u� ����1�C��g� y���M�����ӏ叧� 	��-�?�Q�c����� ����������ǟ��;�M�_����$SCAN_TIM���_%}�R ��(�#((�<0�4d d 
!D�ʣ���u�/�����U��25���@��d5�P�g��]	 ���������dd�x��  P����; ��  8� ҿx�!���D��$� M�_�qσϕϧϹ���������ƿv���F�X��/� ;G�ob��pm���t�_Di�Q̡  � l �|�̡ĥ������� !�3�E�W�i�{��� ������������/� A�S�e�]�Ӈ����� ��������); M_q����� ��r���j�T fx������ �//,/>/P/b/t/��/�/�/�/�/�%�/  0��6��!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O*�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo�O�OJ�o�o �o�o�o�o�o 2 DVhz��������
�7?   ;�>�P�b�t������� ��Ǐُ����!�3� E�W�i�{�������ß �ş3�ܟ�� &�8�J�\�n�������������ɯ�����,� �+�	�1234567�8�� 	� =5���f�x�������������
��.� @�R�d�vψϚ�៾� ��������*�<�N� `�r߄߳Ϩߺ����� ����&�8�J�\�n� �ߒ����������� �"�4�F�u�j�|��� ������������ 0_�Tfx��� ����I> Pbt����� ��!/(/:/L/^/ p/�/�/�/�/�/�/�2�/?�#/9?K?�]?�iCz  B}p˚   ��h�2��*�$SCR�_GRP 1�(��U8(�\x�d�@} � ��'�	 �3�1�2�4(1*�&��I3�F1OOXO}m��D�@�0ʛ�)���HUK�LM�-10iA 89�0?�90;��F;�M61C D�:�CTP��1
\&V�1 	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^�o OUO>oPo#G�/����o'o�o�o�o�oB��0�rtAA�0*  @�Bu&"Xw?��ju�bH0{�UzAF@ F�`�r��o���� �+��O�:�s��mBq�rr����������B� ͏b����7�"�[�F� X���|�����ٟğ�� �N���AO�0�B�CU�
L���E�jqBq>m3󵔯$G@�@pϯ7 B���G�I�
E�0EL_DEFAULT  �T���E���MIPOWERFL  
E*���7�WFDO� �*��1ERVENT? 1���`(��� L!DUM�_EIP��>��j�!AF_INEx�¿C�!FT�������!o:� ���a�!RP?C_MAINb�D�q�Pϭ�t�VIS}��Cɻ����!TP&��PU�ϫ�d��E��!
PMON_POROXYF߮�e4ߐ���_ߧ�f����!�RDM_SRV��߫�g��)�!R��Iﰴh�u�!
�v�M�ߨ�id���!RLSYNC���>�8���!R3OS��4��4��Y� (�}���J�\������� ������7��[" 4F�j|�����!�Eio�I�CE_KL ?%�� (%SVCPRG1n>����3��3���4�//�5./3/�6V/[/�7~/�/��D$�/�9�/�+�@� �/��#?��K?� �s?� /�?�H/�? �p/�?��/O��/ ;O��/cO�?�O� 9?�O�a?�O��?_ ��?+_��?S_�O {_�)O�_�QO�_� yO�_��Os��� �>o�o}1�o�o�o�o �o�o�o;M8 q\������ ���7�"�[�F�� j�������ُď��� !��E�0�W�{�f��� ��ß���ҟ��� A�,�e�P���t�����࿯�ί�y_DE�V ���MC:��_.!�OUT��2�~�REC 1�`e��j� �� 	 �����ȿ೿�׿��!�
 ��PJ�%6 (�޷&�!�a�}���u,��0�  Z�+ 3��3��Ge3�c���V��˒��� � ��$��H�6�l�~�`� �ߐ��ߴ������� � ��V�D�z�h��� ����������
�� R�@�v���j������� ������*N< ^�r����� �&J8Z� b������� "/4//X/F/|/j/�/ �/�/�/��2��/�/�/ ?:?(?^?L?�?�?v? �?�?�?�?�?�? O6O OFOlOZO�O~O�O�O �O�O�O_�O2_ _B_ h_V_�_n_�_�_�_�_ �_
o�_.o@o"odoRo tovo�o�o�o�o�o�o <*`Np� x������� 8�J�,�n�\������� ��Ə�Ώ�����F��4�j�X���`�p�V [1�}� P��m���ܺ)I�� !<��TYPE\���HELL_CFG� �.�F��� � 	�����RSR������ӯ����� ��?�*�<�u�`��������������/  ��!%�3�PE��Q�\���M�Lo�p�����2���d]�K�:�HK 1�H� u����� ��A�<�N�`߉߄� �ߨ������������&�8��=�OMM ��H���9�FTOV_ENB&��!1��OW_REG_U�I��8�IMWAI�T��a���OUTr������TIM��w���VAL��>��_UNIT��K��1�MON_ALI�AS ?ew� ( he�������� ����і��);M ��q����d� �%�I[m �<����� �!/3/E/W//{/�/ �/�/�/n/�/�/?? /?�/S?e?w?�?�?F? �?�?�?�?�?O+O=O OOaOO�O�O�O�O�O xO�O__'_9_�O]_ o_�_�_>_�_�_�_�_ �_�_#o5oGoYokoo �o�o�o�o�o�o�o 1C�ogy�� H����	��-� ?�Q�c�u� ������� ϏᏌ���)�;�� L�q�������R�˟ݟ �����7�I�[�m� �*�����ǯٯ믖� �!�3�E��i�{��� ����\�տ����� ȿA�S�e�wω�4ϭ� �����ώ����+�=� O���s߅ߗߩ߻�f� ������'���K�]� o���>�������� ���#�5�G�Y��}����������o��$S�MON_DEFP�RO ������ �*SYSTEM�*  d=��R�ECALL ?}��� ( �}/�xcopy fr�:\*.* vi�rt:\tmpb�ack7=>in�spiron:11828 Ybt\�� }0.a6�HZ_��
�xyzrate 61 ���n���.M3304 HZ��/��3/s:orde�rfil.dat�<�a/s/�/�/� */mdb:9�Y/�/�/?�	..A� �/n?�?�?�-�G? Y2_?�?OO'/9/�/ ]?nO�O�O�/�?�/[O �O�O_#?5?�?Y?j_ |_�_�?�?D_�?�_�_ oO1O�OUOfoxo�o �O�OJo�O�o�o�o -_�_Q_bt���_ <�_����)����p������N6368�Y����� !o3o�o��a�s����� �oE���Y�����! 3F�ݟn������ 6�H�ŀ^����&� 8���ܟm�������� ȟZ�����"�4�ǯ X�i�{ύϠ���C�֯ ������0�����e��w߉ߜ���U 2112ǏY������!�3� ������n���߷�400G�Y������ !�3�����a�s����� ��E���Y�����!� 3�F�����n���� 6H��^�&� 8�����m����� ��Z��/"4� Xi/{/�/��C/� �/�/?0BTe? w?�?��I?��?�?�OO�$SNPX�_ASG 1�����9A�� P 0 '�%R[1]@g1.1O9?�$3%dO�OsO�O�O�O�O �O�O __D_'_9_z_ ]_�_�_�_�_�_�_
o �_o@o#odoGoYo�o }o�o�o�o�o�o�o* 4`C�gy� ������	�J� -�T���c�������ڏ �����4��)�j� M�t�����ğ������ ݟ�0��T�7�I��� m��������ǯٯ� ��$�P�3�t�W�i��� �����ÿ����:� �D�p�Sϔ�wω��� ���� ���$���Z� =�dߐ�sߴߗߩ��� ���� ��D�'�9�z� ]���������
� ���@�#�d�G�Y��� }�������������* 4`C�gy� �����	J -T�c���� ��/�4//)/j/ M/t/�/�/�/�/�/�/��/?0?4,DPAR�AM �9E�CA �	��:P�4�0$HOFT�_KB_CFG � q3?E�4PIN_SIM  9K��6�?�?�?�0,@R�VQSTP_DS�B�>�21On8J0S�R ��;� &� MULTIR�OBOTTASK�=Oq3�6TOP�_ON_ERR � �F�8�APTN� �5�@�A�BRING_�PRM�O J0V�DT_GRP 1y�Y9�@  	�7 n8_(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 Dkhz���� ���
�1�.�@�R� d�v���������Џ�� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\������� ����ȯگ����"� I�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� tߛߘߪ߼������� ��(�:�a�^�p�� ���������� �'� $�6�H�Z�l�~��������������3VPRG_COUNT�6���A�5ENB��OM=�4J_U�PD 1��;8  
q2��� ��� )$6H ql~����� /�/ /I/D/V/h/ �/�/�/�/�/�/�/�/ !??.?@?i?d?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_�_�_Y?SDEBUG" � ��Pdk	�PSP_�PASS"B?~�[LOG ��+m�P�X�_�  �g�Q
M�C:\d�_b_M�PCm��o�o��Qa�o �vfSAV �m:dUb�U�\gSV�\TE�M_TIME 1]�� (�`#�S�!�o	T1SV�GUNS} #'�k�spASK_OPTION" �g�ospBCCFGg ��| �b�{�}`����a &��#�\�G���k��� ��ȏ������"�� F�1�j�U���y���ğ ���ӟ���0��T�f��UR���S���Ư A������ ��D��n d��t9�l��������� ڿȿ�����"�X� F�|�jϠώ��ϲ��� ������B�0�f�T� v�xߊ��ߦؑ����� ��(��L�:�\�� p�����������  �6�$�F�H�Z���~� ������������2  VDzh��� ������4F dv����� �//*/�N/</r/ `/�/�/�/�/�/�/�/ ??8?&?\?J?l?�? �?�?�?�?�?�?�?O O"OXOFO|O2�O�O �O�O�OfO_�O_B_ 0_f_x_�_X_�_�_�_ �_�_�_oooPo>o tobo�o�o�o�o�o�o �o:(^Ln p�����O�� $�6�H��l�Z�|��� ��Ə؏ꏸ����2�  �V�D�f�h�z����� ԟ����
�,�R� @�v�d���������ί Я���<��T�f� ������&�̿��ܿ� �&�8�J��n�\ϒ� �϶Ϥ���������� 4�"�X�F�|�jߌ߲� ������������.� 0�B�x�f��R����� �������,��<�b� P�������x������� ��&(:p^ �������  6$ZH~l� �������/&/ D/V/h/��/z/�/�/�/�/�&0�$TB�CSG_GRP �2��%��  �1 
 ?�  /?A?+? e?O?�?s?�?�?�?�?��;23�<d�, �$A?1	 �HC���6>���@E�5CL  B�'2^OjH4J��B\)LFY  3A�jO�MB��?�I#Bl�O�O�@�JG_>�@�  D	�15_ __$YC-P{_F_`_j\��_�]@0�>�X �Uo�_�_6oSoo0o�~o�o�k�h�0	�V3.00'2	�m61c�c	�*�`�d2�o�e>�dJC0(�a�i ,p��m-  �0�����omvu1JCFoG ��% 1Y #0vz��rBr�|�|����z � �%��I�4�m�X� ��|��������֏� ��3��W�B�g���x� ����՟������� �S�>�w�b�����'2 A ��ʯܯ������ E�0�i�T���x���ÿ տ翢����/��?� e�1�/���/�ϜϮ� �������,��P�>� `߆�tߪߘ��߼��� �����L�:�p�^� ������������  �6�H�>/`�r���� ������������  0Vhz8��� ���
.�R @vd����� ��//</*/L/r/ `/�/�/�/�/�/�/�/ �/?8?&?\?J?�?n? �?�?�?�?���?OO �?FO4OVOXOjO�O�O �O�O�O�O__�OB_ 0_f_T_v_�_�_�_z_ �_�_�_oo>o,obo Poroto�o�o�o�o�o �o(8^L� p������� $��H�6�l�~�(O�� ��f�d��؏���2�  �B�D�V�������n� ���ԟ
���.�@�R� d����v�������� Я���*��N�<�^� `�r�����̿���޿ ��$�J�8�n�\ϒ� �϶Ϥ�������ߊ� (�:�L���|�jߌ߲� �����������0�B� T��x�f������ �������,��P�>� t�b������������� ��:(JL^ ������ � 6$ZH~l� �^���dߚ // D/2/h/V/x/�/�/�/ �/�/�/�/?
?@?.? d?v?�?�?T?�?�?�? �?�?OO<O*O`ONO �OrO�O�O�O�O�O_ �O&__6_8_J_�_n_ �_�_�_�_�_�_�_"o oFo��po�o,oZo �o�o�o�o�o0 Tfx�H��� ����,�>��b� P���t���������Ώ ��(��L�:�p�^� ������ʟ���ܟ�  �"�$�6�l�Z���~� ����دꯔo��&� ЯV�D�z�h������� Կ¿��
��.��R��@�v�dϚτ�  ���� ��������$TBJOP_�GRP 2ǌ���  �?�������������x�JBЌ��9� �< �X�ƞ�� @���	� �C�� t�b�  C����>ǌ�͘Րդ�>���йѳ33=��CLj�fff?>��?�ffBG���Ќ�����t�ц�>;�(�\)�ߖ��E噙�;��h{CYj��  @h�~�B�  A�����f��C�  D�hъ�1��O��4�N����
:�/��Bl^��j�i��l�l����Aə�3A�"��D���Ǌ=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������<$�6�>B�\��T����Q�tsx�@g33@���C����y�1����>��Dh����������O<{�h�@i�  ��t��	� ��K&�j� n|���p�/��/:/k/�ԇ����!��	V3.0}0J�m61cIԃ*� IԿ��/�'� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�I�!CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;��;Q�UT,8�4` *���?�2���3\�X/�O��ESTPAR�S  ��	���H�R@ABLE 1%����0��
H�7Q 8��9
G
H
H�����
G	
H

H�
HYE��
H
H:
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_�^:BS _� �JGoYo ko}o�o�o�o�o�o�o �o1CUgy ����`#oRL�y�_ �_�_�_�O�O�O�O�O�X:B�rNUM  ����P���� V@P:B_CF�G ˭�Z�h�@���IMEBF_T�T%AU��2@�VE�RS�q��R {1���
 (�/����b� ����J� \���j�|���ǟ��ȟ ֟�����0�B�T�@��x�������2�_����@�
��MI_�CHAN�� � >��DBGLV����������ETHE�RAD ?��
O�������h������ROUT�!���!������SN�MASKD��U�255.���#������OOLOFS_�DI%@�u.�OR�QCTRL � ����}ϛ3rϧϹ��� ������%�7�I�[��:���h�z߯�APE?_DETAI"�G��PON_SVOF�F=���P_MON� �֍�2��S�TRTCHK ��^�����VTCOMPAT��O������FPROG �%^�%MULTIROBOTTݱx���9�PLAY&H���_INST_M�ް ������US8�q��LCK���QUICKME��=���SCREZ�}G�tps� @���u�z����_���@@n�.�SR_GR�P 1�^� �O����
��@+O=sa�� ��
m������ L/C1gU� y�����	/��-//Q/?/a/�/	1234567�0h�/�/@Xt�1����
 �}ipn�l/� gen.htm�? ?2?D?V?�`Panel� setupZ<}�P�?�?�?�?�?�? �??,O>OPObOtO �O�?�O!O�O�O�O_ _(_�O�O^_p_�_�_ �_�_/_]_S_ oo$o 6oHoZo�_~o�_�o�o �o�o�o�oso�o2D Vhz�1'� ��
��.��R�� v���������ЏG����UALRM��G ?9� �1�#� 5�f�Y���}������� џן���,��P���SEV  �����ECFG C��롽�A���   BȽ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �(�� ��3�/SOFTPAR�T/GENLIN�K?curren�t=editpa7ge,��,1���8!�3��� �����menu��962 �߆����K�]�o�36u�
��.�@��� W�i�{���������R� ����/A��e w����N�� +=O�s� �������f�� f//'/9/K/]/` �/�/�/�/�/�/j/�/ ?#?5?G?Y?�/�/�? �?�?�?�?�?x?OO 1OCOUOgO�?�O�O�O �O�O�OtO�O_-_?_ Q_c_u__�_�_�_�_ �_�_��)o;oMo_o qo�o�_�o�o�o�o�o �o%7I[m � ������ �3�E�W�i�{���� ��ÏՏ������� A�S�e�w�����*��� џ�����ooO� a�s���������ͯ߯ ���'���K�]�o� ��������F�ۿ��� �#�5�ĿY�k�}Ϗ� �ϳ�B��������� 1�C���g�yߋߝ߯� ��P�����	��-�?� *�<�u������� ������)�;�M��� �������������l� %7I[�� �����hz !3EWi��� ����v////�A/S/e/P���$U�I_PANEDA�TA 1������!  	�}w/�/�/�/�/?? )?>?� �/i?{?�?�?�?�?*? �?�?OOOAO(OeO LO�O�O�O�O�O�O�O��O_&Y� b� >RQ?V_h_z_�_�_�_ _�_G?�_
oo.o@o Rodo�_�ooo�o�o�o �o�o�o*<#`@G��}�-\�v �#�_��!�3�E�W� �{��_����ÏՏ� ��`��/��S�:�w� ��p�����џ����� �+��O�a����� ����ͯ߯�D���� 9�K�]�o�������� ɿ���Կ�#�
�G� .�k�}�dϡψ����� ����n���1�C�U�g� yߋ��ϯ���4����� 	��-�?��c�J�� ������������ ��;�M�4�q�X���� �������%7 ��[������ �@��3W iP�t���� �/�//A/����w/ �/�/�/�/�/$/�/h ?+?=?O?a?s?�?�/ �?�?�?�?�?O�?'O OKO]ODO�OhO�O�O �O�ON/`/_#_5_G_ Y_k_�O�_�_?�_�_ �_�_oo�_Co*ogo yo`o�o�o�o�o�o�o �o-Q8u�O�O}��������)�>��U-�j� |�������ď+��Ϗ ���B�)�f�M��� �����������ݟ��&�S�K�$UI_�PANELINK� 1�U�  �  ���}1234567890s����� ����ͯդ�Rq���� !�3�E�W��{����� ��ÿտm�m�&����Qo�  �0�B� T�f�x��v�&ϲ��� ������ߤ�0�B�T� f�xߊ�"ߘ������� ���߲�>�P�b�t� ���0��������� ���$�L�^�p����� ,�>������� $�0,&�[gI� m������ �>P3t�i� �Ϻ� -n��'/ 9/K/]/o/�/t�/�/ �/�/�/�/?�/)?;? M?_?q?�?�UQ�= �2"��?�?�?OO%O 7O��OOaOsO�O�O�O �OJO�O�O__'_9_ �O]_o_�_�_�_�_F_ �_�_�_o#o5oGo�_ ko}o�o�o�o�oTo�o �o1C�ogy �����B�	� �-��Q�c�F����� |�������֏�)� �M���=�?��?/ ȟڟ����"�?F� X�j�|�����/�į֯ �����0��?�?�? x���������ҿY�� ��,�>�P�b��� �Ϫϼ�����o��� (�:�L�^��ςߔߦ� ��������}��$�6� H�Z�l��ߐ����� ����y�� �2�D�V� h�z����-������� ��
��.RdG ��}����c� ��<��`r�� ������//&/ 8/J/�n/�/�/�/�/ �/7�I�[�	�"?4?F? X?j?|?��?�?�?�? �?�?�?O0OBOTOfO xO�OO�O�O�O�O�O _�O,_>_P_b_t_�_ _�_�_�_�_�_oo �_:oLo^opo�o�o#o �o�o�o�o ��6 H�l~a��� �����2��V� h�K�������1� U
��.�@�R�d�W/ ��������П����� �*�<�N�`�r��/�/ ?��̯ޯ���&� ��J�\�n�������3� ȿڿ����"ϱ�F� X�j�|ώϠϲ�A��� ������0߿�T�f� xߊߜ߮�=������� ��,�>���b�t�� ����+���� ��:�L�/�p���e��� �������� ��6����ۏ��$U�I_QUICKM�EN  ����}��RE�STORE 1����  �
�8m3\n���G ����/�4/F/ X/j/|/'�/�/�// �/�/??0?�/T?f? x?�?�?�?Q?�?�?�? OO�/'O9OKO�?�O �O�O�O�OqO�O__ (_:_�O^_p_�_�_�_ QO[_�_�_I_�_$o6o HoZoloo�o�o�o�o �o{o�o 2D�_ Qcu�o���� ���.�@�R�d�v���������Џ⏜S�CRE� ?��u1sc� �u2�3�4�5*�6�7�8���USER����TL���ks'���4��U5��6��7��8���� NDO_CFG� ڱ  �  �� PDATE �h��No�ne�SEUFR�AME  �ϖ��RTOL_A�BRT����EN�B(��GRP 1���	�Cz  A�~�|�%|�������į֦��X�� �UH�X�7�MSK � K�S�7�N��%uT�%�����V�ISCAND_M;AXI�I�3����FAIL_IMG�I�z �% #S���IMREGNUMI�9
���SIZI�� ��ϔ,�ONOTMOU'�K�Ε��&����a���a��s��FR:\�� � MC:\(��\LOGh�B@Ԕ !{��Ϡ������z MCyV����UD1 ֓EX	�z ��POO64_�Q���n6��PO!�L!I�Oڞ�e�V�N��f@`�I�� =�	_�SZVmޘ���`�WAImߠ�S?TAT �k�% !@��4�F�T�$#�x���� �2DWP  ?��P G��=��͎����_JMPERR �1ޱ
  �p2�345678901���	�:�-�?� ]�c������������������$�MLOWp�ޘ�����_TI/��˘'��MPHA�SE  k�ԓ|� ��SHIFT%�k1 Ǚ��< z��_���� F/|Se�� �����0/// ?/x/O/a/�/�/�/�/�/����k�	V�SFT1\�	V:��M+3 �5�Ք� p����A�  �B8[0[0�Πp�g3a1Y2�_3Y�7ME��K�͗	6e���W&%��M����b��	��$��TDINEND3�4��4AOH�+�G1�OS2O�IV I���]LRELEvI��4.�@�~�1_ACTIV�IxT��B��A �m�0�/_��BRDBГO�Z�YBOX �Xǝf_\��b�2�T�I190.�0.�P83p\N�V254p^�Ԓ�	 �S�_�[b���robot�84q_   �p�9o\�pc �PZoMh�]Hm�_Jk@1��o�ZABCd��k�,���P\�Xo}�o 0);M�q� �������>��aZ�b��_V