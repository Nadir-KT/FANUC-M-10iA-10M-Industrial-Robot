��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�O�AUTOBA�CKU0 ?$ENAB��!oEVIC�TI� � D� DX�!2ST� ?0B�#$�INTERVAL�!2DISP_UNsIT!20_DOn6�ERR�9FR_F�!2IN,GRE5S�!0Q_;3!4�C_WA�471�:O�FF_ N�3DELHLOGn25A�a2?i1@N?�� -M��A�W+0�$Y $D�B� 6COMW!2MO� "0G_A.o	 \rVE�1�$F��A{$�O��D�B�CTMP�1_F�E2�G1_��3�B�2GXD��#
 d $�CARD_EXI�ST4$FSS�B_TYPuAH�KBD_S�B�1A�GN Gn $�SLOT_NUM�JQPREV,DB�U� g1G ;1_ED�IT1 � *1G=� S�0�%$EP�$�OP�AEToE_OKRUS�oP_CRQ$;4x�V� 0LACIw�1�RAPk �1x@M}E@$D�V��Q�Pv�A{oQLv� OUzR ,mAЧ0�!� B� LM�_O�^eR�"CAsM_;1 xr~$ATTR4�NP� ANN�@5I�MG_HEIGH|Q�cWIDTH4�VT� �UU0F_�ASPECQ$�M�0EXP��@A�X�f�CFT ?X $GR� � �S�!�@B@NFL�I�`t� UIREx 3dTuGITCHCj�`N� S�d_L�`2�C�"�`EDlpE
� J�4S�0� �zsa�!ip;G0 �� 
$WARNM��0f�!,P� �s�pN{ST� CORN�"�a1FLTR�uTRkAT� T�p H0ACCa1���{��ORI
`"S={R�T0_S�B�qHG�,I1 [ Thp�"3I9�TY�D(,P*2 �`w@� X�!R*HD�cJ* TC��2��3��4��U5��6��7��8���94�qO�$ <� $6xK3 1w`�O_M�@�C t� � E#6NGP�ABA� �c��ZQ ���`���@nr���� ��P�0����x�p�PzPb26��4��"J�_R��B�C�J��3�JV P��tBS��}Aw��"v�tP_*0OFSzRw @� RO_K8̨��aIT�3��NO�M_�0�1ĥ3vFCPT �� �$���AxP��K}EX �� �0g0I01��p��
$TFa��C$M�D3��TO�3�0U�� �� �H�w2�C1|�EΡg0@wE{vF�vF���hp@�a2 
P$A`�PU�3N)#�dR*�AX�!sDEwTAI�3BUFV8��p@1 |�p۶��pPIdT� PP�[�MZ�Mg�Ͱj�F>[�SIMQSI�"�0��A.������lw Tp|zM��P�B^�FACTrbHPEW7�P1Ӡ��v���MCd� �$�*1JB�p<�*1DE�CHښ�H��(�c�� � +PNS_wEMP��$GP����,P_��3�p�@Pܤ��TC��|r��0 �s��b�0�� �B���!�
���JR� ��SE�GFR��Iv �aRʟTkpN&S,�PV�F���� &k�Bv�u�cu��aEЀ� !2��+�MQ��E�SCIZ�3����T���P�����aRSINF�����kq��������LX�����F�gCRCMu�3CClp G��p���O}���b�1@�������2�V�DxIC��C���r����P���{� EV �zF*_��F�pNB0��?������A�! �r�Rx����V� lp�2��aR�t�,�g���RTx @#�5�5"2��uAR��:�`CX�$LG�p���B�1 `s�P�t�aA�0{�У+0R���t�ME�`!BupCrRA 3tAZ�л�pc�OT�FC�b�`�`�FNp���1��ADI+�a%��b�{�@�p$�pSp�c�`S�P���a,QMP6�`Y$�3��M'�pU��a�U  $>�TITO1�S�S�!��$��"0�DBPXWO���!��$SK@��2�P� �"�"v@�PR8� 
� 8���# >�q1�$��$��+�LB9$?(�V�%@?�R4C&_?R4ENE��'~?(�� �RE�pY2(H ��OS��#$L�3$$3R��;3��MVOk_D@!V�ROScrr�w�S���C�RIGGER2FP�A�S��7�ETUR�N0B�cMR_��T�Uː[��0EWM%���GN>`��R#LA���Eݡ�P�O&$P�t�'�@D4a��C�DϣV�DXQ���4�1��MVGO_oAWAYRMO#��aw!�DCS�_)  `IS#� �� �s3S�AQ汯 4Rx�ZSW��AQ�p�@1UW��cTNTV)�5RV
a���� |c�éWƃ��JB��<x0��SAFEۥ�V�_SV�bEXCL�UU�;��ONLĆ�cYg�~az�OT<�a{�HI_V? ��xR, M�_ *�0�� ��_z�2� �CdSGO  + �rƐm@�A�c~b����w@��V�i�b�fAN�NUNx0�$�dIDY�UABc�@Sp�i��a+ �j�f��ΰAPI:x2,��$F�b�$�ѐOT�@A ?$DUMMY��Ft���Ft±� 6U-o ` !�HE��|s��~bc�B@ SU�FFI��4PCUA�Gs5Cw6Cq��DMSWU. =8!�KEYI��5�TM�1�s�qoA�vI�Nޱw��", / �D��HOST�P!4���<���<�°<��p<�EM'���Z�� �SBL� UL��0  �	�����DT�01 �� $��9USAMPLо�/���決��$ I@갯 $SUBӄ��w0QS�����#��SAV������c�S< 9�`�fP$��0E!� YN_Bn�#2 0�`DI�db�pO|�m��#$F��R_IC� �E�NC2_Sd3C  ��< 3�9���@� cgp����4�"Ȼ�2�A��ޖ5����`ǻ�@Q@K�&D-!�a�AVERp�q����DSP
���PC_�q��"�|��ܣ�VALU3�HiE�(�M�IP)î��OPPm �T!H�*��S" T�/�Fb�;�d����d �D�qЗ16 }H(rLL_DUǀ��a�@��k���֠OaT�"U�/����R_NOAUTO70�$}�x�~�R@s��|�C� ��YC� 2w�L�� 8H *��L� ���Բ@sv��` � �� ÿ���Xq��cq����q���q��7��8J��9��0���1�U1 �1-�1:�1G�U1T�1a�1n�2|ʩ2��2 �2-�2�:�2G�2T�2a�2*n�3|�3�3� �U3-�3:�3G�3T�3a�3n�4|�ia����9 <���z�ΓKI����H硵Ba�FEq@{@: ,<��&a? P_P�?h`$>�����E@�@���qQQ��;fp�$TP�$V�ARI����,�UP�2Q`< W�߃TD ��g���`������ ���BAC�"= T2����$)�,+r³�p IFI��p�� �q M�P"<��F�l@``>t ;h��6����ST� ���T��M ����0	��i���F����������kRt ����FOR�CEUP�b܂FL+US
pH(N��� ���6bD_CM�@E �7N� (�v�P��REM� Fa���@j���
K�	N���EFF/���@3IN�QOV���OVA�	TROV� DT)��DTMX:e �P:/���Pq�vXpCL�N _�p��@ ��	_�|��_T: �|�J&PA�QDI����1��0�Y0RQDm�_+qH���M���CL�d#�RIV�{�ϓN"EAR/�I�O�PCP��B�R��CM�@N 1b =3GCLF��!�DY�(��a�#5T��DG���� �%	?(�FSS� )��? P(q1�1��`_1"811�E�C13D;5D6�GSRA���@�����PW�ON2EBUG�S�2�C`g�ϐ_E A ���?����TERMr�5B�5 �ORIw�0C�5���SM_�-`���0D�5&��TA�9EIUP>��F� -Qϒ�A�P�3�@B$S�EGGJ� EL�UU�SEPNFI���pBx��1@��4>DC$sUF�P��$����Q�@C���G�0T������SNSTj�P�ATۡg��APTH	J�A�E*�Z%qB\`@F�{E��F�q�pARxP<Y�aSHFT͢qA|�AX_SHOR$��>��6 @$GqPE���OVR���aZP�I@P@$U?r *aAGYLO���j�I�"���Aؠ��ؠERV ��Qi�[Y)��G�@R���i�e��i�R�!P�uASYM���uqA#WJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P���WkOR�@M��k0�SMT��G��GR��3�aPA�@��p|5�'�H � j��A�TOCjA7pP<]Pp$OPd�O�P�C�%�p�O!���RE.pR�C�AOX�?��Be5pR�E�ruIx'QG�e$PW�R) IMdu�RR_p$s��5��B Iz2�H8�=�_ADDR~H�H_LENG�BP�q�q:�x�R��So�mJ.�SS��SK������� ��-�SEh*���rSN�MN1K	�j�5�@r�֣OL��\�WpW�Q�>pACRO�p���@�H ����Q� ��OSUPW3�b_>�I��!q�a1�������� |��������-���X:���iIOX2S=��D�e��]���L� $��p�!_OFyF[r_�PRM_炽�rTTP_�H��M (�pOBJر"��G�$H�LE��C��ٰN � �9�*�AB_�T���
�S�`�S��LV漣KRW"duHIT�COU?BGi�LO�q����d� �Fpk�GpSS� ����HWh�wA��O.���`INCPUX2VISIO��!��¢�.�á<�á-� �IwOLN)�P 87�yR'�[p$SL�b�d PUT_��	$dp�Pz �� �F_AS2Q/��$LD���D�aQT U�0]P�A������P�HYG灱Z�DS9�4�UO� 3R ` F���H�Yq�Yx�ɱvpP�Sdp���x��,ٶ�1UJ��S����;NE�WJOG�G �'DIS��&�KĠ��&3T |��AV��`�_�CTR!S^�FL�AGf2AP�LG�dU �n�:��3?LG_SIZ��`�ň��=���FD��I����Z �ǳ��0�� ��@s��-ֈ�-�=�-����-��0-�ISCHy_��Dq �LN?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHrܵ�I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn���_BWUFF1XY��PT�$�� �v���f���װA�rYY���P �����pOS1*�2�3�L�>0Z �  ��apiE�*��IDX�d	P�RhrO�+��A&+ST��R��Yz�<!� Y$EK&C K+���Z&m&�5�0[ L��o�0�� ]PL�6pwq�t^����w���7�_ \ ��`��瀰�7��#�0C��] ��CLD�P��;eTRQLI��jd.�094FLG z�0r1R3�DM�R7Ɩ�LDR5<4R5ORG.���e2(`���V�8�.��T<�3�d^ A�q�<4��-4R5S�`�T00m��0DFRCLMC!D�?�?3I�@��MIC��d_ Yd���RQm�q��DSTB	�  ؏Fg�HAX;b |�H�LEXCESZr��rBMup�a`�@�B;d�!rB`��`a��F_A�J��$[�Ot�H0K�db \���ӂS�$MB��LI�Б}SREQUIR��R>q�\Á�XDEB�U��oAL� MP�c@�ba��P؃ӂ!BoA#ND���`�`d�҆��c�cDC1��IN@�����`@�(h?Nz��@q��o��UPST�8� e�rLOCf�RI�p�EX�f�A�p��AoAODA�QP�f X��ON��[rMF�����f)@�"I��%�e��T���FX�@IGG� g �q��"E�0�h�#���$R�a%;#�7y��Gx��VvCPi�D'ATAw�pE:�y���RFЭ�NVh t_ $MD�qIёA)�v+�tń�tH�`��P�u�|��sANSAW}��t�?�uD��)�b�	@Ði �@CU��V�T0�ewRR2�j Dɐ��Qނ�Bd$CALII�@F�G�s�2⠧RIN��v�<�I'NTE���kE����,��b����_Nl@��ڂ��kDׄRm�7DIViFDH�@ـ:n�$V��'cv!$��$Z������~�[��o�H �$BEL�Tb��!ACCEL�+��ҡ��IRC��t����T/!���$PS�@#2L� q�Ɣ83������� ��PATH��������3̒Vp�A_�Q�.��4�B�Cᐈ�_M=Gh�$DDQ���G�$FWh��p���m�����b�DE��P�PABNԗROTSPEED����00�J�Я8��@����$USE_��P���s�SY��c�A �kqYNu@Ag��OsFF�q�MOUN�3NGg�K�OL�H�INC*��a��q��Bxj�L@�BENCS���q�Bđ���D��IN�#"I̒��4�\BݠV�EO�w�Ͳ23_UyPE�߳LOWLA���00����D��@�BwP��� �1RCʀ�ƶMOSIV�JRM�O���@GPERC7H  �OV�� ^��i�<!�ZD<!�c@��d@�P��V1�#P͑��L���EW�ĆĸUP������T�RKr�"AYLOA'a�� Q-�(�<�1�8�`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H�����b�DUM2(�S_�BCKLSH_C (���>�=�q�#�U��������2�t�]ACLA�LvŲ�1n�P�C�HK00'%SD�RT�Y4�k��y�1�q_�6#2�_UM$Pj�C�w�_�SCL��ƠLMT_J1_LO�"�@���q��E������๕�幘SPC`��7������PCo�B��H� �PU�m�C/@��"XT_�c�CN_b��N��e���SFu���V�&#����9�(�d��=�C�u�SH6# ��c����1�Ѩ�o�0�0͑
��_�PAt�h�_Ps�W�_10��4֠R�01D�VG�J� L��@J�OGW���ToORQU��ON*ɀMٙ�sRHљ��_	W��-�_=��C��TI��I�I�II�	F�`�JLA.�1[��VC��0�D�BO1�U�@i�B\JRK�U��	@DBL_�SMd�BM%`_D9LC�BGRV��0C��I��H_� �*COS+\�(LN�7+X>$C�9)�I�9)u*c,)�Z2 HƺMY@!�( "�TH&-�)THET=0�NK23I��"l=�A CB6CB=�C�A�B(261C�61�6SBC�T25GT	S QơC��aS$�" �4c#�7r#$DUD�EX�1s�t��B�6䆱�AQ|r�f$NE�DpIB U�\B5��	$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2��&�C�J�&!�VAHV�6H3�YLVhJVuKV��KV�KV�KV�KV�IHAHZF`RXM��wX�uKH�KH�KH�KH��KH�IO2LOAHOT�YWNOhJOuKO�KUO�KO�KO�KO�&�F�2#1ic%�d4GS�PBALANCE�_�!�cLEk0H_�%SP��T&�bc&�b>r&PFULC�hr��grr%Ċ1ky�U�TO_?�jT1T2Cy��2N&�v�ϰ ctw�g�p�0Ӓ~����T��O���� IN�SEGv�!�REV8�v!���DIF�鉳1l�w�1m
�OaB�q
����MIϰ�1��LCHWAR̭���AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|�n��ROBR�CR(����N��'�MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD�0�ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDX�Р  ��MOR^��t $-�U�� )��r�B���(�����Gؒu � $SIMULT ��~�x�� ���OBJE�`> �ADJUS>�1�OAY_Ik��D_�����C�_FIF�=�T� ��Ұ��{���p� �����p�@��DN�FRI��ӥT�ՓRO� ��E�{��͐OPWO�ŀv�0��SYSBU<�@ʐ$SOP�����#�U"��pPRUYN�I�PA�DH��D����_OU��=��qn�$}�IMKAG��ˀ�0P�q3IM����IN�q�~��RGOVRDȡ:���|�P~���Р�0�L_6p���i��R)B���0��M���SEDѐF� ��N`�M*����̰SL��`ŀw x $�OVSL�vSDI��DEXm�g�e�9Hw�����V� ~�N����w����Ûǖȳ�M��
͐�q<��� �x HˁE�F�AWTUS���C�08àǒ��BTM����If���4����(�.ŀy DˀEz�g���PE�r�����
���EXE��V��E�pY�$Ժ ŀz @ˁf��UP{�h�$�p��XN���9�H�� �PG"�{ h $SUB���c�@_��01\�MP�WAI��P����L�O��<�F�p�$�RCVFAIL_9C�f�BWD"�F����DEFSPup | Lˀ`�D��8� U�UNI���S���R`���_LZ�pP��͐P�ā}��� B�~���|�t�`ҲN�`KET��Jy���P� $�~��=�0SIZE] �h��{���S<�OR��?FORMAT/p 㰷 F���rEMR���y�UX���@�P�LI7�ā  �$�P_SWI���Ş_PL7�A�L_ �ސR�AR��B�(0C��Df��$Eh����C�_=�U� � �� ���~�J3x�0����TIA4��u5��6��MOM��@���� �B��AD��*��* PU70NRW��W� ��V����� A$PI�6���	� �)�4l�}69�Q���c�SPEED�PGq�7�D�> D����>tMt8[��SAM�`�p�>��MOV�� �$��p�5��5�D�	1�$2��������{�Hip�IN ?,{�F(b+=$�H*��(_$�+�+GAMM��f�1{�$GETH��ĐH�D����
^pOLIBR�ѝI��$HI��_��Ȑ*B6E��*8A$>G086LW=e6\<G9�686б�R��ٰV��?$PDCK�Q�"H�_����;"�� z�.%�7�4*�9�� �$IM_SRO�D�s"���H�&"�LE�O�0\H��6@�췀U� �ŀ��P�qUR_S�CR�ӚAZ��S_?SAVE_D�E��NO��CgA�Ҷ� �@�$����I��	�I � %Z[� ��RX"  ��m���"�q�'" �8�Hӱt�W�UPpS��рM��O� ��.'}q��Cg���@�ʣ����S�M�AÂ� � $PY���$WH`'�NG p���H`��Fb��Fb��Fb��PLM���	� 0(h�H�{�X��O��z��Z�eT�M���� pS��C��O__�0_B_�a��_%�� |S����@	�v��v@ �@���w�v��EM���%ˑS�fr�B�ːt��ftP��PM���QU� �U�Q���Af�QTH=�H{OL��QHYS�3ES�,�UE��B���O#��  -�P�0�|�gAQ���ʠu���O��ŀ�ɂv�-�8�A;ӝROG��a2D�E�Âv�_�Ā^Z�INFO&��+�h���bȜ�OI��� ((@SLEQ@/�#����@O�$o���S`c0O�0�j01EZ0NUe��_�AUT�Ab�CO�PY��Ѓ�{��@M��N�����1�P�
�M ��RGI�����3X_�Pl�$�����`�W��P��j@��G���EXT_CYCtb���p�����h�_NA�1!$�\�<�RO�`]�?� � m���POR�ㅣ���S�RVt�)����DI �T_l���Ѥ{�ۧP��ۧ �ۧ5٩6٩%7٩8���AS�B�-���$�F6����PL�A�A^�TAR��@E `�Z������<��d� ,(@F1Lq`h��@YNL����M�C���PWR�Ѝ�쐔e�DELiAѰ�Y�pAD#q��RQSKIP��� ĕ�x�O�`NT2!� ��P_x��� ǚ@�b�p1�1� 1Ǹ�?� �?��>���>�&�>�3�>�9��J2R;쐖 46��EX� TQ���� ށ�Q���[�KFд��w�RDCIf� �U`�X}�R�#%M!�*�0�)��$RGEA�R_0IO�TJBFcLG�igpERa�TC݃������2T�H2N��� 1�� �Gq TN�0 ����M����`Ib���EF:�1�� l�h���ENAB��lcTPE?@���!(ᭀ�� ��Q�#�~�+2 H�W���2�Қ���"�P4�F�X�j�3�қ{�@��������j�4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:Lj�7�ҟo@�����j�8�����"4Fj��SMSK�� � �+@��E�A�QR�EMOTE�������@ "1��Q�IIO�5"%I��tRd�9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C�ШP^��S232%�Sb��iDEVICEU�S#�R�RPARI�T�!OPBIT��Q��OWCON�TR��Qⱓ�RC�U� M�SUXTA�SK�3NB��0�$T�ATU�P�S�@@쐦F�6�_�PC�}�$FREEF�ROMS]p�ai�GsETN@S�UPDl��ARB73P%0����� !m$US�A���az9�L�ER1I�0f��pRY�5~"�_�@f�P�1�!�6WRK��D9�F9�~�FRIEND�Q�4bUF��&�A@TO�OLHFMY5�$�LENGTH_VT��FIR�pqC�@��E� IUFINt�R���RGI�1��AITI:�xGX���I�FG2�7G1`a����3�B�GPRR�DA��O_� o0e�I1�RER�đ�3&���T�C���AQJV�G(|�.2���F��1�!�d�9Z�8+5K�+5���N�y�L0�4�XS �0m�LN�T�3�Hz��89��%�4�3G���W�0�W�RdD �Z��Tܳ��K�a3d���$cV 2����1��I1H�02*K2sk3K3Jci �aI�i�a�L��SL���R$Vؠ�BV�EVDk��A bQ*R��� �,6Lc���9V2F{X/P:B��PS_�E���$rr�C�ѳ$A0��wPR���v�Ub�cSk�� {��6���� 0���VX`�!�tX`��0P��ꁂ
�5SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V��� �S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD��<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C���:c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQkfC�ѷ =	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�qG �X��ȑ����$.A$�1$�c1Ó���� x~�EGvpݓ��q!AR����09p>B�%��AXE���ROB��W�A4�_�-֣SY���!6��&MS�'WR���-1���STR��5�9�E�� 	5B��=QB90�@6������kOT�0o 	$�ARY8�w20����	%�FI��;�$�LINK�H��1��a_63�5�q�2XYZ"��;�q�3�@��1�2�8{0B�{D��� CFI��6G��
�{�_J��6��3a'OP_O4Y;5�Q#TBmA"�BC
�z��DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ ��@�5<:7�� +1�?0K�Mc�6�8Cb�vrb�4�ORQ��X�>8�#op�� ����wq�Uf�����T'OVE�Q��M;�@E#�UK#�UQ"�VW�Z Q�W���Tυ� ;� ���QH�!`�ҽ��U�Q��WkeK#kecXER��	GE	0��S�dAWaǢ:D���7!�!AX�rB! {q��1uy-!y �pz�@z�@z6Pz \Pz� z1v�y �y�+y�;y�Ky �[y�ky�{y��y��q�yDEBU��$����L�!º2WG�� AB!�,��S9V���� 
w��� m���w����1���1�� �A���A��6Q��\Q����!�m@��2CLAB3B�U�����So  ÐER��>�� � $�@� mAؑ!p�PO���Z�q0w�^�_MR}Aȑ� d  9T�-�ERR��TYz�B�I�V83@�cΑTOQ�d:`!L� �d2�]�X�}C[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	�SFZ�N_CFG_!� 4��?º�|�ų����@�ȲW ���\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(����$�!s�Q�g�P{RV �HELLĥ�� 56�B_BAS�!�RSR��ԣo ��#S��[��1r�%���2ݺ3ݺ4ݺ5*ݺ6ݺ7ݺ8ݷ���ROOI䰝0�0NLK!�CAB� ���ACK��IN��T�:�1�@�@ z�m�_�PU!�CO� ��OU��P� Ҧ) ��޶���TPFWD_�KARӑ��RE�~��P��(��QU�E�����P
��CSTOPI_AL������0&���㰑�0S#EMl�b�|�M��dЛTY|�SOK�}�D�I�����(���_�TM\�MANRQ�ֿ0E+�|�$K�EYSWITCH�&	���HE
�B�EAT����E� LQEҒ���U��FO������O_HOM��O�REF�PPARz��!&0��C+�9OA�ECO��B<�rIOCM�D8׆��]���8�` �# D�1����U��&��MH�»P�CFOR�C��� �P��O}M�  � @V�T�|�U,3P� 1-�T`� 3-�4�]��NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F�Ҿ���` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�r��J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7s�'��VP��UPD�� � ��|�԰��YS�LOǢ� �  z��и���o�E��`>�8^t��АALUץ�����CU���wFOqIgD_L�ӿuHI�z�I�$FILE_����t��$`�JvS�A��� h���E_BLCK�#�C>,�D_CPU<�{� <�o����tJr���R ��
PWl O� ��LA���S��������RUN F�Ɂ��Ɂ����F�����ꁬ��TBC�u�C� �X ;-$�LENi���v������I��G�L�OW_AXI�F)1��t2X�M����hD�
 ��I�� ���}�TOR����Dh��� L=��⇒�8s���#�_MA`�8ޕ��ޑTCV����T���&��ݡ�����J�����J����MDo���J�Ǜ ����
���2��� v���l��F�JK��VKi�hΡv�Ρ3��J0㤶ңJJڣJJ�A�ALң�ڣ��42�5z�&�N1-�9�(��␅�L~�_Vj�������� ` �GROU�pD��}B�NFLIC�����REQUIREa�EBUA��p����2¯�����c�ޞ� \��APKPR��C���
�;EN�CLOe�ɇS_M v�,ɣ�
����� ���M�C�&���g�_MG�q�C� �{�9����|�BRKz�NOL��|ĉ R��_LI�|��Ǫ�k�J����P 
���ڣ�����&���D/���6��6��8���r���� ���8�%�W�2�e�PATHa�z�p�z�=�hvӥ�ϰ�x�CN=��CA�����p�INF�UC��bq��CO�UM��YZ������q�E%���2������P�AYLOA��J2=L3pR_AN��<�L��F�B�6�R�{�R_F2LSHR��|�LOG��р��ӎ�>��ACRL_u��Ր����.���H�p��$H{���FLEX�
��J�� :�/����6�2�`����;�M�_�F16� ����n���������ȟ��Eҟ�����,� >�P�b���d�{�������������5�T��X��v���E ťmFѯ����� ��&�/�A�S�e�+p|�x�� � ��0����j�4pAT����6n�EL  �%ø�J���ʰJE��C�TR�Ѭ�TN��F�&��HAND_V�B[
�pK�� $F2{�6� �r�SWi��("U���� $$Mt�h�R ��08��@<b 35��^6�A�p3�k��q{9t�A(�̈p��A��A�ˆ0���U���D��D��P2��G��IST��$A4��$AN��DYˀ� {�g4�5D���v�6�v瀑�5缧�^�@��P �����#�,�5�>�(#�� &0�_��ER!V9�SQASYM$��] �����x�������_SHl����� ��sT�(����(�:�JA���S�cir��_VI�#Oh9�``V_UNI��td�~�J���b�E�b��d ��d�f��n�������H��uN���(!2�H������"Cq3EN� a�DI��>��ObtC�Dpx�� ��2IxQA����q ��-��s �� s������ ��OMMEB��rr/�TVpPT�P ���qe�i�A���P�x ��yT�P�j� $DUM�MY9�$PSm_��RFq�  ��:� s���!~q�� X����K�ST�s�ʰSBR��M�21_Vt�8$S/V_ERt�O��z����CLRx�A  O�r?p? Oր �� D $GLOB���#LO��Յ�$�o��P�!SYS�ADR�!?p�pT�CHM0 � ,x����W_NA���/�e���D�SR~��l (: ]8:m�K6�^2m�i7 m�w9m��9���ǳ��� ����ŕߝ�9ŕ�� �i�L���m��_�_��_�TD�XSCRE��ƀ�� ��ST�F���}�pТ6��C�] _v AŁ� 9T����TYP�r�@K��u�!u���-O�@IS�!��tvC�UE{t� �����H�S���!RSM�_�XuUNEXCcEPWv��CpS_�� {ᦵ�ӕ���÷����COU ��� [1�O�UET�փr|���PROGM� {FLn!$CU��cPO*q��c�I_�p}H;� � 8��.N�_HE
p��Q�~�pRY ?����,�J�*��;�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� D�C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!$��VSHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3�����w�2u�P{t9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+��t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2$��2���5��`�? ��ZAB�CS��  $��2��J�
���$$�CLAS������AB���'@@V�IRT��O.@AB�S�$�1 <E�� < *AtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v�����M@[�AXLրK�*B��dC  ���IN8��ā��PRE������LARM�RECOV �<I䂥�NG�� �\K	 A   �J�\�M@PPLIC��?<E�E��HandlingTool ��� 
V7.50�P/28[�  ��X0��
�_�SW�� UP*A� ��F0ڑ�����A���� 2)0��*A���:����(<FB �7DA5�� �'@Y0@<��None������� ��T��K*A4I/xl�_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ�:�i�n�����#B)B ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��e��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���oe�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� �0�5 	 �9 O�?$OO HO6K�2	���=9"��Q?55��C�PK��D3P������a�-4�O__|Z
�OG_�7�PO�� ȕ�6_��,xV�ADB���='�)
mc�:cpmidbgX�_`��S:�(�����Yp�_)o�S`��BBi�P�_mo8j��(�Koo�o9i�(��og�o�o�m�of�oGq:I�Z?DEF f8���)�R6pbuf.txtm�]n�@��Y��# 	`(Ж�Ao=L���zMC�21�=��9���4��=�n׾�Cz � BHBCCo��C|��Cq�D��C����C�{iSZE@D���F.��F���E⚵F�,E�ٙ�E@F��N�IU��I�?O�I<#I6�I�SYR���vqG���E�m�(�.��(�b(��<�q�G�x2ʄ�Ң �� a�D��j���E�e��EX��EQ�EJP� F�E�F�� G�ǎ^F� E�� FB�� H,- Ge�߀H3Y��� � >�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE d�O c
�(�;�"�G  <�6�z�R���?�j�C4��SZm� W��{�m��C��B-G�C�`@�$�q��T{�FP?ROG %i����c�I��� �Ɯ�f��KEY_TBL � �vM�u� �	
��� !"�#$%&'()*+,-./01c��:;<=>?@A�BC�pGHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������p����͓���������������������������������耇���������������������!j�LCK��.�j����STAT���_AUTO_DO����W/�INDT_'ENB߿2R��9��+�T2w�XSTO�P\߿2TRLl�L�ETE����_S�CREEN ~ikcsc���U��MMENU �1 i  <g\��L�SU+�U�� p3g���������� ��2�	��A�z�Q�c� ��������������. d;M�q� �����N %7]�m�� �/��/J/!/3/ �/W/i/�/�/�/�/�/ �/�/4???j?A?S? y?�?�?�?�?�?�?O �?O-OfO=OOO�OsO �O�O�O�O�O_�O_�P_Sy�_MANU�AL��n�DBCO�U�RIG���DB'NUM�p��<����
�QPXWORK 1!R�ү�_o�O.o@oRk�Q_AW�AY�S��GCP� ��=��df_AL�P�db�RY��������X_�p 1"�� , 
�^���o( xvf`MT�I^�rl�@�:sONTIM6������Zv�i�
õ�cMOTNE�ND���dRECO_RD 1(R�a��ua�O��q�� sb�.�@�R��xZ��� ����ɏۏ폄��� #���G���k�}����� <�ş4��X���1� C���g�֟�������� ӯ�T�	�x�-���Q� c�u����������>� ���)Ϙ�Mϼ�F� ࿕ϧϹ���:����� ��%�s`Pn&�]�o��� ��~ߌ���8�J���� ��5� ��k����ߡ� ��J�����X��|�� C�U�����������0�����	��dbTO�LERENCqdB�Ⱥb`L�͐PC�S_CFG )��k)wdMC:�\O L%04d.'CSV
�Pc�)s[A �CH� z�P�)~���hMR�C_OUT *��[�`+P SGN� +�e�r��#��10-MAY-�20 09:21~*V17-FEBj�19:09�k PQ�8��)~��`pa�m�?�PJPѬ�VERSION �SV2.�0.8.|EFLO�GIC 1,�[ 	DX�P7)�P�F."PROG_E�NB�o�rj ULS�ew �T�"_WRSTJNEp�V�r`d�EMO_OPT_�SL ?	�es
� 	R575 )s7)�/??*?<?'>�$TO  �-�l�?&V_@pEX�W�d�u�3PATHw ASA\�?��?O/{ICT�aF�o`-�gds�egM%&AST?BF_TTS�x�Y�^C��SqqF�PM�AU� t/XrMSWR.�i6.|S/�Z!D_N�O0__�T_C_x_g_�_�tSB�L_FAUL"0��[3wTDIAU 1�6M6p�A�12345678#90gFP?Bo Tofoxo�o�o�o�o�o �o�o,>Pb��S�pP�_ �� �_s�� 0`��� ��)�;�M�_�q��� ������ˏݏ��|)gUMP�!� �^��TR�B�#+�=�P�MEfEI�Y_TE{MP9 È�3@8�3A v�UNI�.(�YN_BRK �2Y)EMGDI�_STA�%WЕN�C2_SCR 3��1o"�4�F�X� fv���������#��ޑ14����)��;�����ݤ5�����x�f	u�ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/߭P�b�t��  ��xߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N���r������� ��������&8 J\n����� ���"`�FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/4 ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O?�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�O�O�o�o�o 
.@Rdv� �������� *�<�N�`�r����o�� ��̏ޏ����&�8� J�\�n���������ȟ�ڟ����H�ETM�ODE 16��]� ��ƨ�
R�d�v�נRRO�R_PROG �%A�%�:߽�  ���TABLE  A������#�L��RRSEV_NU�M  ��Q���K�S���_AU�TO_ENB  q��I�Ϥ_NOh�� 7A�{�R��  *������������^�+��Ŀֿ迄�HISO�͡I��}�_ALM 18.A� �;�����+�e�wωϛϭ����_H���  �A���|��4�TC�P_VER !�A�!����$EXTLOG_REQ�s�{�V�SIZ_�~Q�TOL  ͡{Dz��A Q�_BWD����r����n�_DI�� 9��}�z�͡m���STEP����4��_OP_DO����ѠFACTORY�_TUN�dG�E�ATURE :�����l�H�andlingT�ool ��  -� CEngl�ish Dict�ionary��O�RDEAA �Vis�� Mas�ter���96 �H��nalog �I/O���H55�1��uto So�ftware Update  ���J��matic �Backup��P�art&�gr�ound Edi�t��  8\ap�Cameraz��F��t\j6R��ell���LOA�DR�omm��sh�q��TI" ��cyo��
! o����pane�� �
!��tyle select��H59��nD���o�nitor��48�����tr��Rel�iab���adi�nDiagn�os"����2�2 u�al Check� Safety �UIF lg\a���hanced �Rob Serv> q ct\��lUser FrU���DIF��Ext�. DIO ��f�iA d��en]dr Err L@���IF�r��  �П�90��FCT�N MenuZ v�'��74� TP �In��fac � SU (G�=�p��k Exc�n g�3��Hig�h-Sper Sk]i+�  sO�H9 ~� mmunic!��onsg�teurh� ����V����^conn��2��{EN��Incr�stru���5.�fdKARE�L Cmd. L�?uaA� O�R�un-Ti� EnIv����K� ��+%��s#�S/W��74���License|T�  (Au* �ogBook(S�y��m)��"
�MACROs�,V/Offse6��ap��MH� �����pfa5�Mec�hStop Pr3ot��� d�b =i�Shif���/j545�!xr ��#��,[>b o�de Switc]h��m\e�!oz4.�& pro��4��g��Mul�ti-T7G��n�et.Pos Regi��z�}P��t Fun����3 Rz1��Nu!mx �����9m�1>�  Adjuj��O1 J7�7�* ��<���6tatuq1EIKRDMt�ot��scove�� ��@By- }Ouest1�$Go� �� U5\SNPX b"���YA�"Libr����#b�� �$~@h�pd]0��Jts in VCCM�����0�q  �u!��2 R�0��/I�08��T�MILIB�M J�92�@P�Acc�>�F�97�TPT�X�+�BRSQelZ0�M8 Rm��q%��692��Une�xceptr mo�tnT  CVV�P���KC����+�-��~K  II)��VSP CSXC��&.c�� e�"�� =t�@Wew�gAD Q�8bvr �nmen�@�iP�� a0y�0�pfG�ridAplay !� nh�@*�3R�1�M-10iA(B�201 �`2V" y F���scii��load��83 �M��l����Gua=r�d J85�0�maP'�L`���stua�Pat�&]$Cyc8���|0ori_ x%oData'Pqu���ch�1��g`� mj� RLJam�5����IMI De�-B(\A�cP" #�^0C  etk}c^0asswo%q.�)650�ApU��Xnt��Pven��CTqH�5�0�YELLOW BqO?Y��� Arc�0�vis��Ch�W�eldQcial44Izt�Op� ��gs�` 2@�a��p�oG yRjT1� NE�#HT� xyWb��! �p�`!gd`���p\� =P���JPN ARCP�*PR�A�� �OL�pSup̂f�il�p��J�� ��cro�670�1C~E��d��SS�pe�t�ex�$ �P� Soz7 t� ssagN5� <Q�BP:� �9 �"0�QrtQC��P�l0dpn�笔�r�pf�q�e�ppm�ascbin4p�syn�' ptx�]08�HELNC�L VIS PK�GS �Z@MB �&��B J8@I�PE GET_V�AR FI?S (�Uni� LU�OO�L: ADD�@2/9.FD�TCm���E�@DVp���`A��ТNO WTWTOEST �� f�!���c�FOR ��E�CT �a!� AL�SE ALA`�CPMO-130���� b D: HAN?G FROMg���2��R709 D�RAM AVAI�LCHECKS �549��m�VPC�S SU֐LIM�CHK��P�0x�F_F POS� F��� q8-12� CHARS�ER>6�OGRA ��Z@wAVEH�AME��G.SV��Вאn$���9�m "y�TR}Cv� SHADP��UPDAT k�0>��STATI���? MUCH ����TIMQ MOTN-003��@�OBOGUIDE? DAUGH���b8��@$tou� �@�C� �0��PATH|�_�MOVET��� R64��VMX�PACK MAY ASSERTjS޴�CYCL`�TA���BE COR �71�1-�AN��R�C OPTION�S  �`��APSwH-1�`fix��2�SO��B��XO򝡆��_T��	�i��0j���du�byz p cwa��y�٠HI������U�pb XSP�D TB/�F� \�hchΤB0���EmND�CE�06\Q��p{ smay In@�pk��L ���traff#�	� ���~1from �sysvar s�cr�0R� ��d�DJU���H�!A���/��SET ER�R�D�P7����N�DANT SCR�EEN UNRE�A VM �PD�D���PA���R�I�O JNN�0�F�I��B��GROUNנD Y�Т٠��h�SVIP 5�3 QS��DIGI?T VERS��k���NEW�� P0�6�@C�1IMAG��ͱ���8� DIx`���pSSUE�5���EPLAN J=ON� DEL���1�57QאD��CALLI���Q��m����IPND}�IMG� N9 PZ�19޴�MNT/��ES� ���`LocR HCol߀=��2�Pn� �PG:��=�M��c�an����С: �3D mE2vie�w d X��e�a1 �0b�pof �Ǡ"HCɰ�AN�NOT ACCE�SS M cpite$Et.Qs a� {loMdFlex)a�:��w$qmo G
�sA9�-'p~0��h0�pa��eJ AU�TO-�0��!ip�u@Т<ᡠIABL�E+� 7�a FPL�N: L�pl lm� MD<�VI�����WIT HOCv�Jo~1Qui�t�"��N��USB�@��Pt & rem�ov���D�vAxi�s FT_7�PG�ɰCP:�OS-�144 � h s� 268QՐOST��p  CRASH� DU��$P��W�ORD.$�LOgGIN�P��P:	��0�046 iss�ueE�H�: Solow st��c�`6����໰I�F�IMPR��SPOT:Wh4���N1�STY��0VMGqR�b�N�CAT��-4oRRE�� � 58�1��:%�R�TU!Pe -M a�SE:�@pp���AGp�L��m@al�l��*0a�OCB �WA���"3 CN�T0 T9DWro>O0alarm�ˀm0d t�M�"0�2�|� o�Z@OME�<�� ��E%  #1�-�SRE��M�st�}0g     �5KANJI5n�o MNS@�I�NISITALI�Z'� E�f�we���6@� dr�@ f�p "��SCII� L�afails� w��SYSTaE[�i��  � tMq�1QGro8�m n�@vA����&���n�0q��RWR=I OF Lk���� \ref"�
�u�p� de-rel}a�Qd 03.�0�SSchőbet�we4�IND e�x ɰTPa�DOȬ l� �ɰGi�gE�soperawbil`p l,��aHcB��@]�le�Q0cflxz�Ð���OS {����v4pwfigi GLA�$��c2�7H� la�p�0ASB� Ifz��g�2 l\c�0��/�E�� EX'CE 㰁�P���$i�� o0��Gd`]���fq�l lxt��EFal��#0��i�O�Y�n�CLOSn��SRNq1NT^��F�U��FqKP�AN�IO V7/ॠ1p�{����DB �0ء�ᴥ�ED��DE�T|�'� �bF�N�LINEb�BUG�T���C"RLIB���A��ABC J�ARKY@��� r7key�`IL���P�R��N��ITGAR
� D$�R �Er�� *�T��a�U�0��h�[�ZE V� �TASK p.vr�P2" .�XfJ��srn�S谥dIB�P	c���B/��B�US��UNN�  j0-�{��cR'���LOE�DIVS�C�ULs$cb����BW!��R~�W`P���&��IT(঱tʠ�{OF��UNEXڠ�+���p�FtE��S�VEMG3`NML� 505� D*�C?C_SAFE�P*�p �ꐺ� PET��8'P�`�F  !���IR����c i S�>� K��K�H �GUNCHG��S^�MECH��M��T*�%p6u��tP�ORY LEAKr�J���SPEg�D��2V 74\G�RI��Q�g��CTLN��TRe @�_��p ���EN'�IN�������$���r��T�3)�i�STO�A$�s�L��͐X	����q��Y� ��TO2�J m��0F<�K�����DU�S��O��3$ 9�J F�&�����SSVGN-18#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRKC�TR/"� �q\j5���_�Q�S�qINVJ0D ZO�Pݲ�� �s��г�Ui ɰ̒�a��DUAL� J�50e�x�RVO1/17 AW�TH!�Hr%�N�247%�5q2��|�&aol ���R���at�Sd�cU8���P,�LER��i�x�Q0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�cб���{�U��RO�P 2�b�pB��ITP4M��b !�AUt c0< � pl�ete�N@� �z1^qR635 (�AccuCal2zkA���I) "�(ǰ�1a\�Ps��ǐ � bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etaca2��AT���PC�`��슰�_p�.pc�!Ɗ��:�circB���5�tl��Bɵ��:�fm+�Ί�V�b��ɦ�r�upfrma.����ⴊ�xed�8�Ί�~�pedA�D ��}b�ptlib0B�� �_�rt�߄	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆�D����c�Ӳ�5�j>ʌ����tcȐ��	�r(����mm 1��T�#sl^0��T�mѡ�&#�rm3��ub Y��q�std}��pl�;�&�ckv�=�r�vaf�䊰��9�vi������ul�`�0fp�q� �.f��� d�aq; i Data� Acquisi
��n�
��T`���1�89��22� DMCM RR[S2Z�75��9 ?3 R710�o�59p5\?��T{ "��1 (D�T� nk@���������E Ƒȵ��Ӹ�et3dmm ��ER����gE��1�q\mo?۳�=(G����[(

�2�` ! ��@JMACRO���Skip/Of�fse:�a��V�4�o9� &qR662����s�H�
 6�Bq8����9Z�4_3 J77� 6�J783�o ���n�"v�R5IK�CBq2 PTLC�Zg R�3 (�s, ��������03�	зJԷ\�sfmnmc "MNMC����ҹ�%wmnf�FMC"�Ѻ0ª etmcr�� �8����� ,[>Df>�   874�\prdq>,jxF0���axisH�Process �Axes e�rol^PRA
�Dp� �56 J81j�5-9� 56o6� ��l�0w�690 98� �[!IDV�1��2(8x2��2ont�0�
 ����m2���?C���etis "I�SD��9�� FpraxRAM�P� D��defB�,�G�isbasicH�B�@޲{6�� 70U8�6��(�Acw: ������D
�/,��AMOX�� ��DvE��?�;T��>Pi� RAFM';�]�!PAM�V�W��Ee�U�Q'
bU�7y5�.�ceNe� �nterfaceh^�1' 5&!54�K<��b(Devam±��/�#���/<�Tane`"DNEWE���btpdnui �A�I�_s2�d_rsCono���bAsfj|N��bdv_arFv�f�xhpz�}w��hkH9xstc��gAp�onlGzv{�ff ��r���z�3{�q'Td>pcha�mpr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�!��pcchmp]aM�P&B�� �mpe�v�����pcs���YeS�� MacKro�OD��16Q! )*�:$�2U"_,��Y�(PC ��$_;�������o��J�geg{emQ@GEMSW�|~ZG�gesndy�<�OD�ndda��Sƕ�syT�Kɓ�su^Ҋ���n�m���L��O  ���9:p'�ѳ޲��spotplusp���`-�W�l�J�s��t[�׷p�key�ɰ�$��s��-Ѩ�m���\fea;tu 0FEAWD�oolo�srn '!2 p���a�As3���tT.� (N. A.)��!e!(�J# (j�,��o�BIB�oD -�.�n6��k9�"K��u[�-�_���p� "P�SEqW����wop "sEЅ�&�:� J������y�|��O8� �5��Rɺ���ɰ[� �X�������%�(
 ҭ�q HL�0k� 
�z�a!�B�Q�"(g�Q�����]�'� .�����&���<�!ҝ_�#��tpJ�H�~Z�� j�����y������2 ��e������Z����V� �!%���=�]�͂���^2�@iRV� on��QYq͋JF0� 8�ހ�`�	(^�dQueue���X\1����`�+F1tpvtsen��N&��ftpJ0v �RDV�	f���J1 Q���v�eyn��kvstk���mp��btkcl�rq���get�����r��`k�ack�XZ�st1rŬ�%�stl��~Z�np:!�`�� �q/�ڡ6!l�/Yr$�mc�N+v3�_`� ����.v�/{\jF��� �`�Q�΋ܒ�N50 (�FRA��+��͢f?raparm��Ҁ��} 6�J643�p:V�ELSE
�#�VAR $SG�SYSCFG.$��`_UNITS �2�DG~°@�4Jgfqr��4A�@FRL-� �0ͅ�3ې���L�0 NE�:�=�?@�8�v�9~Qx304��;�B�PRSM~QA�5T�X.$VNUM_�OL��5��DJ50�7��l� Functʂ"qwAP��琉�G3 H�ƞ�kP9jQ��Q5ձ� ��@jLJ zBJ[�6N�kAP�����S��"TPPRp���QA�prna�SV�ZS��AS8Dj5k10U�-�`cr�`8 ��ʇ�DJR`jYȑH  �Qm �PJ6�a21���48AAVM3 5�Q�b0 lB�`�TUP xbJ�545 `b�`61�6���0VCA�M 9�CLI�O b1�5 ����`MSC8�
rP� R`\sSTYL MNIN�`oJ628Q  �`�NREd�;@�`SC�H ��9pDCSU� Mete�`OR�SR Ԃ�a04 �kREIOC ��a5�`542�b9 vpP<�nP�a�`�R�`�7�`�MAS�K Ho�.r7 <�2�`OCO :��r�3��p�b�p���r0�X��a�`13\mn��a39 HRM"��q�q��LCH}K�uOPLG B��a03 �q.�pH�CR Ob�pCpP�osi�`fP6 i=s[rJ554�òp'DSW�bM�D�pqR��a37 }Rjr0 L�1�s4 �R6�7���52�r5 �2�r7� 1� P6���Re�gi�@T�uF�RDM�uSaq%�4�`930�uSNB�A�uSHLB̀\�sf"pM�NPI��SPVC�J5�20��TC�`"M�NрTMIL�I=FV�PAC W�poTPTXp6.%��TELN N M�e�09m3U�ECK�b�`UFR��`��VCOR��V�IPLpq89qSX9C�S�`VVF�J��TP �q��R62]6l�u S�`Gސ~�2IGUI�C���PGSt�\ŀH863�S�q�����q�34sŁ684`���a�@b>�3 :B抂1 T��96 :.�+E�51 y�q353�3�b1 ���b31 n�jr9 ���`�VAT ߲�q75� s�F��`�sAWSyM��`TOP u��ŀR52p���a809 
�ށXY q���s0 ,b�`885�QXрOLp}�"pE�v��tp�`LCMDў�ETSS���6� �V�CPE o�Z1�VRCd3
�NuLH�h��001m2�Ep��3 f��p��4� /165C��6�l���7PR��00�8 tB��9 -2[00�`U0�pF�1&޲1 ��޲2L"����p��޲4��5 �\hmp޲6 RB�CF�`ళ�fs�8� �Ҋ��~�J�7 OrbcfA�L�8\P0C����"�32m0u��n�K�Rٰn�5 5oEW
n�9 zΊ�40 kB��3 ��6ݲ�`00iB%/��6�u��7�u���8 µ������sU0��`�t �1 05\;rb��2 E��K���j���5˰��6A0��a�HУ`:�63�`jAF�_���F�7 ڱ�݀H�8�eHЋ��cUI0��7�p��1u��8u��9 73�������D7� ��5\t�97 ��8U�Q1��2��1�1:����h��1np�"��8�(�U1��\pyl���,࿱v ��B�85E4��1V���D�4��im��1�<���$>br�3pr�4@pGPr�6 B���цp���1����1�`͵15=5ض157 �2�у62�S����1�b��2����1Π"�2L���B6`�1<cf�4 7B�5 DR���8_�B/��18�7 uJ�8 06��90 rBn�1 �(��202 0E�W,ѱ2^��2��9�0�U2�p�2��2 �b��4��2�a"RiB����9\�U2�`xw�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`ڰR,:7 �2��V�2��5���2^��a^9���qr�����n�5����5᥁"�8Ha�Ɂ}�5B���5������`UA���� ��8�6 �6 S�0��5��p�2�#�529 ��2^�b1P�5�~�2`���&P5���8��5��u�!�5\��ٵ544��5��	R�ąP nB^z�c (�4�����SU5J�V�5��1�1@^��%�����5 �b21��gA��5m8W82� rb��95N�E�5890r�: 1�95 �"�� ����c8"a��|�L (���!J"5|6��^!"�6��B�"8�`#���+�8%�6B�AM�E�"1 iC��622�Bu�6V��d� �4��84�`ANR�SP�e/S� �C�5� �6� ��� \@� �6� �V� 3t��?� T20CA�R���8� Hf� 1DH��� AOE� ��w ,[|�� �0X\�� �!64K��ԓ�rA� �1 (M-7�!/50T�[PM��P�Th:1�C�#P�e� �3�0� 5`M�75T"� �D8p�! �0Gc� u�4��i1�-710i�1� S�kd�7j�?6�:-HS,� �RN�@�UB��f�X�=m75sA*A6an���!/CB�B2.6A �0;A�C�IB�A�2�QF1�UB2:�21� /70�S� �4����Aj1�3p����r#0 B2\m*A@C��;bi"i1K��u"A~AAU� imm7c7��ZA@I�@�Df�A�D5*A�E� #0TkdR1�35Q1�" *�@�Q�1�QC)P�1 *A�5*A�EA�5B�4>\77
B7=Q�D�2H�Q$B�E7�C�D/qA	HEE�W7�_|`jz@@� 2�0�Ejc7(�`�E"l7�@7�A
1��E�V~`�W2%Q�R9\ї@0L_�#��� �"A���b��H3s=rA/2�R5nR4�7�4rNUQ1ZU�A�s\m9
1M92L2�!F!t^Y�ps� 2ci��-?�qhimQ�t  w0 43�C�p2�mQ�r�H_ �H20�Evr�QHsXBFSt62�q`s����� ��Pxq350_�*A3I)�2�d�u0X�@� '4TX�0�pa3i1A3sQ25L�c��st�r�VR1%e�q0
��j1��O 2 �A�UEiy�.�‐� �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ�� qA!Pvs� 5	15aU ���?PŅ���ဝQG9A6�zS*�7�q�b5�1����Q��00	P(��V7]u�aitE1 ���ïp?7� !?�z���rbUQRB1P�M=�Qa9��H��QQ�25L�������Q���@L��8ܰ��y0�0\ry�"R2B�L�tN  ��w� �1Df>�2�qeR�5���_bx�3�X]1m1lcqP!1�a�E�Q� 5F����!5���@M-16 Q�� f���r��Q�e�� ��� PN�LT_`�1��i1��9453�p�@�e�|�b1l>�F1u*AY2�
��R8`�Q����RJ�J3�D}T� 85
Qg�/0�� *A!P�*A�Ð𫿽�Y2ǿپ6t�6=Q����Pȓ��� AQ� g�*ASt]1^u�a jrI�B����~�|I��b��yI�\m�Qb�I �uz�A�c3Apa9q� B6S��S��m����}�85`N�N�  �(M���f1����6����161��5�s`�SC��U��A�����5\set036c����10�y�#h8��a6��6��9r�2HS ���Er���W@}�a��I�lB� ��Y�ٖ�m�u�C������5�B��B��h `�F���X0���A:���C�M��AZ��@��4��6i����� e�O�- 	���f1��F ������1F�Y	���T6HL3��U66~`���Ur�dU�9D20Lf0 ��Qv� ��fjq��N� �����0v
� ��i	��	��72lqQ2�������� \chngmove.V���d���@2l_arf	�f~�� 6������9C�Z��0�~���kr41 S���0��V��t����8��U�p7nuqQ%��A]��V�1\�Qn�BJ�2W�E�M!5���)�#:�648��F�e50S�\� �0�=�PV���e�� ����E������m7shqQSH" U��)��9�!A��(����� ,[s>�ॲTR1!�L��,�60e=�4F�d����2��	 R-�� ���������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2��"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D�� �5V��@2cVE��pȖ�T��pt갖�1L ~E�#�F�Q��9E�#Dce/��RT��59�� �	�A�EiR�������9\m20�20 ��+�-u�19r4�`� E1�=`O9`�1"ae��O�2��_$W}am41�4�3�/d?1c_std��1�)�!�`_T��r�_ 4\jdg�a�q�P J%!~`-�r�+bg8B��#c300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W �"PsA��e��� �t�i�P�W.�� c�FX.�e�kE1�4�44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�A Pf��coWo!\�[2a��2A;_2��QW2�bF�(�V11ă23�`��X5�Ra2�1�J*9�a:88�J9X�l5�m1a`첚��*���(85�& �������P6����R,52&A����,8fA9IfI50\u�z��OV
�v��}E֖J0���Y>� 16r�C �Y��;��1��L���A q�&ŦP1��vB)e��m�����1p� .�1Df>�27�F��KAREL Us�e S��FCTN<��� J97�FA+�� (�Q޵�p%�L)?�Vj9F?(�j�R�tk208 "Km�6Q�y�j��iæP�r�9�s#��v�kr;cfp�RCFt3����Q��kcctme��!ME�g����6�mWain�dV�� ��Cru��kDº�c��0�o����J�dt�F9 �»�.vrT�f�����E%�!��5�FR�j73B�K���UtER�HJ�O  J��# (ڳF���F�q� Y�&T��p�F�z��19�tkvBr���V�h�9p�E�y�<�k������p��;�v���"CT�� f����)�
І��)� V	�6���!��qFF ��1q���=�����O�@?�$"���$��je����TCP Aut��r�<520 H5n�J53E193��9��96�!8��9���	 �B574��5�2�Je�(�� Se%!Y�����u��ma>�Pqtool�ԕ������conr�el�Ftrol �Reliable��RmvCU!��H51������ a55�1e"�CNRE ¹I�c�&��it��l\sfutst "UTա��"X�\u��g@�i�6Q]V�0�B,Eѝ6A�  �Q�)C���X��Yf�hI�1|6s@6i��T6IU��vR�d�
$ae%1��2�C58�E6��8�Pv�iV4OFH�58SOeJ� mvBM6E~O58�I�0�E �#+@�&�F�0���F �P6a���)/++�</>N)0\tr1������P ,[>ɶ�rmwaski�msk�a$A���ky'd�h	A	��P�sDispla�yIm�`v����J887 ("A��+Hyeůצprds�ҨIϩǅ�h�0pl�2"�R2��:�Gt�@��PRD�TɈ�r�C�@�Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@��^Sp��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@�P�firmQ����P@p�2�=bk�6�r�3��6��tppl��PAL���O�p<b�ac�q 	��g1J�U�d�J��gait_9e��Y��&��Q���	�Sha�p��eratio�n�0��R674�51j9(`sGen@�ms�42-f��r�p`�5����2�rsgl��E��p�G���qF�20�5p�5S���Ձ�re�tsap�BP�O�\}s� "GCR��z�? �qngda�AG��V��st2ax�U��Aa]��bad��_�btputl�/�&�e���tpli1bB_��=�2.����5���cird�v�sqlp��x�hex���v�re?�Ɵx�key�v�pm��x�sus$�6�gcr���F������[�q27j9�2�v�ollis�mqSk�9O�ݝ� �(pl.���t��p!o��29$Fo8��cg�7no@�tptcls` CLS�o�b�F\�km�ai_
�s>�v�o	�t�b���ӿ�E�H��6�1e_nu501�[m���utia|$cal�maUR��CalMwateT;R51%�i=1]@-��/V� ���Z�� �fq1�9 "�K9E�L����2m�CLMTq�S#��3et �LM3!}t �F�c�nspQ�<c���c_moq��� ��c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 �̆�N�ve��C�cl�m�&Ao# �|$fi�nde�0S�TD ter FiLANG���R��
��n3���z0Cen���r, ������J����� � ��K��Ú�=���_�����r� "FNCDR�� 3��f��tguid�䙃N�."��J�tq�� ��� ����������J����_������c��	m��Z��\fndrA.��n#>
B2p��>Z�CP Ma������38A��� c��6� (���N�B���@���� 2�$�81�B�m_���"ex� z5�.Ӛ��c��0bSа�efQ���	��RBT;�OPTN �+#Q� *$�r*$��*$r*$%/ s#C�d/.,P�/0*ʲDPN��$����$*�Gr�$k E�xc�'IF�$MA�SK�%93 H5��%H558�$548 H�$4-1�$�d�#1(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9j0�"M�49�4  ���4�4tpsh���4�P�4- DQ�� �3�Q�4�R�4�pR@%0�2�r�4.b
E\���5�A�4��3adq}\�5K979":E��ajO l "DQ ^E^�3i�Dq ��4�ҲO ?R�? ��q@�5��T��3rAq�OF�Lst�5~��7p�5`��REJ#�2�@av^E�ͱ�F���4��.�5y� N� �2il(iqn�4��31 JH1��2Q4�251ݠ�4r'mal� �3)�RE o�Z_�æOx����4��8^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4$�REM���4yݱ"u<@�RER5932fO��47Z��5lity�,�U��e"Dil�\�5��o ��79�87�?�25 �3hk910�3��FE�0�=0P_�Hl\mhm �5��qe�=$�^��
E��u�IAympt�m�U��BU��vst e�y\�3��me�b�Dv I�[�Qu�:F�Ub�*_0�
E,�su��_	 Er��ox���4huse�E-�?�sn�������FE��,�Gbox�����c݌ ,"�������z���M��g��pdspw )�	��9���b���(��1���c�� Y�R�� �>�P���W�@�������'�0ɵ��[��͂��� � � ,[@�� �A�bu�mpšf��B*�BCox%��7Aǰ60�pBBw���MC� (6��,f�t I�s� ST��*��}B������w��"BBF�
�>�`���)��\�bbk968 "��4�ω�bb�9�va69����etb�Š��X�����ed�	�F��u�f� �s�ea"������'�\���,���b�ѽ�oH6�H�
�x�$�f����!y���Q[�! toperr�fd� �TPl0o� Rec�ov,��3D��R/642 � 0��C@�}s� N@��(U�rro���yu2r���  �
 � ����$$CL~e� ������������$z�_�DIGIT��������.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�o$j��+c:PR�ODUCTM�0\�PGSTKD��V�&ohozf99��D����$FEAT_INDEX���xd�� � 
�`ILEC�OMP ;����#��`�cSET�UP2 <�e��b�  N ��a�c_AP2BC�K 1=�i G �)wh0?{%&c����Q�xe% �I�m���8� �\�n����!���ȏ W��{��"���F�Տ j���w���/�ğS�� �������B�T��x� �����=�үa����� �,���P�߯t���� ��9�ο�o�ϓ�(� :�ɿ^���Ϗϸ� G���k� �ߡ�6��� Z�l��ϐ�ߴ���U� ��y����D���h� �ߌ��-���Q����� �����@�R���v�� ��)�����_����� *��N��r�� 7��m�&��3\�i
pP }2#p*.VRc�*��� /��PC/1/�FR6:/].��/+T�`�/�/F%��/�,�`r/?�*#.F�8?	H#&?�e<�/�?;STM� �2�?�.K �?�=�iPenda�nt Panel�?;H�?@O�7.O�?8y?�O:GIF�O�O��5�OoO�O_:JPG _J_�56_�O_�_��	PANEL1'.DT�_�0�_�_�?O�_2�_So�W Ao�_o�o�Z3qo�o@�W�o�o�o)�Z4�o�[�WI��
�TPEINS.XSML��0\����qCustom� Toolbar�	��PASSW�ORDyFR�S:\L�� %�Password Config�� �֏e�Ϗ�B0��� T�f����������O� �s������>�͟b� �[���'���K��� �����:�L�ۯp��� ��#�5�ʿY��}�� $ϳ�H�׿l�~�Ϣ� 1�����g��ϋ� ߯� ��V���z�	�s߰�?� ��c���
��.��R� d��߈���;�M��� q������<���`��� ����%���I������ ��8����n��� !��W�{" �F�j|�/ �Se��/�/ T/�x//�/�/=/�/ a/�/?�/,?�/P?�/ �/�??�?9?�?�?o? O�?(O:O�?^O�?�O �O#O�OGO�OkO}O_ �O6_�O/_l_�O�__ �_�_U_�_y_o o�_ Do�_ho�_	o�o-o�o Qo�o�o�o�o@R �ov��;�_ ���*��N��G� �����7�̏ޏm�� ��&�8�Ǐ\�돀�� !���E�ڟi�ӟ��� 4�ßX�j�������� įS��w������B��#��$FILE_�DGBCK 1=���/���� ( �)�
SUMMARY�.DGL���MD�:�����Di�ag Summa�ry��Ϊ
CONSLOG��������D�ӱConso?le logE�ͫ���MEMCHECCK:�!ϯ���X��Memory D�ata��ѧ�{�)��HADOW�ϣϵ�J���Sh�adow Cha�ngesM�'�-��)	FTP7�Ф�3ߨ���Z�mment TBD���ѧ0=4)ET?HERNET��������T�ӱEth�ernet \�f�iguratio�nU�ؠ��DCSV�RF�߽߫������%�� veri?fy all��'��1PY���DIF�F�����[���%=��diff]�������1R�9�K���c ���X��CHGD������cB��r����2Z8AS� ��GD���k��qz��FY3b8I[� �/"GD���s/�����/*&UPDATES.� �/��?FRS:\�/�-�ԱUpdate?s List�/���PSRBWLD.CM(?���"<?�/�Y�PS_ROBOWEL��̯�?�?� �?&�O-O�?QO�?uO OnO�O:O�O^O�O_ �O)_�OM___�O�__ �_�_H_�_l_o�_�_ 7o�_[o�_lo�o o�o Do�o�ozo�o3E �oi�o���R �v���A��e� w����*���я`��� ������O�ޏs�� ����8�͟\����� '���K�]�쟁���� 4���ۯj������5� įY��}������B� ׿�x�Ϝ�1���*� g�����Ϝ���P��� t�	�ߪ�?���c�u� ߙ�(߽�L߶��߂� ��(�M���q� �� ��6���Z������%� ��I���B�����2�����h����$FoILE_� PR� ���������MDO?NLY 1=.��? 
 ���q ����������~ %�I�m �2��h��!/ �./W/�{/
/�/�/ @/�/d/�/?�//?�/ S?e?�/�??�?<?�? �?r?O�?+O=O�?aO �?�O�O&O�OJO�O�O �O_�O9_�OF_o_
?VISBCKL6>[*.VDv_�_>.PFR:\�_�^�.PVisio�n VD file�_�O4oFo\_joT_ �oo�o�oSo�owo �oB�of�o� +������� +�P��t������9� Ώ]�򏁏��(���L� ^�������5���ܟ k� ���$�6�şZ���~�����
MR_�GRP 1>.�L��C4  B���	 W������*u����RHB ���2 ��� ��� ���B����� Z�l���C���D��������Ŀ��K��N�J��I���T��:F�5U�P�򶲿�ֿ �E�M.G��E$��;n���:G��@O����@�Tf@���fy�@���m@���*λ?� F@ ��������J��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<,6\b�π+�&�(�a�L߅�p�A��A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�PS@�P��J����߿�#�B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�O�гߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������0u[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U�� 
//./�v���/ ���/�/�/�/�/� !?3?E?W?i?�/?�? �?�?�?�?�?��� AO�?eO�/�O�O�O�O �?�O�O__+_NO�O J_s_�_�_�_�_
OO .OoB_'ovOKo]ooo �oP_>o�o�o�o�oo �o5GYk}�_ �_�_��8o�� 1�C�U�$y������� �ӏf���	��-�?� ����Ə���ϟ �����;�M�_� q���.�(���˯ݯ� �P�b�t�����m��� ������ǿٿ����� !�3�E�h��{ύϟ� �����$�6�H�J�/� ~�S�e�w߉ߛ�jϿ� �������*߬�=�O��a�s��YT_ER�R J5
���P�DUSIZ  j��^J����>��?WRD ?t���  guest}��%�7��I�[�m�$SCDMNGRP 2Ktw�������V$�K�� 	�P01.14 8~��   y�����B   � ;����� ����������
 �������?�����~����C.gR|����  i  ��  
��������� +�������
���l �.r���"�l��� m
d����|��_GROU��]L�� �	�����07EQUPD'  	պ�J��TYa ����T�TP_AUTH �1M�� <!iPendany���6�Y!K?AREL:*��
-KC///A/ �VISION �SETT�/v/� "�/�/�/#�/�/
? ?Q?(?:?�?^?p>�CTRL N�����5�
�F�FF9E3�?��FRS:DEFA�ULT�<FA�NUC Web �Server�:
 �����<kO}O�O�O��O�O��WR_CONFIG O��� �?��IDL_CPU_PC@��B��7P�BHUMIN(\��<T?GNR_IO�������PNPT_S_IM_DOmVw[�TPMODNTO�LmV �]_PRT�Y�X7RTOLNK 1P����_o�!o3oEoWoio�RMA�STElP��R�O�_CFG�o�iUO���o�bCYCLE��o�d@_ASG s1Q����
 ko ,>Pbt��� ������sk�bNUM����K@�`�IPCH�o��`R?TRY_CN@oR<��bSCRN����Q��� �b�`�b�R���Տ��$J�23_DSP_E�N	����OB�PROC�U�iJ[OGP1SY@��?8�?�!�T��!�?*�POSRE��zVKANJI_@�`��o_�� ��T�L��6͕����CL_�LGP<�_���EYL_OGGIN�`�����LANGU�AGE YF7ReD w���LG��YU�?⧈�x� ������=P��'�0��$ NM�C:\RSCH\�00\��LN_D?ISP V��
�0�������OC�R.R�DzVTA{�OGB?OOK W
{��`i��ii��X������ǿٿ�����"��6	h������e�?�G_BUF/F 1X�]��2	աϸ������� ����!�N�E�W߄� {ߍߺ߱�����������J���DCS� Zr� =����^�+�ZE������|��a�IO 1[
{G ُ!� �!� 1�C�U�i�y������� ��������	-A Qcu�����z��EfPTM  �d�2/ASew �������/ /+/=/O/a/s/�/�/���SEV���.�TYP�/0??y͒�RS@"�|�×�FL 1\
������?�?�?�?0�?�?�?/?TP6���">�NGNA�M�ե�U`�UPSF��GI}�𑪅mA�_LOAD�G �%�%DF_�MOTN���O�@MAXUALRM<���J��@sA�Q����(WS ��@C �]m�-_����MP2�7�^
{k ر�	�!P��+ʠ�;_/��Rr�W�_�WU�W�_�� �R	o�_o?o"ocoNo so�o�o�o�o�o�o�o �o;&Kq\� x������� #�I�4�m�P���|��� Ǐ���֏��!��E� (�i�T�f�����ß�� ӟ���� �A�,�>� w�Z�������ѯ���� د���O�2�s�^� ������Ϳ���ܿ��'��BD_LDXD�ISAX@	��ME�MO_APR@E {?�+
 �  *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT�� Q�c�Ϝ߇��ߧ��� ��w����>�)�b�t� [����{������� ���:���I�[�/��� ���������o����� 6!ZlS�� s����2� AS'�w��� �g��.//R/d/��_MSTR �`�-w%SCD 1am͠L/�/H/�/�/ ?�/2??/?h?S?�? w?�?�?�?�?�?
O�? .OORO=OvOaO�O�O �O�O�O�O�O__<_ '_L_r_]_�_�_�_�_ �_�_o�_�_8o#o\o Go�oko�o�o�o�o�o �o�o"F1jU g������� ��B�-�f�Q���u�𮏙�ҏh/MKCF/G b�-㏕"�LTARM_��c�L�� �σQ�N�<�METP�UI�ǂ���)N�DSP_CMNT�h���|�  d�.��ς�ҟܔ|�_POSCF�����PSTOL 1e�'�4@�<#�
 5�́5�E�S�1�S�U� g�������߯��ӯ� ��	�K�-�?���c�u������|�SING_?CHK  ��;�/ODAQ,�f��Ç���DEV 	�L�	MC:!�HOSIZEh��-��TASK %6��%$123456�789 �Ϡ��T�RIG 1g�+ l6�%���ǃ��0���8�p�YP[� ���EM_INF �1h3� �`)AT&F�V0E0"ߙ�)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ�����ԁH�����A���A�I�q�,��|����  ���ߵ�����J��� n������W������� ����"����X�� /����e���� ��0�T;x�= �as��/�,/ c=/b/�/A/�/�/ �/�/��?��� ^?p?#/�?�/�?s?}/ �?�?O�?6OHO�/lO ?1?C?U?�Oy?�O�O 3O _�?D_�OU_z_a_��_�ONITORG ?5�   �	EXEC1TɃ�R2�X3�X4�XQ5�X���V7�X8�X9Ƀ�RhBLd�RLd �RLd�RLd
bLdbLd "bLd.bLd:bLdFbLcU2Sh2_h2kh2whU2�h2�h2�h2�hU2�h2�h3Sh3_h�3�R�R_GRP?_SV 1in����(����C?B�PP�A4�>%���gY�>r3��x�_D=R^���PL_NAME� !6��p�!�Default� Persona�lity (from FD) ��RR2eq 1j)TUX)TX��q��X dϏ8�J�\� n���������ȏڏ� ���"�4�F�X�j�|������2'�П��� ��*�<�N�`�r��<��������ү������,�>�P�b� �R�dr 1o�y �\��, �3��~�� @D�  ��?�����?䰺�㱏A'�6����;��	lʲ	 �xJ����� ��< �"�� ��(pK�K� ��K=*�J����J���J�V���Z�����rτ́p@j��@T;f���f���ұ]�l��I�o��������������b��3���o�  ��`�>�����bϸ�z��{Ꜧ���Jm��
� B�H�˱]����q�	� p��  P�pQ�p�>�p|  Ъ�g����c�	'� �� ��I� ��  ����:��È
�È=����"�nÿ�	�ВI�  �n @@B�cΤ�\��ۤ���q�y�o�N���  �'�����@2��@�����/��C��C�C�@� C������
��A�W�@<�*P�R�
h�B�b�A��j�����:����Dz۩��߹������j��( ?�� -��C�`��'�7�����q��Y����� �?�ff ��gy ����o��:a��
>+�  PƱj�(����7	����|�?���xZ�p<
6b�<߈;܍��<�ê<� �<�&Jσ�A�I�ɳ+���?ff�f?I�?&�k�@��.��J<?�`�q�.�˴ fɺ�/��5/���� j/U/�/y/�/�/�/�/��/?�/0?q��F �?l??�?/�?+)��?�?�E�� E��I�G+� F� �?)O�?9O_OJO�OXnO�Of�BL޳B� ?_h�.��O�O��%_�O L_�?m_�?�__�_�_x�_�_�
�h�Îg>��_Co�_`goRodo�o�GA�ds�q�C�o�o�o|����$]Hq�m��D��pC����pCHmZZ7t����6q�q��ܶN'�3�A�A�AR1�AO�^?�$��?�K/�±
�=ç>�����3�W
=�#�\W��e��9������{����<���(�B��u��=B�0�������	L��H�F�G����G��H��U`E���C��+���I#��I��HD��F��E��R�C�j=��
�I��@H�!�H�( E<YD0q�$��H� 3�l�W���{������� �՟���2��V�A� z���w�����ԯ���� ����R�=�v�a� �����������߿� �<�'�`�Kτ�oρ� �ϥ��������&�� J�\�G߀�kߤߏ��� ��������"��F�1� j�U��y������� �����0��T�?�Q�t���(���3/�E����u�������q3�8�x����q4Mgs�&IB+2D�a���{�^ ^	������u%P2P7Q4_A���M0bt��R�������/   �/�b/P/�/ t/�/ *a)_3/�/�/�%1a?�/?;?8M?_?q?  �?�/��?�?�?�?O 2 �F�$�vGb��/�A��@�a�`�qC��C@�o�Ot���K�F� DzH@��� F�P D�!��O�O�ys<O!_�3_E_W_i_s?��W�@@pZ�42�2!2~
 p_�_�_�_	oo -o?oQocouo�o�o�o��o��Q ��+���1��$MSK�CFMAP  ��5� ��6�Q�Q"~�cONR�EL  
�q3�bEXCFE�NB?w
s1uXqF�NC_QtJOGO/VLIM?wdIpMr]d�bKEY?w�u]�bRUN�|�u��bSFSPDT�Y�avJu3sSIG�N?QtT1MOT��Nq�b_CE_�GRP 1p�5s\r���j����� T��⏙������<� �`��U���M���̟ ��🧟�&�ݟJ�� C���7�������گ��������4�V�`TC�OM_CFG 1�q}�Vp�����
�P�_ARC_\r�
jyUAP_CP�L��ntNOCHE�CK ?{ 	r��1�C� U�g�yϋϝϯ����������	��({NO_?WAIT_L�	u6M�NTX�r{�[�m�_ERRY�29sy3� &�������r�c� �촯T_MO��t��,� �5j�2�PA�RAM��u{��	�[���u?�� �=9@345678901��&���E� W�3�c�����{������������=��UM_RSPA�CE �Vv��$?ODRDSP����jxOFFSET_�CARTܿ�DI�S��PEN_FILE� �q��c֮��OPTION_I�O��PWORK� v_�ms  �P(�R�Q
�j.j	 ��Hj&6$�� RG_DSBOL  �5Js�\���RIENTT5O>p9!C��Pq�fA� UT_SIM�_D
r�b� V~� LCT ww��bc��U)+$_PEsXE�d&RATp Тvju�p��2X�j)TUX)TX�##X d-�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	OO-O?O�H2�/oO�O �O�O�O�O�O�O�O_]�<^O;_M___q_�_ �_�_�_�_�_�_o���X�OU[�o(ҿ�(���$>o�, ��Ip~B` @D�  Ua?�[cAa?p]a]��DWcUa쪋l;��	lmb�`�xoJ�`�p����a�< ���`� ��b��H�(��H3k7H�SM5G�22G���Gp
��
���'|��C%R�>�>q�Gsua|T�3���  �4spBpyr  ]o��*SB_���{�j]��t�q� ��rna �,����6  ���PQ�|�N�M�,k���	'�� � ��I�� �  �=�%�=��ͭ����ba	���I  ?�n @��~ ���p��Y����*�9N	 W�  '!o�t:q�pC	 C�@@s�Bq�|��� m�
��!�h@ߐ�nH����*�B	 �A���p� �-�qbz��P��t�_�������( �� -��恊�n��ڥ[A]Ѻ�b4�'!�5�(p �?�ff � ��
����OZ�DR*�85�z���>΁'  Pia��(5����@���ک�a�c�dF#?���5�x��*�<�
6b<߈;�܍�<�ê<� <�&�o&�)�A�lcΐI�*��?fff?�?&�c���@�.u?J<?�`��Y ђ^�nd��]e��[g�� Gǡd<����1��U� @�y�dߝ߯ߚ����� ��	���-������&����"�E�� E�~�G+� Fþ� ����������&��PJ�5��bB��AT� 8�ђ��0�6���>��� J�n�7��[m<�0��h��1��>�M�I
0�@��A�[���C-�)��?���� /�Y�Ē��Jp��vav`CH/������}!�@I�Y�'�3�A�A�AR1�AO�^?�$��?����±
�=ç>�����3�W
=�#�\���+e��ܒ������{����<���.(�B��u��=B�0�������	�*H�F�G����G��H��U`E���C��+�-I#��I��HD��F��E��R�C�j=U>
�I��@H�!�H�( E<YD0/�?�?�?�? �?O�?3OOWOBOTO �OxO�O�O�O�O�O�O _/__S_>_w_b_�_ �_�_�_�_�_�_oo =o(oaoLo�o�o�o�o �o�o�o�o'$ ]H�l���� ���#��G�2�k� V���z���ŏ���ԏ ���1��U�g�R��� v�����ӟ�������t-��(���������a�����Q�c�,!3�8�x}���,!4Mgs�����ɢIB+կ篴a���{�� �A�/�e�S���w��%P!�P��������7��ӯ�ϑ�R�9�Kτ�oχϓϥ�  ���χ����)� �M������z���{��ߛ���ߒߤ���8����  )�G��q�_���2 �F�$�&Gb����n�[ZjM!C�s�@j/�A�S�=�F� Dz���� F�P D�!�W����)������������x?��W�@@
9�=�=��=��
 v���� ���*<N�`�*P ���˨��1��$PAR�AM_MENU �?-���  DE�FPULSEl�	WAITTMO{UT�RCV�� SHELL�_WRK.$CU�R_STYL��,OPT�/P�TB./("C�R_DECSN���, y/�/�/�/�/�/�/? 	??-?V?Q?c?u?�?��USE_PRO/G %�%�?�?.�3CCR������7_HOST �!�!�44O�:T ̰�?PCO)ARC�O>�;_TIME�XB�  �GDE�BUGV@��3GI�NP_FLMSKĵO�IT`��O�EPG�AP �L��#[CyH�O�HTYPE����?�?�_�_�_ �_�_oo'o9obo]o oo�o�o�o�o�o�o�o �o:5GY�} ����������1�Z��EWORD� ?	7]	R}S`�	PNS��$��JOE!>��TEs@WVTRACECTL 1x-�� ������ɆDT �Qy-���Do � ��,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�T� (�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_j��_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\�n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�_����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv��������//"#�$PG�TRACELEN�  #!  �_�" �8&�_UP z����g!o S!�h 8!_CFG �{g%Q#"!x!��$J �#|"DEFS_PD |�,!!�J �8 IN T_RL }�-" �8�%�!PE_CO�NFI� ~g%'�g!�$�%�$WLID�#�-74?GRP 1�7Q!��#!A ����&ff"!A+3�3D�� D]� CÀ A@+6
�!�" d�$�9�9*1~*0� 	 +9p�(�&�"�? ´	C�?�;B@3AO�?O�IO3OmO"!>�T?�
5�O�O�N�O� =��=#�
�O_�O_J_5_n_ Y_�O}_�_y_�_�_�_�  Dzco" 
 oBo�_Roxoco�o�o �o�o�o�o�o>�)bM��;
V�7.10beta�1�$  A��E�rӻ�Ay " �p?!G��q/>���r��0�q��ͻqBQ��qA\�p�q�4�q�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏��� 4��1�j�U���y��� ��֟������0�� T�?�x�c�������ү ����!o�,�ۯP�;� M���q�����ο��� ݿ�(��L�7�p�+9<��sF@ �ɣ� �ϥ�g%������+� !6I�[߆������ߵ� ����������!��E� 0�B�{�f������ �������A�,�e� P���t���������� ��=(aL^ ������� '9$]�Ϛ��ϖ �������/<�5/ `�r߄ߖߏ/>�/�/ �/�/�/?�/1??U? @?R?�?v?�?�?�?�? �?�?O-OOQO<OuO `O�O�O�O�O���O_ �O)__M_8_q_\_n_ �_�_�_�_�_�_o�_ 7oIot���o�o� ��o�o�o(/!L/^/ p/�/{*o���� �����A�,�e� P�b����������Ώ ��+�=�(�a�L��� p������Oߟ񟠟�  �9�$�]�H���l�~� ����ۯƯ���#�No `oro�on��o�o�o�o Կ���8J\n g����vϯϚ����� ��	���-��Q�<�u� `�r߫ߖ��ߺ����� ��;�M�8�q�\�� ������z������%� �I�4�m�X���|��� ��������:�L�^� ��Z��������� ��$�6�H�S wb������ �//=/(/a/L/�/ p/�/�/�/�/�/?�/ '??K?]?H?�?��? �?f?�?�?�?O�?5O  OYODO}OhO�O�O�O �O�O�O&8J4_F_ ����_�_��_�_ "4-o�O*ocoNo �oro�o�o�o�o�o �o)M8q\� �������� 7�"�[�m��?����R� Ǐ���֏�!��E� 0�i�T���x������� �_$_V_ �2�l_~_�_�����R�$PL�ID_KNOW_�M  �T������SV ���U͠�U��
��.�ǟ�R�=�O�����mӣM_GRP 1�પ!`0u��T@ٰo�ҵ�
���Pз j��`���!�J�_� W�i�{ύϟϱ����ϰ����߱�MR���b��T��s�w� s� �ߠ޴߯߅��ߩ߻� ����A���'��� ������������ =���#���������`}������S��ST���1 1��U# �v��0�_ A . ��,>Pb��� �����3( iL^p������2*���<-/3/)/;/M/4f/x/�/�/A5�/�/�/�/6??(?:?7S?e?w?�?8�?�?�?�?�MAD  d�#`PARNU/M  w�%O�SCH?J ME
��G`A�Iͣ�EUPD�`OrE
a�OT_C�MP_��B@�P@'�˥TER_CHK'U��˪?R$_�6[RSl�¯��_M�OA@�_�U_�_RE__RES_G � �>�oo8o+o\oOo �oso�o�o�o�o�o�o �o�W �\�_% �Ue Baf�S� � ���S0����S R0��#��S�0>�]��b��S�0}������RV� 1�����rB@c�]��t�(@c�\����D@c�[�$���RTHR_INRl�DA��˥�d,�MASS9� �ZM�MN8�k�MO�N_QUEUE ����˦��x� *RDNPUbQN{�P[���END���_ڙEcXE�ڕ�@BE�|ʟ��OPTIOǗ��[��PROGRAoM %��%���ۏ�O��TASK_�IAD0�OCFG ����tO��ŠDA�TA���Ϋ@��27�>�P�b�t��� ,�����ɿۿ������#�5�G���INFO
Uӌ�������ϭ� ����������+�=� O�a�s߅ߗߩ߻��ߠ�����^�jč� �yġ?PDIT ��ίc���WER�FL
��
RGA�DJ �n�AЄ���?����@���I�ORITY{�QV�>��MPDSPH������Uz����OT�OEy�1�R� _(!AF4�E�P�]���!tcp|h���!ud�>�!icm��ݏn6�XY_ȡ�R�{�ۡ)� *+/ ۠�W: F�j����� �%7[Bz�*��PORT#��BC۠����_CARTREP
�|R� SKSTAz�^�ZSSAV���n��	2500H8�63���r�$!�*R����q�n��}/�/�'� URGE��B��rYWF� DO{�rUVWV��$�A��WRUP_DE?LAY �R��$�R_HOTk��%�O]?�$R_NOR�MALk�L?�?p6S�EMI?�?�?3AQ�SKIP!�n�l#x 	1/+O+  OROdOvO9Hn��O�G �O�O�O�O�O_�O_ D_V_h_._�_z_�_�_ �_�_�_
o�_.o@oRo ovodo�o�o�o�o�o �o�o*<Lr�`���n��$R�CVTM������pDCR!�L�ЈqB��C*�J�C$�>��$ >5?-;���04M¹�O���ǃ��������~��9On�Y�<�
6b<߈;�܍�>u.�?!<�&{� b�ˏݏ��8����� ,�>�P�b�t������� ��Ο���ݟ��:� %�7�p�S������ʯ ܯ� ��$�6�H�Z� l�~�������ƿ��� տ���2�D�'�h�z� ���ϰ���������
� �.�@�R�d�Oψߚ� �߾ߩ��������� <�N��r����� ��������&�8�#� \�G�����}������� ����S�4FXj |������� ��0T?x� u����'// ,/>/P/b/t/�/�/�/ �/�/�/�?�/(?? L?7?p?�?e?�?�?� �?�? OO$O6OHOZO lO~O�O�O�?�?�O�O �O�O __D_V_9_z_ �_�?�_�_�_�_�_
o o.o@oRodovo�X�q�GN_ATC 1��� A�T&FV0E/� �ATDP/6�/9/2/9�h�ATA�n,�AT%G1%B9�60/�+++��o,�aH,�qI�O_TYPE  ��u�sn_�oRE�FPOS1 1�>P{ x�o�Xh_�d_���� �K�6�o�
���.����R����{{2 1�P{���؏V�ԏz�<���q3 1��$��6�p��ٟ���S4 1�����˟����n���%�S5 1� <�N�`�����<���S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB�-�|f��S8 1������Y�������y�SMASK 1�P�  
9�G��XN	OM���a~߈Ӂq?MOTE  h�~t���_CFG ������рrPL_R�ANG�ћQ��PO�WER ��e���SM_DRY�PRG %i�%���J��TART ��
�X�UME_�PRO'�9��~t_�EXEC_ENB�  �e��GSP�D������c��TD�B���RM��MKT_!�T���`�OBOT_NAM/E i���i�OB_ORD_N_UM ?
�\q�H863 � �T���������bPC_TIME�OUT�� x�`S�232��1��k� LTEAC�H PENDAN �ǅ�}���`�Mainten�ance Con�s�R}�m
"{�dKCL/Cg��Z ��n� No Use}�	��*NPO��х����(CH�_L�������	��mMAVAI�L��{��ՙ�S�PACE1 2��| d��(>���&���p��M,8�?�ep/e T/�/�/�/�/�W// ,/>/�/b/�/v?�?Z? �/�?�9�e�a�=?? ,?>?�?b?�?vO�OZO@�?�O�O�Os�2�/O*O<O�O`O�O �_�_u_�_�_�_�_[3_#_5_G_Y_o}_ �_�o�o�o�o�o[4.o@oRodovo$ �o�o����"�	�7�[5K]o�� A����	�̏�?�&�T�[6h�z����� ��^�ԏ���&��;�\�C�q�[7������ ��͟{���"�C�� X�y�`���[8���� Ưدꯘ��0�?�`��#�uϖ�}ϫ�[G ;�i� �ϋ
G� ����$� 6�H�Z�l�~ߐ��8 ǀ������߈��d (���M�_�q��� ���������?��� 2�%�7�e�w������� �������������!� RE�W������ ����?Qw `�� @0���ߖrz	�V _�����
/L/ ^/|/2/d/�/�/�/�/ �/�/?�/�/�/*?l? ~?�?R?�?�?�?�?�? �?�?2O�?
��O�[_MODE  y�˝IS ���vO,*ϲ�O�-_��	M_v_#dCW�ORK_AD�M��A�%aR  ���ϰ�P{_�P_I�NTVAL�@�����JR_OPTIO�N�V �EBpV�AT_GRP 2ݭ���(y_Ho �e_vo�o �oYo�o�o�o�o�o *<�bOoNDpw ������	�� �?�Q�c�u�����/� ��ϏᏣ����)�;� ��_�q���������O� ɟ���՟7�I�[� m�/�������ǯٯ� ���!�3���C�i�{� ��O���ÿտ���� ��/�A�S�e�'ωϛ� ��oρ�������+� =���a�s߅�Gߕ߻� ���ߡ���'�9�K� ]��߁����y��� �������5�G�Y��E��$SCAN_T�IM�AYuew�R� �(�#((��<0.a�aPaP
Tq >��Q��o������OO2H/��:	d/JaR��WY��^����^R^	r  P���� �  �8�P�	�D��GYk}� �������Qp/@/R//<)P;�o\T���Qpg-�t��_DiKT��[  � lv%����� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OWW�# �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_olO ~Od+No`oro�o�o�o �o�o�o�o&8 J\n������u�  0�"0g�/ �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q�����$o�� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E����� Do��������ҿ��� ��,�>�P�b�tφ� �Ϫϼ���������w
�  58�J�\�n� �ߒߜկ��������� 	��-�?�Q�c�u��8���� ��- ����� �2�D�V�h� z�������������������& ���%	1234�5678�" 	��/� `r�������� (:L^p� ������ // $/6/H/Z/l/~/��/ �/�/�/�/�/? ?2? D?V?h?�/�?�?�?�? �?�?�?
OO.O@Oo? dOvO�O�O�O�O�O�O �O__*_YON_`_r_ �_�_�_�_�_�_�_o oC_8oJo\ono�o�o �o�o�o�o�oo" 4FXj|���������	��s�3�E�W�{�Cz�  Bp��   ���2���z�$�SCR_GRP �1�(�U8(ӿ\x^ �@  �	!�	 ׃��� "�$� ��-��+���R�w����D~�����#����O����M-10iAo 8909905 �Ŗ5 M61C �>4��Jׁ
� ���0�����#�1�	"�z�����h��¯Ҭ ��� c���O�8�J�� �����!�����ֿ.��B�y����������A��$�  @��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ�� ��������%��I�4� m��<�l߃ߕߧ���B���\����1� �U�@�R��v��� ��������;���*<=�
F���?�d��<�>7�����@��:��� B����ЗЙ���EL_�DEFAULT � �����B�MIPO�WERFL  ��$1 WFDO� $��ERV�ENT 1������"�pL!DUM_EIP���8��j!AF_�INE �=�!�FT���!���4 ��[!�RPC_MAI�N\>�J�nV�ISw=���!7TP�PU��	�d�?/!
PMON_PROXY@/��e./�/"Y/�f�z/�/!RDM_'SRV�/�	g�/#?G!R C?�h?�o?!
pM�/�i�^?�?!RLSY3NC�?8�8�?O�!ROS�.L�4�?SO"wO�#DOVO �O�O�O�O�O_�O1_ �OU__._@_�_d_v_ �_�_�_�_o�_?oo�coiICE_KL� ?%y (%�SVCPRG1@ho8��e���o�m3�oD�o�`4 �`5(D-�`6PU�`7x }�`���l9��{�d:?��a�o��a �oE��a�om��a�� �aB���aj叟a� ��a�5��a�]��a ����a3����a[�՟ �a�����a��%��aӏ M��a��u��a#����a K�ů�as���a��mo b�`�o�`8�}�w��� ����ɿ���ؿ��� 5�G�2�k�VϏ�zϳ� �����������1�� U�@�y�dߝ߯ߚ��� ��������?�*�Q� u�`��������� ���;�&�_�J��� n�����������sj_DEV y	��MC:�w�_OUT"�,REC �1�Z� d  �  	�    ��@�� ����A�����
 �PSD�#6 r��O*� �� �� `�� Q�Z�{� �� 9*�  +X- U� I- �- !- �� �X�YZ�PWSJ;4 ��?  (� � � ��R V��� E- � ��/e/�l�4�/��� X� (,/>/P/�/�/�"�"4� =�!� �
 ؀  ?"S1���'!�/���("- ��\?�?$=�=�? �?�?"OOFO4OjO|O ^O�O�O�O�O�O�O�O _ __T_B_x_f_�_ �_�_�_�_�_�_oo oPo>oto�oho�o�o �o�o�o�o(
L :\�p���w,����4�"� X�F�|���p�����֏ ď����0��@�f� T���x�����ҟ�Ɵ ���,��<�b�P��� h�z������ί�� (�:��^�L�n�p��� ����ܿ�п� �6� $�Z�H�jϐ�rϴϢ� ���������2�D�&� h�Vߌ�z߰ߞ����� ������
�@�.�d�R�x��ZjV 1�w� P����j 
�� ����
TYPEVF�ZN_CFG ��5d�~4�GRP 1�A�^c ,B� A�~ D;� B����  B4�RB21HELEL:�(
��?�<��<%RS'! ��H3lW�{ ������2�Vh�������%w����#!a�1�����7��2�0d����H�K 1���  �k/f/x/�/�/�/�/ �/�/�/??C?>?P?�b?�?�?�?�?��OM�M ����?��FTOV_ENB ����+�HOW_RE�G_UIO��IM/WAITB�JK�OUT;F��LIT�IM;E���OV�AL[OMC_UNI�TC�F+�MON_�ALIAS ?e~�9 ( he�� _&_8_J_\_B_�_ �_�_�_j_�_�_oo +o�_Ooaoso�o�oBo �o�o�o�o�o'9 K]n���� t���#�5��Y� k�}�����L�ŏ׏� �����1�C�U�g�� ��������ӟ~���	� �-�?��c�u����� ��V�ϯ������ ;�M�_�q�������� ˿ݿ����%�7�I� ��m�ϑϣϵ�`��� ����ߺ�3�E�W�i� {�&ߟ߱������ߒ� ��/�A�S���w�� ���X�������� ��=�O�a�s���0��� ����������'9 K]����b ���#�GY k}�:���� ��/1/C/U/ /f/ �/�/�/�/l/�/�/	? ?-?�/Q?c?u?�?�? D?�?�?�?�?O�?)O ;OMO_O
O�O�O�O�O �OvO�O__%_7_�C��$SMON_D�EFPRO ����`Q� *SYS�TEM*  d=�OURECALL� ?}`Y ( ��}
xyzra�te 61 >1�92.168.4��P46:6244} �W7956 �U��_�_�_n}�W=�]792�_�_aoso��od9copy �frs:orde�rfil.dat� virt:\tmpback\*o�<a�o�o�ol0�bm?db:*.*�o�o� �obt�c4x�d:\)�p;<aU���
� }5�ua ��7f�g�y����Z +�=�O�����o)o6580 ��ҏc� u����o�o56�ٟ� ��"��5�џb�t�䆯�6����emp>:�1652 W��t����.��*.d���Ʈϯ`�r�����1  +�=�O�����)� Ҳ��ҿc�uχϚ��� 5�ͧ�������"��� ̨��b�t߆ߙ���� K�V����������� >���h�z��ϱ�:� ������
�߸�A��� d�v�����.�;����� ������O�`r ����2����� �'��K�\n��� ��8�����# �G/j/|/����3/�E/W/�/�/�/ϱW5012?��/b?t?�? ��458�?�?�? "�?58�?bOtO�O����?���P8188  WO�O�O�O��O�I�O `_r_�_�/��;_M_�_ �_o?'?�T�_�_co uo�o�?�?5O�G�o�o �oO"O�o�I�ocu ���/�/RbU�� 
�/��Ta�h�z� ��o�o:����
� ��Aӏd�v�������$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1����?���%֟ ��&�	��\�?�f� ��u��������ϯ�� "��F�)�;�|�_��� ����ֿ��˿��� B�%�f�I�[Ϝ�Ϧ� �ϵ�������,��6� b�E߆�i�{߼ߟ��� ��������L�/�V� ��e��������� ���6��+�l�O�v� �������������� 2V9K�o� ������& R5vYk��� ��/��<//F/ r/U/�/y/�/�/�/�/ ?�/&?	??\???f? �?u?�?�?�?�?�?�? "OOFO)O;O|O_O�O �O�O�O�O�O_�O_ B_%_f_I_[_�__�_ �_�_�_�_�_,oo6o boEo�oio{o�o�o�o �o�o�oL/V �e������ ��6��+�l�O�v��������PARAM� ����� ��	��P�����OFT_K�B_CFG  �⃱���PIN_S_IM  ����C�U�g�����RVQSTP_DSB,��򂣟����SR ��/�� & � AR�����T�OP_ON_ER�ސ���PT�N /�@��A	�RINGo_PRM� ���VDT_GRP �1�ˉ�  	 ������������Я� ����*�Q�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߣߠ߲� ����������0�B� i�f�x�������� �����/�,�>�P�b� t��������������� (:L^p� ������  $6HZ�~�� �����/ /G/ D/V/h/z/�/�/�/�/ �/�/?
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8___\_��VP�RG_COUNT���@���REN�BU��UM�S��__�UPD 1�/�8  
s_�oo *oSoNo`oro�o�o�o �o�o�o�o+&8 Jsn����� ����"�K�F�X� j���������ۏ֏� ��#��0�B�k�f�x� ��������ҟ����� �C�>�P�b������� ��ӯί�����UYSDEBUG�P��P�)�d�YH�SP�_PASS�UB�?Z�LOG �V�U�S)�#��0�  ��Q)�
�MC:\��6���_MPC���U���Q�ñ8� �Q�SA/V �����ǲ�%�ηSV;�T�EM_TIME �1��[ (�P��T��ؿT1SV�GUNS�P�U'��U���ASK_OPTION�P�U�Q��Q��BCCFGg ��[u� n�X�G�`a�gZo��� �ߕ��߹������� :�%�^�p�[���� ������ �����6�!� Z�E�~�i���������%�������&8�� nY�}�?�� ԫ ��(L :p^����� ��/ /6/$/F/l/ Z/�/~/�/�/�/�/�/ �/�/2?8 F?X?v? �?�??�?�?�?�?�? O*O<O
O`ONO�OrO �O�O�O�O�O_�O&_ _J_8_n_\_~_�_�_ �_�_�_�_o�_ o"o 4ojoXo�oD?�o�o�o �o�oxo.TB x��j���� ����,�b�P��� t�����Ώ��ޏ�� (��L�:�p�^����� ��ʟ��o��6� H�Z�؟~�l������� د���ʯ ��D�2� h�V�x�z���¿��� Կ
���.��>�d�R� ��vϬϚ��Ͼ����� ��*��N��f�xߖ� �ߺ�8��������� 8�J�\�*��n��� ���������"��F� 4�j�X���|������� ������0@B T�x�d���� �>,Ntb ������/� (//8/:/L/�/p/�/ �/�/�/�/�/�/$?? H?6?l?Z?�?~?�?�? �?�?�?O�&O8OVO hOzO�?�O�O�O�O�O �O
__�O@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<o^o�oro �o�o�o�o�o�o  J8n$O��� ��X���4�"��X�B�v��$TBC�SG_GRP 2��B�� � �v� 
 ?�  ������׏ �������1��U�g��z���ƈ�d,� ���?v�	 H�C��d�>�����e�CL  B�p��Пܘ������\)��Y  A��ܟ$�B�g�B�Bl�i�X�ɼ���X��  D	J���r�����C����үܬ	���D�@v�=�W�j� }�H�Z���ſ���������v�	�V3.00��	�m61c�	*`X�P�u�g�p�>���2v�(:�� ��p���  O�����p�����z�JCFG� �B��� ,���������=��=�c�q�K� qߗ߂߻ߦ������ ��'��$�]�H��l� ������������#� �G�2�k�V���z��� �����������p *<N���l�� �����#5G Y}h���� v�b��>�// /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?d?R? t?v?�?�?�?�?�?O �?*OO:O`ONO�OrO �O�O��O�O�O_&_ _J_8_n_\_�_�_�_ �_�_�_�_�_�_oFo 4ojo|o�o�oZo�o�o �o�o�o�oB0f T�x����� ��,��P�>�`�b� t�����Ώ������ �&�L��Od�v���2� ����ȟʟܟ� �6� $�Z�l�~���N����� دƯ�� �2��B� h�V���z�����Կ¿ ����.��R�@�v� dϚψϪ��Ͼ����� ��<�*�L�N�`ߖ� �ߺߨ����ߚ��� ����\�J��n��� ��������"���2� X�F�|�j��������� ������.TB xf������ �>,bP� t�����/� (//8/:/L/�/�ߚ/ �/�/h/�/�/�/$?? H?6?l?Z?�?�?�?�? �?�?�?O�?ODOVO hO"O4O�O�O�O�O�O �O
_�O_@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<oro`o�o �o�o�o�o�o�o& �/>P�/��� ������4�F� X��(���|�����֏ ����Ə0��@�B� T���x�����ҟ���� ��,��P�>�t�b� ������������� �:�(�^�L�n����� ��2d�����̿� $�Z�H�~�lϢϐ��� �����Ϻ� ��0�2� D�zߌߞ߰�j����� �����
�,�.�@�v� d����������� ��<�*�`�N���r� ������������& J\�t��B ������F 4j|��^��p��/�  2 �6# 6&J/6"��$TBJOP_G�RP 2����  ?i�X,i#�p,� ��x�J� �6$�  �_< �� �6$� @2 �"	 ߐC�� �&b � Cق'�!�!>�c��
559>�0�+1�33=�{CL� fff?+0?�ffB� J1�%�Y?d7�.��/>��2\)?0�5����;��hC=Y� �  @� �!?B�  A�P?�?��3EC�  Dp�!�,�0*BOߦ?��3JB��
:���Bl�0��0�$�1��?O6!Aə�A�ДC�1D�G6��=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH��1ts�A@333@?1� C�� �@�_�_&_8_>��D��UV_0�LP�Q30<'{�zR� @�0�V �P!o3o�_<oRifoPo ^o�o�o�oRo�o�o�o �oM(�ol�pP~��p4�6&�q�5	V3.00��#m61c�$�*(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�N�aF���F�^�lF���F�:�
F�)F���3G�G���G��G,I�R�CH`�C��dTDU�?D���D��DE(�!/E\�E���E�h�E��ME��sF�`F+'\FD���F`=F}�'�F��F��[
F���F���M;S@;Q�*�|8�`rz@/&�
8�6&<��1�w��^$ESTPARS�  *({ _#HR���ABLE 1̒p+Z�6#|�Q� (� 1�|�|�|�5'T=!|�	|�
|�|�T˕6!|�|�|����RDI��z!�ʟܟ� ��$���O ������¯ԯ�����	S��x# V���˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �U-����ĜP�9�K� ]�o��-�?�Q�c�u����6�NUM  V�z!� > � Ȑ����_CFGG �����!@b �IMEBF_TT�����x#��a�VER腣b�w�a�R 1=�p+
 (3�6"	1 ��  6!���� ������ �9�$�:�H� Z�l�~����������� ����^$��_���@x�
b MI_CWHANm� x� k�DBGLV;0o��x�a!n ETHER_AD ?�� �y�$"�\&n oROUT��!p*�!*�SNM�ASK�x#�255.h�fx^$�OOLOFS_D�I��[ՠ	ORQCTRL �p+ ;/���/+/=/O/ a/s/�/�/�/�/�/���/�/�/!?��PE_�DETAI��P�ON_SVOFF��33P_MON ��H�v�2-9ST�RTCHK ����42VTCOMPATa8�24:0�FPROG %�%CA)&O�3?ISPLAY��L:_INST_MPe GL7YDUS���?�2LCK�LPKQ?UICKMEt �O��2SCRE�@>�
tps��2 �A�@�I��@_Y����9�	SR_GRP� 1�� ���\�l_zZg_�_ �_�_�_�_�^�^�o j�Q'ODo/ohoSe� �oo�o�o�o�o�o�o !WE{i�������	1?234567���!���X�E1�V[
� �}ipnl�/a�gen.htmno��������ȏ~��Panel _setup̌}�?���0�B�T�f�  ��񏞟��ԟ��� o����@�R�d�v��� ���#�Я����� *���ϯůr������� ��̿C��g��&�8� J�\�n�����϶��� ������uϣϙ�F�X� j�|ߎߠ����;��߀����0�B��*NU�ALRMb@G ?�� [���� �������� ��%�C��I�z�m�������v�S�EV  �����t�ECFG �Ձ=]/BaA$ �  B�/D
  ��/C�Wi{�� ����� PRց; �To\�o�I�6?K0(% ����0����� //;/&/L/q/\/�/0�/�/l�D �Q��/I_�@HIST� 1ׁ9  �(  ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1?pv?�?�?�?�� >?P=962c?�?
OO0.O�?�?�136�?|O �O�O�OAOSOeO�O_ _0_�HM___q_�_�_ �_�_H_�_�_oo%o 7o�_[omoo�o�o�o Do�o�o�o!3E ��a81�ou�� ����o���)� ;�M��q��������� ˏZ�l���%�7�I� [���������ǟٟ h����!�3�E�W�� ��������ïկ�v� ��/�A�S�e�Pb ������ѿ������ +�=�O�a�s�ϗϩ� ��������ߒ�'�9� K�]�o߁�ߥ߷��� �����ߎ�#�5�G�Y� k�}���������� �����1�C�U�g�y� ��v�����������	 �?Qcu�� (����) �M_q���6 ���//%/�I/ [/m//�/�/�/D/�/ �/�/?!?3?�/W?i? {?�?�?�?�����?�? OO/OAOD?eOwO�O �O�O�ONO`O�O__ +_=_O_�Os_�_�_�_ �_�_\_�_oo'o9o Ko�_�_�o�o�o�o�o �ojo�o#5GY �o}������?���$UI_PA�NEDATA 1�������  	�}��0�B�T�f�x��� )����mt�ۏ��� �#�5���Y�@�}��� v�����ן��������1��U�g�N������ �1��Ïȯگ ����"�u�F���X� |�������Ŀֿ=��� ���0�T�;�x�_� �Ϯϕ��Ϲ������,ߟ�M��j�o߁� �ߥ߷������`�� #�5�G�Y�k��ߏ�� ������������� C�*�g�y�`������� ��F�X�	-?Q c����߫��� �~;"_F ��|����� /�7/I/0/m/���� �/�/�/�/�/�/P/!? 3?�W?i?{?�?�?�? ?�?�?�?O�?/OO SOeOLO�OpO�O�O�O �O�O_z/�/J?O_a_ s_�_�_�_�O�_@?�_ oo'o9oKo�_oo�o ho�o�o�o�o�o�o�o #
GY@}d� �&_8_����1� C��g��_�������� ӏ���^���?�&� c�u�\�������ϟ�� �ڟ�)��M��� ��������˯ݯ0�� ���7�I�[�m���� ������ٿ�ҿ��� 3�E�,�i�Pύϟφ�`�Ϫ���Z�l�}���@1�C�U�g�yߋ�)� ��#������� ��$� 6��Z�A�~�e�w�� ����������2���V�h�O�����v�p���$UI_PANELINK 1�v��  ��  ��}1�234567890����	-?G  ���o����� a��#5G�	�����p&���  R�����Z ��$/6/H/Z/l/~/ /�/�/�/�/�/�/�/ 
?2?D?V?h?z??$? �?�?�?�?�?
O�?.O @OROdOvO�O O�O�O �O�O�O_�O�O<_N_``_r_�_�_�0,�� �_�X�_�_�_ o2oo VohoKo�ooo�o�o�o �o�o�o��,> r}�������� ����/�A�S�e� w��������я��� tv�z����=�O� a�s�������0S��ӟ ���	��-���Q�c� u�������:�ϯ�� ��)���M�_�q��� ������H�ݿ��� %�7�ƿ[�m�ϑϣ� ��D��������!�3� Eߴ_i�{�
�߂��� �߸������/��S� e�H���~��R~'� '�a��:�L�^�p� ��������������  ��6HZl~� ��#�5���  2D��hz��� ��c�
//./@/ R/�v/�/�/�/�/�/ _/�/??*?<?N?`? �/�?�?�?�?�?�?m? OO&O8OJO\O�?�O �O�O�O�O�O�O[�_ ��4_F_)_j_|___�_ �_�_�_�_�_o�_0o oTofo��o��o� �o�o�o,>1 bt����K� ���(�:���� {O������ʏ܏�uO �$�6�H�Z�l����� ����Ɵ؟����� � 2�D�V�h�z�	����� ¯ԯ������.�@� R�d�v��������п ���ϕ�*�<�N�`� rτ��O�Ϻ�Io���� �����8�J�-�n߀� cߤ߇����߽���� o1�oX��o|��� �����������0� B�T�f���������� ����S�e�w�,>P bt��'��� ��:L^p ��#���� / /$/�H/Z/l/~/�/ �/1/�/�/�/�/? ? �/D?V?h?z?�?�?�? ??�?�?�?
OO.O�� ROdO�߈OkO�O�O�O �O�O�O_�O<_N_1_ r_�_g_�_7OM��m�$UI_QU�ICKMEN  }��_�AobRESTOR�E 1�  �|��Rto�o�im�o�o�o �o�o:L^p �%������o ����Z�l�~��� ��E�Ə؏���� � ÏD�V�h�z���7��� ����/���
��.�@� �d�v�������O�Я �����ßͯ7�I� ��m�������̿޿�� ��&�8�J��nπ� �Ϥ϶�a�������Y� "�4�F�X�j�ߎߠ� �������ߋ���0�xB�T�gSCRE`�?#mu1�sco`u2��3���4��5��6��7��8��bUSER�q�v��Tp���ksT����4��5��6���7��8��`NDO_CFG �#k�  n` `PD�ATE ����NonebS�EUFRAME � �TA�n�RTOL_ABRTy��l��ENB����G�RP 1�ci/a?Cz  A�����Q�� $6HRd��`U�����?MSK  ������Nv�%�U�%����bVISCA�ND_MAX��I��FAILO_IMG� �PݗP�#��IMREG�NUM�
,[S�IZ�n`�A��,VONTMOU4��@���2���a��a�����FR:\� � M�C:\�\LOGn�B@F� !��'/!+/O/�Uz �MCV�8#7UD1r&EX{+�S��PPO64_t��0'fn6PO��LIb�*r�#V���,f@�'޻/� =	�(SZ�V�.����'WA�I�/STAT ����P@/�?�?��:$�?�?��2D�WP  ��P� G@+b=���� H�O_JMP�ERR 1�#k
�  �2345678901dF�ψO {O�O�O�O�O�O_�O *__N_A_S_�_
� MLOWc>
 �g_TI�=�'�MPHASE  ���F��PSH�IFT�1 9�]@<�\�Do�U#o Io�oYoko�o�o�o�o �o�o�o6lC U�y������ ��	�V�-�e2�����	VSFT1��2	VM�� S�5�1G� ���%�A�  B8̀�̀�@ pكӁ˂�у��z�ME@�?�q{��!c>&%�a�M1��k�0�{ ��$`0TDINEND��\�O� �z�����S��w��P�{��ϜRELE�Q��Y���\�_AC�TIV��:�R�A ��e���e�:��RD� ���YBO�X �9�د�6���02����190.0.�8�3��254t��QF�	 ��X�j��1�r�obot���   p�૿�5pc��̿������7�����-�f�ZA+BC�����,]@U� �2ʿ�eϢωϛϭ� ������ ���V�=� z�a�s߰�E�Z��1�Ѧ