��   D�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���C�ELLSET_T�   w$�GI_STYSEL_P 7_T  7ISAO:iRibDi�TRA�R��I_INI; ���t�bU9ARTaRSRPNS1Q�2345*678Q
�TROBQACKSNO��) �7�E�S�a@�o�z2 U3 4 5 6 �7 8awn&GINm'D�&��)%� �)4%��)P%��)l%3SN�{(OU��!|7� OPTNA�73�73.:B<;}a6�.:C<;CK;CaI?_DECSNA�38R�3�TRY1���4��4�PTHC�N�8D�D�INCYC@HG�KD�?TASKOK�{D �{D�7:�E�U:�C h6�E�J�6�C�6U�J��6O�;0U��:IAT�L0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T��T�@REQ�d��drG�:Mf�GJO_HFAUL�Xd�dvgALE� �g�c�g�cvgE� �H�dvg�NDBR�H�dgR�GAB�Xtb  �CLMLIy@�   $�TYPESIND�EXS�$$CL�ASS  ����lq��;pupapV?IRTUALi{q�'61ION  ~����q��t+ UP0 �u�q�Style �Select 	�  ��r�uReq. /Echo���yAck����sInitiat(�p�r�s�t@�O��a�p���	��  U�����������q�������q���sOption� bit A���B����C�Dewcis�cod;���zTryout �mL��Path �segJ�ntin5.�II�yc:��Task OK���!�Manual _opt.r�pA�ԖBޟԖC�� d�ecsn ِ�R�obot int�erlo�"�>� Oisol3��C���i/�"�z�ment���z�ِ����_�s�tatus�	M�H Fault:<��ߧAler���%��p@r 1�z �L��[�m�+�; L�E_COMNT �?�y�    ��䆳�Ŀֿ���� �0�B�T�g�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼�@�����������U�������   ��E�NAB  �� �u�����������MENU>�y��NAME ?%��(%$*4���D��p 2�k�V���z������� ������1U@ Rdv����� ��*<u` �������� /;/&/_/J/f/n/�/ �/�/�/�/?�/%?? "?4?F?X?j?�?�?�? �?�?�?�?�=