��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ��'�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�
  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"�SBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� �21� _A.	 \vrVE�1$F��A{$O��D�B~�CTMP1_F�E2�G1_�3�B�2��XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�0@� �zsa�!ip;G0� � 
$WARNM�0f�!,P� ܁s�pNST� CO�RN�"a1FLTR^�uTRAT� T�p; H0ACCa1�p��{�ORI
`l"S={RT0_S�BְqHG,I1 E[ Tp�"3I9�CTY�D,P*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7���8��94�qO�$ <� $6x8K3 1w`O_M�@�C_ t � E#f6NGP�ABA�  �c��ZQ���`���@n!r��� ��P�0��,��x�p�PzP�b26����"J�_)R��BC�J��3�JVP��tBS��}�Aw��"�tP_*0O�FSzR @� RcO_K8���aIT�3���NOM_�0�1�ĥ3�p��T Ԑ� $���AxP��K}EX�� �0g0I01��p��
$TFa��C$7MD3��TO�3�0yU� �� �)Hw2�C1|�EΡg0wE{vF�vF�40�CPp@�a2 
P�$A`PU�3Nc)#�dR*�AX�!�sDETAI�3BU�FV��p@1 |X�p۶�pPIdT� +PP[�MZ�Mg�Ͱ�j�F[�SIMQS�I�"0��A.����PNkx Tp|zM�x�P�B�FACTrbHPEW7�P1Ӡ��v��MCd� �$*1JB�p<�*1DECHښ�H���b�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF4��� &k�Bv�u�cu��a E�� !2��+�MQ��EчSIZ�3����T��P�����aRSINF�����kq��������LX������F�CRCMu�3CC lpG��p���O}���b��1�������2�V�D
xIC��C���r����0P��{� EV �zUF_��F�pNB
0�?������A�! �r�Rx���� V�lp�2��aR�t�,��g�RTx �#�5�5"2��uARt���`CX�$LG�p��B�1 `s�P�t�a!A�0{�У+0R���tME�`!BupCr3RA 3tAZ�л4�pc�OT�FC�b�`��`FNp���1��ADI+�a%��b��{��p$�pSp�c�`S0�P��a,QMP6�`IY�3��M'�pU���aU  $>�TITO1�S�S�!���$�"0�DBPXW�O��!��$S1K��2�DB��"�"@�PR8� �
� ���# l>�q1$��$��
+�L9$?(�V�)%@?R4C&_?R4gENE��'~?�(�� RE�pY2(�H �OS��#$L�3$$3R�h�;3�MVOk_D@!V�ROScrr�w�S����CRIGGER�2FPA�S��7�ET�URN0B�cMR_���TUː[��0EkWM%���GN>`���RLA���Eݡ<�P�&$P�t�'�@4a��C�DϣV��DXQ��4�1��MVG�O_AWAYRM�O#�aw!�D�CS_)  `IS#� �� �s 3S�AQ汯 4Rx�@ZSW�AQ�p�@1UW��NcTNTV)�5RV
a����|c�éWƃ��J�B��x0��SAFE�ۥ�V_SV�bEX�CLUU�;��ONL��cYg�~az��OT�a{�HI_V�? ��R, M�_ �*�0� ��_z�2�� 
CdSGO  +�rƐm@�A�c~b���w@��V�i�b�fANNUNx0�$�dKIDY�UABc�@@Sp�i�a+ �j�f1�!��pOGIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�� 6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6Cq�!MS�WU. 8��KE3YI��5�TM�1�s�qoA�vINޱE��!�, / D��HOST�P!4���<����<�°<��p<�EMp'���Z�� SBL� �UL��0  p�	����DT�0~1 � $��>9USAMPLо� /���決�$ I@�>� $SUBӄ���w0QS�����#��SAV�����c�S< 9�,`�fP$�0E!� �YN_B�#2 0&��DI�d�pO|�m�v�#$F�R_IC�� �ENC2_9Sd3  ��< 3�9���� cgp�����4�"��2�A��ޖ5���`���@Q@K&D-!�a�AVER�q����gDSP
���PC_��q��"�|�ܣ�VA�LU3�HE�(�M��IP)���OPPm �TH�*��"��S" T�/�Fb�;�d����d D�q�1�6 H(rLL_DUǀ�a�@��k���֠OT�"U�/����q@@NOAUT5O70�$}�x�~�@s��|�C ����C� 2 �z�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|¶�'����9 A<���z�ΓKI��0��H硵FEq@{@�: ,��&a?3 P_P?��>�J����E�@��r��RP��;fp$T�P�$VARI�����,�UP2Q`< W�߃TD��g���П`��������BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P�"u�Fl@``>Gt ;��6����ST����T��M ����0	��i���F� ��������kRt ����FORCEUP�b^܂FLUS
pH(�N��� ��6bD_CM�@E�7N� (��v�P��REM� F a��@j���
�K�	N���EFF�/���@IN�QO�V��OVA�	TgROV DT)��DTMX:e � P:/��Pq�vXpCLN _�p��@d ��	_|��_T: T�|�&PA�QDI���1��0�&Y0RQm�_+qH�2��M���CL�d#��RIV{�ϓN"EAmR/�IO�PCPd��BR��CM�@�N 1b 3GCLF��!DY�(�q6�#5T�DG���8� �%%�FSS� )��? P(q1�1��`_1"811�E�C13D;5D6�GSRA���@�����PW�ON2EBUG�S�2�C`g�ϐ_E A ���@a �TER�M�5B�5���OR�Iw�0C�5/���SM_-`���0D\�5p��TA�9E�5�E  �UP��F�� -QϒA��P�3�@B$SEG�GJ� EL�UUSE.PNFI��pBx���1@��4>DC$UF�P��$���Q�@"C���G�0T������SNSTj�PATxۡg��APTHJ�A�E*�Z%qB\`F�{E��F�q�pARxPY�aSHFT͢qA�AX_SHOR$�>��6% @$GqPE���GOVR���aZPI@P�@$U?r *aAYLO���j�I�"��A8ؠ��ؠERV��Q i�[Y)��G�@R��i�e��i�R�!P�uA�SYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C��%UP���P���WORڒ@M��k0SM5T��G��GR��3�aPA�@��p5�'�_H � j�A�'TOCjA7pP]Pp$OPd�O��C��%�p�O!��R%E.pR�C�AO�?��Be5pR�EruIx|'QG�e$PWR) 3IMdu�RR_$s��\5��B Iz2H8��=�_ADDRH�H_LENG�B�q�qT:�x�R��So�J.�SS��SK�����0� ��-�SE*��ھrSN�MN1K�	�j�5�@r�֣O�L��\�WpW�Q�>pACRO�p���@H �����Q� ��OUPW3�b_>�I��!q�a1��������|�� ������-���:���ViIOX2S=�D��e��]���L $x��p�!_OFF[r�_�PRM_�^�aTTP_�H��wM (�pOBJ�"l�pG�$H�LE�C���ٰN � \9�*�AB_�T��b
�S�`�S��LV���KRW"duHITC�OU?BGi�LO�q����d� Fp�k�GpSS� ���HQWh�wA��O.��`�INCPUX2VISIO��!��¢.��á<�á-� �IO�LN)�P 87�R�'�[p$SL�b�d PUT_��$�dp�Pz �� F�_AS2Q/�$ALD���D�aQT U�0�]P�A������PH�YG灱Z���5�UO� 3R `F���H�@Yq�Yx�ɱvpP�S�dp���x��ٶBP��UJ��S����NEΊWJOG�G �DI�S��r�KĠ��3T� |��AV��`_�C�TR!S^�FLAG�f2 �LG�dU� �n�:��3LG_SIZ��ň�X��=���FD��I�� ��Z �ǳ��0�Ʋ�@s ��-ֈ�-�=�-���-�x�0-�ISCH_��Dq��N?���V���EE!2�C��n�Uȡ����`L�Ӕ�DAU��EA��Ġt�����GHr��I�BO}O)�WL ?`��� ITV���0\�R;EC�SCRf 0��a�D^�����MARG��`!P�)�T�/ty�$?I�S�H�WW�I�ܩ�T�JGM��MN�CH��I�FNKEuY��K��PRG���UF��P��FWDv��HL�STP���V��@�����RS"S�H�` �Q�C�T1� ZbT�R ���U����@��|R��t�i���G��8PPO��6�F�1�Mޘ�FOCU��RG�EXP�TUI��IЈ�c��n��n ����ePf���!p6�ePr7�N���CANAI��jB��VAIL��C�Lt!;eDCS_H!I�4�.��O�|!"�S Sn�}��_BUFF1�XY��PT�$ �� �v��f�L6q
1YY��P ������pOS1�2�3���� 0Z �  ��aiE�*���IDX�dP�RhrO��+��A&ST��R���Yz�<! Y$EK&CK+���Z&pm&��E�1[ L�� o�0��]PL�6pwq�t�^����w��7�_ \ �`��瀰�7�t�#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3�1DM�R7��LDR5<4R5ORG.���e2(` ���V�8.��T<�4�d^ �q�<4��-4R5�S�`T00m��0D>FRCLMC!D�?0�?3I@��MIC��dg_ d���RQm�=q�DSTB	� c �Fg�HAX;b� �H�LEXCE�SZr/oEMup�a`� �B;d�rB`��`5a��F_A�J���$[�O�H0K�db q\��ӂS�$MB���LIБ}SREQU�IR�R>q�\Á�XD�EBU��oAL� MP�c�ba��P؃ӂ!B�oAND���`�`d0�҆�c�cDC1��IN�����`@�(h?�Nz�@q��o��UP�ST8� e�rL�OC�RI�p�E�X�fA�p��AoAOwDAQP�f X��3ON��[rMF���� �f)�"I��%�e��T�v�!FX�@IGG� g �q��"E��0��#���$R�a% ;#7y��Gx��VvCPi�ODATAw�pE:��y��RFЭ�NVh �t $MD�qI�ё)�v+�tń�tH��`�P�u�|��sAN�SW}��t�?�uD��)�b�	@Ði -�@CU��V�T0�eRR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2N�RIN��v�<��'NTE���kE����,��b����_Nl@��ڂ��kDׄRm�7DIViFDH�@ـ:n�$V��'cv!$��$Z������~�[��o�H �$BEL�Tb��!ACCEL�+��ҡ��IRC��t����T/!���$PS�@#2L� q�Ɣ83������� ��PATH��������3̒Vp�A_�Q�.��4�B�Cᐈ�_M=Gh�$DDQ���G�$FWh��p���m�����b�DE��P�PABNԗROTSPEED����00�J�Я8��@����$USE_��P���s�SY��c�A �kqYNu@Ag��OsFF�q�MOUN�3NGg�K�OL�H�INC*��a��q��Bxj�L@�BENCS���q�Bđ���D��IN�#"I̒��4�\BݠV�EO�w�Ͳ23_UyPE�߳LOWLA���00����D��@�BwP��� �1RCʀ�ƶMOSIV�JRM�O���@GPERC7H  �OV�� ^��i�<!�ZD<!�c@��d@�P��V1�#P͑��L���EW�ĆĸUP������T�RKr�"AYLOA'a�� Q-�(�<�1�8�`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H�����b�DUM2(�S_�BCKLSH_C (���>�=�q�#�U��������2�t�]ACLA�LvŲ�1n�P�C�HK00'%SD�RT�Y4�k��y�1�q_�6#2�_UM$Pj�C�w�_�SCL��ƠLMT_J1_LO�"�@���q��E������๕�幘SPC`��7������PCo�B��H� �PU�m�C/@��"XT_�c�CN_b��N��e���SFu���V�&#����9�(�d��=�C�u�SH6# ��c����1�Ѩ�o�0�0͑
��_�PAt�h�_Ps�W�_10��4֠R�01D�VG�J� L��@J�OGW���ToORQU��ON*ɀMٙ�sRHљ��_	W��-�_=��C��TI��I�I�II�	F�`�JLA.�1[��VC��0�D�BO1�U�@i�B\JRK�U��	@DBL_�SMd�BM%`_D9LC�BGRV��0C��I��H_� �*COS+\�(LN�7+X>$C�9)�I�9)u*c,)�Z2 HƺMY@!�( "�TH&-�)THET=0�NK23I��"l=�A CB6CB=�C�A�B(261C�61�6SBC�T25GT	S QơC��aS$�" �4c#�7r#$DUD�EX�1s�t��B�6䆱�AQ|r�f$NE�DpIB U�\B5��	$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2��&�C�J�&!�VAHV�6H3�YLVhJVuKV��KV�KV�KV�KV�IHAHZF`RXM��wX�uKH�KH�KH�KH��KH�IO2LOAHOT�YWNOhJOuKO�KUO�KO�KO�KO�&�F�2#1ic%�d4GS�PBALANCE�_�!�cLEk0H_�%SP��T&�bc&�b>r&PFULC�hr��grr%Ċ1ky�U�TO_?�jT1T2Cy��2N&�v�ϰ ctw�g�p�0Ӓ~����T��O���� IN�SEGv�!�REV8�v!���DIF�鉳1l�w�1m
�OaB�q
����MIϰ�1��LCHWAR̭���AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|�n��ROBR�CR(����N�'�MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD�0�ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDX�Р  ��MOR^��t $-�U�� )��r�B���(�����Gؒu � $SIMULT ��~�x�� ���OBJE�`> �ADJUS>�1�OAY_Ik��D_�����C�_FIF�=�T� ��Ұ��{���p� �����p�@��DN�FRI��ӥT�ՓRO� ��E����͐OPWO�ŀv�0��SYSBU<�@ʐ$SOP�����#�U"��pPRUYN�I�PA�DH��D����_OU��=��qn�$}�IMKAG��ˀ�0P�q3IM����IN�q�~��RGOVRDȡ:���|�P~���Р�0�L_6p���i��R)B���0��M���SEDѐF� ��N`�M*����̰SL��`ŀw x $�OVSL�vSDI��DEXm�g�e�9Hw�����V� ~�N����w����Ûǖȳ�M��@��q<��� �x HˁE�F�AT+US���C�0à�ǒ��BTM����I
f���4����(�ŀy DˀEz�g���PE�r�����
���EXE��V��E�Y�8$Ժ ŀz @ˁ��3UP{�h�$�p��XN���9�H�� �PG"�{ h? $SUB��c��@_��01\�MPW�AI��P����LO��<�F�p�$R�CVFAIL_C�f�BWD"�F����DEFSPup | Lˀ`�D�� U�UNI��S�b��R`���_L�pAP��̐���ā}���� B�~���|��`ҲNN�`KET��y���P� $�~���0SIZE] ଠ{����S<�OR��FORMAT/p � F��ᖫrEMR��y�UqX���@�PLI7�~ā  $�P_SWI��Ş�_PL7�AL_ S�ސR�A��B��(0C��Df�$E�h����C_=�U�� � � ���~�J3�0�����TIA4��5��6��MOM������h �B�AD��*��* PU70NARW��W R������ A$PI�6���	�� )�4l�}69��Q����c�SPEED�PG q�7�D�>D�� ��>tMt[��SAM�`痰>��MOV���$��p �5��5�D�1�$2�������{�Hip�IN?,{� F(b+=$�H*�(_$�+�+GAMM�f�1{�$GET��ĐH��D����
^pLIB�R�ѝI��$HIB��_��Ȑ*B6E��b*8A$>G086LW= e6\<G9�686��R���ٰV��$PGDCK�Q�H�_����;"��z�.%�7��4*�9� �$IM_SRO��D�s"���H�"�LE��O�0\H��6@�qR� �ŀ�P�q?UR_SCR�ӚA�Z��S_SAVEc_D�E��NO��CgA�Ҷ��@�$��� �I��	�I� %Z[�  ��RX" ��m���" �q�'"�8�H ӱt�W�UpS���Q�M��O㵐.'}q�� Cg���@ʣ����S��M�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PL�M���	� 0h�H�{�X��O��z�Z�eT�M����� pS��C ��O__0_B_�a��_%�� |S����@ 	�v��v �@���w�v��EM��%O�fr�B��ː��ftP���PM��QU� ŉU�Q��Af�QT�H=�HOL��QH�YS�ES�,�U�E��B��O#��  -�P0�|�gAQ����ʠu���O��ŀ��ɂv�-�A;ӝROG��a2D�E�Â�v�_�ĀZ�INFOB&��+����bȜ�OI킍 ((@SLEQ/�#�������o���S`c0O��0�01EZ0N9Ue�_�AUT�Ab�COPY��Ѓ�{�
�@M��N�����1�4P�
� ��RGI��͏��X_�Pl�$P�����`�W��P���j@�G���EXT/_CYCtb����p����h�_NAƹ!$�\�<�RO��`]�� � m��POR�ㅣ�.��SRVt�)����DI �T_l���Ѥ@{�ۧ��ۧ �ۧ5٩�6٩7٩8����S��B쐒��$�F6���PL�A�A^�TAR��@E `�Z�����<��d� ,�(@FLq`h��@YN�L���M�C���P�WRЍ�쐔e�D�ELAѰ�Y�pA�D#q�RQSKIPN�� ĕ�x�O�`�NT!� ��P_ x���ǚ@�b�p1� 1�1Ǹ�?� �?���>��>�&�>�3�>�9��J2R;쐖� 4��EX� TQ ����ށ�Q���[�K�Fд�'�RDCNIf� �U`�X}�R�#%M!*�0�)��$�RGEAR_0I9O�TJBFLG�i&gpERa��TC݃��|����2TH2N���� 1�b��G:q T�0 ���ЉM���`Ib��v�R�EF�1�� l<�h��ENAB��lcTPE?@���!(� ������Q�#�~�+2P H�W���2�Қ��@�"�4�F�X�j�3���{��������j�4�Ҝ��
��.�@�R�j�5�ҝu�����P������j�6�Ҟ���(:L�P��7�ҟo�����
j�8�Ҡ��"x4Fj�SMSK������a��E�A���MOTE������@ "1��Q�IO�5"%I��P�����POWi@쐣  �����X�gpi������Y"$DSB_SIGN4A�Qi�̰�C�ШP�ARS23�2%�Sb�iDEVICEUS#�R�R�PARIT�!O�PBIT�Q��O?WCONTR��QXⱓ�RCU� M�S�UXTASK�3NxB��0�$TATU�PK��S@@쐦F��6�_�PC}�$F�REEFROMS8]p�ai�GETN@S��UPDl�ARBA"S�P%0���� !>m$USA���a8z9�L�ERI�0f�&�pRY�5~"_�@f�qP�1�!�6WRK�D9�F9ХFR�IEND�Q4bUFx��&�A@TOOLHF�MY5�$LEN�GTH_VT��FCIR�pqC�@�E� �IUFIN�R����RGI�1�AITI:�xGX��I�FG2�7G1a����3��B�GPRR�DA��Oa_� o0e�I1RER�0đ�3&���TC���AQJV �G|�.2���F��1�!d�9Z�8 +5K�+5��E�y�L0�4��X �0m�L
N�T�3Hz��89��%��4�3G��W�0�W�RdD�Z��Tܳ���K�a3d��$cV �2���1��I1TH�02K2sk3K3Jci�aI�i�a�0L��SL��R$Vؠ�B�V�EVk�]V*R��� �,6Lc���9V2�F{/P:B��PS_�E���$rr�C�ѳ3$A0��wPR���v�U�cSk�� {��$�1���� 0���VX`�!�tX`��0P��ꁂ
�5SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V����S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD�<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C���:c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQ�pfC�ѷ =	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�q� �X��ȑ� �o .A$�1$�c1 Ē���7� x~�EG�0ݓ��q!AR����0�9>B�%��AXE.��ROB��W�A4�_�-֣SY���!6���&S�'WR���-1���STR��5�:9�E�� 	5B��=QB90�@6�������OT�0o 	$�ARY8�w20�Ԛ�	%�FI��;�$LINK�H��1%�a_63�5�q�2XYZ"��;�qH�3@��1�2�8{0	B�{D��� CFI��6G��
�{�_J��6��3NaOP_O4Y;5�FQTBmA"�BC
�z�DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ �@�5<:7�� W1�?0K�Mc��68Cb�vrb�4�ORQ��X�>8�#op ������wq�Uf����N�TOVE�Q��M;����E#�UK#�UQ"�VW �ZQ�W���Tυ� ;� ����QH�!`�ҽ��U��Q�WkeK#kecXE)R��	GE	0��S�dAWaǢ:D���0�7!�!AX�rB !{q��1uy-! y�pz�@z�@z6P z\Pz� z1v� y�y�+y�;y� Ky�[y�ky�{y�x�y�q�yDEBU��$����L�!º2WG`  AB!�,�r�SV���� 
w� ��m���w����1���1 ���A���A��6Q��\Q����!�m@��2CLAB3B�U������S  V ER|���� � $�@ڳ Aؑ!p�PO���Z�q0w�^�_M�RAȑ� d r T�-�ERR�L�TYz�B�I�qV3@�cΑTOQ�dB:`L� �d2�]��X�C[! � p��`T}0i��_V1��r�a'�4�2-�2<����@P�����F�G$W��g��V_!�l�$�P����c蝢q"�	V FZN�_CFG_!� 4 ��?º�|�ų����@��ȲW ���\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(�����!�s�Q�g�P{R	��SHELLĥ�� 56�B_BAS!�RSR��ԣo E�#S��[��1r�U%��2ݺ3ݺ4ݺU5ݺ6ݺ7ݺ8ݷ��ROOI䰝0�03NLK!�CAB� n��ACK��IN��T:�1�@�@ z�m�7_PU!�CO� ��OU��P� Ҧ) ���޶��TPFWD�_KARӑ�@��R�E~��P��(��Q�UE�����P
��C�STOPI_AL �����0&���㰑�0GSEMl�b�|�M��6d�TY|�SOK�}�DI�����(����_TM\�MANR�Q�ֿ0E+�|�$�KEYSWITCaH&	���HE
�OBEAT����E� �LEҒ���U��F�O�����O_HOuM�O�REF�P�PRz��!&0��Cr+�OA�ECO��xB�rIOCM�D�8׵�\���8�` �# D�1����U��&��MH�»P�CFOR�C��� ��O}M�  � @V�T�|�U,3P� 1-��`� 3-�4��N�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��C@�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fi]7s�'� P��UPD��  ���|�԰��YSL}OǢ� � z� �и���o�E��`>�^t��АALUץ�����CU���wFOqID�_L�ӿuHI�zI~�$FILE_�Ì�t��$`�,pMsS�A��� h���E_BLCK�#�C>,�D_CPU<�{� <�o����tJr���R ��
PWl O� ��LA���S��������RUN F�Ɂ��Ɂ����F�����ꁬ� �TBC�u�C� �X ;-$�LENi���v������I��G�L�OW_AXI�F)1��t2X�M����hD�
 ��I�� ���}�TOR����Dh��� L=��⇒�8s���#�_MA`�8ޕ��ޑTCV����T���&��ݡ�����J�����J����MDo���J�Ǜ ����
���2��� v���l��F�JK��VKi�hΡv�Ρ3��J0㤶ңJJڣJJ�A�ALң�ڣ��42�5z�&�N1-�9�(��␅�L~�_Vj�������� ` �GROU�pD��}B�NFLIC�����REQUIREa�EBUA��p����2¯�����c�ޞ� \��APKPR��C���
�;EN�CLOe�ɇS_M v�,ɣ�
����� ��M�C�&���g�_MG�q�C� �{�9����|�BRKz�NOL��|ĉ R��_LI�|��Ǫ�k�J����P 
���ڣ�����&���D/���6��6��8���r���� ���8�%�W�2�e�PATHa�z�p�z�=�hvӥ�ϰ�x�CN=��CA�����p�INF�UC��bq��CO�UM��YZ������q�E%���2������P�AYLOA��J2=L3pR_AN��<�L��F�B�6�R�{�R_F2LSHR��|�LOG��р��ӎ�>��ACRL_u��Ր����.���H�p��$H{���FLEX�
��J�� :�/����6�2�`����;�M�_�F16� ����n���������ȟ��Eҟ�����,� >�P�b���d�{�������������5�T��X��v���E ťmFѯ����� ��&�/�A�S�e�+p|�x�� � ��0����j�4pAT����6n�EL  �%ø�J���ʰJE��C�TR�Ѭ�TN��F�&��HAND_V�B[
�pK�� $F2{�6� �r�SW�D�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�(#�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������$uN���(!찙H������"CqE�N� a�DI��>�O�btD�Dpx�� ��2IxQA����q ��-��s �� ������ ��OMMEB��rr�QTVpPT�P ���qe�i�A���P�x ��yT�P�j� $DUM�MY9�$PS�_��RFq�0$:� ���!~q�� X����K�ST�s�ʰSBR��M�21_Vt�8$S/V_ERt�O��z����CLRx�A  O�r?p? Oր �� D $GLOB���#LO��Յ�$�o��P�!SYS�ADR�!?p�pT�CHM0 � ,x����W_NA���/�e�3�TS�R��l  (:]8:m�K6�^2m� i7m�w9m��9���ǳ� �ǳ���ŕߝ�9ŕ� ��i�L���m��_��_�_�TD�XSCR�E�ƀ�� ��STF���}�pТ6��sq] _v AŁ�s T����TYP�r��K��u�!u��Z�O�@IS�!��tsqUE{t� �Ȯ��H�S���!RS�M_�XuUNEX�CEPWv��CpS_ ��{ᦵ�ӕ���÷�ӎ�COU ��� �1�O�UET����r���PROGM�� FLn!$CUƕ�PO*q��c�I_��pH;� � 8\��N�_HE
p���Q��pRY ?����,�J�*��;�O�US�� � @�d���$BUTT��R@���COLU�M�íu�SERV<c#=�PANEv Ł�� � �PGE�U�!�F��9�)$�HELP��WRETER��)״���Q ������@� P��P �IN��s��PNߠw v�1������ ���L�N�� ����_���k�$H��M T�EX�#����FLA�n +RELV��DP4p�������M��?,��ӛ$����P�=�USRVIE�WŁ� <d��pU:�p0NFIn i��FOCU��i�PR�ILPm+�q��T�RIP)�m�U9Njp{t� QP��XuWARNWud�S�RTOLS�ݕ�t����O|SORN��'RAUư��T��%���VI|�zu�� $�PATH�g��CACHLsOG6�O�LIMyb�M���'��"�HOS�T6�!�r1�R��OBOT5���I%Ml� D�C� g!���E�L���i�VCPU_AVAILB�VO�EX7�!BQNL��(���A�� Q��Qq ��ƀ�  Qp�C���@$TO�OL6�$�_JM�P� �I�u�$SS�!$sqVS�HIF��|s�P �p�6�s���R���OSURW�pRGADIz��2�_�q��h�g! �q)�L�Uza$OUTP�UT_BM��I�ML�oR6(`)�@T;IL<SCO�@Ce�;��9��F�� T��a��o�>�3�P����w�2u���P{t��%�DJU���|#�WAIT�������%ON�E��YBOư �� $@p�%�C�SBn)TPE��NEC��x"�$t$\���*B_T��R��@�%�qR� ���sB�%�tM�+��t�.�F��R!݀��OPm�MA]S�_DOG�OaT	�D����C3S�	�>O2DELAY���e2JO��n8E��Ss4 '#J�aP6%�����Y_��O2$��2���5��`? sqZ�ABCS��  �$�2��J�
sp��$$CLAS�����AB�sp'@@VIRT��O.@gABS�$�1 <E�� < *AtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v�p����M@[�AXLրtK�*B�dC  ����IN��ā��PRE������LA�RMRECOV c<I䂥�NG��� \K	 A �  J�\�M@PPL�IC�?<E��E�Hand�lingTool� �� 
V7.�50P/28[� � �X���
��_SW�� UPn*A� ��F0ڑ䢒��A����� 20��*A����:���(�FB 7DA5��� '@Y��@��None엃���� ���T��*A4I�Wxl�_��V��t��g�UTOB��ค����HGAPCON8@��LA��U��oD 1<EfA���������� /Q 1שI Ԁ��Ԑ�:�i�n�����#B)B g���\�HE��Z�r�HTTHKY��$BI�[�m��� ��	�c�-�?�Q�o�u� �ϙϫϽ�������� _�)�;�M�k�q߃ߕ� �߹��������[�%� 7�I�g�m����� ��������W�!�3�E� c�i�{����������� ����S/A_e w������� O+=[as� ������K// '/9/W/]/o/�/�/�/ �/�/�/�/G??#?5? S?Y?k?}?�?�?�?�? �?�?COOO1OOOUO gOyO�O�O�O�O�O�O ?_	__-_K_Q_��(��TO4�s���DO_CLEAN��e��S�NM  9� �9oKo]ooo�o�DSPDRYR�_&%�HI��m@&o�o �o#5GYk} ����"���p�Ն# �ǣ�qXՄ���ߢ��g�PLUGGpҠ�Wߣ��PRC�`B`9��o�=��OB��oe�SEGF��K������o%o�����#�5�m���LAP�oݎ���������� џ�����+�=�O�|a���TOTAL�|.���USENUʀ�׫ �X���R(�R�G_STRING� 1��
�kM��Sc�
���_ITEM1 �  nc��.�@�R�d� v���������п������*�<�N�`�r��I/O SIG�NAL��Tr�yout Mod�e�Inp��S�imulated��Out���OVERR�` =� 100�In� cycl����Prog Abo�r�����Sta�tus�	Hea�rtbeat��MH FaulB�K�AlerUم�s� �ߗߩ߻��������� �S���Q� �f�x�������� ������,�>�P�b��t�������,�WOR ������V��
. @Rdv���� ���*<N`PO��6ц�� o�����// '/9/K/]/o/�/�/�/��/�/�/�/�/�DEV�*0�?Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O>�OPALTB��A ���O�O__,_>_P_ b_t_�_�_�_�_�_�_��_oo(o:o�OGRI�p��ra�OLo�o�o �o�o�o�o*< N`r������`o��RB���o� >�P�b�t��������� Ώ�����(�:�L��^�p����PREG �N��.�������� *�<�N�`�r������� ��̯ޯ���&��Ϳ�$ARG_��D ?	���i���  �	$��	[�}�]}���Ǟ�\�S�BN_CONFIOG i��������CII_SA_VE  ��۱�Ҳ\�TCELLSETUP i��%HOME_I�O�͈�%MOVq_�2�8�REP����V�UTOBAC�K
�ƽ�FRA:\�� ��Ϩ���'` ��������  ����$�6�c�Z�lߙ��Ĉ���������� ���!凞��M�_�q� ����2�������� �%�7���[�m���� ����@�������!3E$���Jo��������INI��@��ε��MESSAG����|q��ODE_D$����O,0.��P�AUS�!�i� ((Ol��� ����� /�/ /$/Z/H/~/l/�/�'�akTSK  �q�����UPDT�%�d0;WS�M_CF°i��еU�'1GRP Y2h�93 |�B���A�/S�XSCRDv+11
1; ����/�?�?�? OO $O��߳?lO~O�O�O �O�O1O�OUO_ _2_�D_V_h_�O	_X���G�ROUN0O�SU�P_NAL�h�	��ĠV_ED� 1�1;
 �%-BCKEDT-�_0`�!oEo$���a(��o�����ߨ���e2no_˔o�o�b���ee�o"�o�oED3�o�o ~p[�5GED4� n#�� ~�j���ED5Z��Ǐ6� ~p���}���ED6�� ��k�ڏ ~G���!�3�ED7��Z��~� ~p�V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W��Ư
}3�����CRo�����3�տ@�����P�PNO_D�EL�_�RGE_U�NUSE�_�TLA�L_OUT �q�c�QWD_AB�OR� �΢Q��IT_R_RTN����ONONSe����CAM_PAR�AM 1�U3
� 8
SONY� XC-56 2�34567890��H � @����?���( SАV�|[r؀~�X�HR5k�|U�Q��߿�R57����A�ff��KOW�A SC310M�|[r�̀�d @6�|V��_�X� ����V��� ���$�6���Z�l��CE_R�IA_I857�F�1��R|]]��_LIO4W=V� ��P<~�F<��GP 1�,����_GYk*Cg*  ��C1� �9� @� G� �CVLC]� d� l� Es�R� ��[�Um� v� � �� _�� C�� �"��|W��7�HEӰO�NFI� ��<G_�PRI 1�+ P�m®/���������'CHKPA�US�  1E� ,�>/P/:/t/^/ �/�/�/�/�/�/�/?�(??L?6?\?�?"OƩ����H�1_MkOR�� �Xa�Biq-���5 	 �9 O�?$OOHOZK�2	���=9"�QI?55��C�PK�D�3P������a�-4�O__|Z
�OG_�7�PO�� ��d6_��,xV�ADB����='�)
mc:cpmidbg�_�`��S:�  Y�PZ���Up�_)o�S�  �C@# 	�f�P�_mo8j�  ߏ`y�QiXo�o9i�(�U(��� Qig�o�o�lw
�xOkf�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@R����Ja`(Ж�Ao=L���zMC�21�=��9���4��=�n׾�Cz � BHBCCPUe�B�_B�y�;��>C����CnSZE@E?�{hD]^Dٿ�?r����D���^��G	���F��F���Cm	fF�O�OF�ΫSY���vJqG���Em�(�%.���1(��<�qѪG�&q��Ң �̢ a�D�j���E�S\��X�EQ��EJP F�E��F� G����F^F E��� FB� H,�- Ge��H3�Y���  >�?33 ���xV�  n2xQ@��5�Y��8B� A�AST<7#�
� �_'��%��wRSMOFSb���~2�yT1�0�DE �O@b �
�(�;�"�  Q<�6�z�R���?,�j�C4��SZm�E &q�{�m�C��)B-G�Cu�@$�q���T{�FPROG %i����c��I��� �Ɯ�f�KEY_TBL  �v�M�u� �	
��� !"#$�%&'()*+,�-./01c�:;�<=>?@ABC��pGHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����p����͓��������������������������������������������������?������!j��LCK��.�j���S�TAT���_AU_TO_DO���W�/�INDT_EN�B߿2R��9�+�Ty2w�XSTOP\��2TRLl�LET�E����_SCR�EEN i_kcsc��U���MMENU 1 ~i  <g\ ��L�SU+�U��p3g� ������������2� 	��A�z�Q�c����� ����������. d;M�q��� ���N%7 ]�m���/ ��/J/!/3/�/W/ i/�/�/�/�/�/�/�/ 4???j?A?S?y?�? �?�?�?�?�?O�?O -OfO=OOO�OsO�O�O �O�O�O_�O_P_Sy��_MANUAL���n�DBCOU�R�IG���DBNUIM�p��<���
�Q�PXWORK 1!R�ү�_oO.o�@oRk�Q_AWAYz�S��GCP ��9=��df_AL�P߄db�RY�������X_�p 1"�� , 
�^���o �xvf`MT�I^�rl@|�:sONTIM�כ����Zv�i
�õ�cMOTNEN�D���dRECOR/D 1(R�a��ua�O��q��sb �.�@�R��xZ���� ���ɏۏ폄���#� ��G���k�}�����<� ş4��X���1�C� ��g�֟��������ӯ �T�	�x�-���Q�c� u����������>�� ��)Ϙ�Mϼ�F�� �ϧϹ���:������� %�s`Pn&�]�o��ϓ� ~ߌ���8�J����� 5� ��k����ߡ�� J�����X��|��C� U����������0������	��dbTOL�ERENCqdB�ܺb`L�͐PCS_CFG )�k�)wdMC:\�O L%04d.C�SV
�`c�)sA� �CH� z�`�)~���hMRC_OUT *�[��nSGN �+�e�r��#�1�0-MAY-20� 08:56*V1�5-JANj10�:51�k P/Vt��)~�`�pa�m��P�JPѬVE�RSION �SV2.0.�8.|EFLOGI�C 1,�[ 	DX�P7)�PF."�PROG_ENB��o�rj ULSew ��T�"_WRST�JNEp�V�r`dEM�O_OPT_SL� ?	�es
 ?	R575)s7)��/??*?<?'�$TO  �-��?&[V_@pEX�Wd�u��3PATH ASA\�?�?O�/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C��SqqF�PMAU�� t/XrMSWR.D�i�a.|S/�Z!D_N�O0__T_C_�x_g_�_�tSBL_/FAUL"0�[3w/TDIAU 16M�a�p�A12�34567890gFP?BoTofo xo�o�o�o�o�o�o�o ,>Pb�S�p-P�_ ���_s �� 0`����� )�;�M�_�q����������ˏݏ��|)UM�P�!� �^�T�R�B�#+�=�PME�fEI�Y_TEMP9 È�3@�3A �v�UNI�.(YN_BRK 2Y�)EMGDI_S�TA�%W!bՐNC�2_SCR 3��1o"�4�F�X�fv ���������#��ޑ14����)�;������ݤ5��� ��x�f	u�ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/߭P�b�t�� �� xߞ߰���������
� �.�@�R�d�v��� �����������*� <�N���r��������� ������&8J \n������ ��"`�FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/4? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O ?�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�O�O�o�o�o
 .@Rdv�� �������*� <�N�`�r����o���� ̏ޏ����&�8�J� \�n���������ȟڟ�����H�ETMO�DE 16���� ��ƨ
�R�d�v�נRROR�_PROG %fA�%�:߽�  ���TABLE  �A������#�L�R�RSEV_NUM�  ��Q���K�S���_AUT�O_ENB  ���I�Ϥ_NOh� �7A�{�R� W *���������	���^�+��Ŀֿ���HISO�͡I�}�_ALM 18A�� �;�����+�e�wωϛϭϿ�r�_H���  A����|��4�TCP_VER !A��!����$EXTL�OG_REQ�9�{�V�SIZ_�QԿTOL  ͡D�z��A Q�_BWD����r���n�w_DI�� 9���}�z�͡m���S�TEP����4��O/P_DO���Ѡ�FACTORY_�TUN�dG�EATURE :�����l�Ha�ndlingTo�ol ��  - �CEngli�sh Dicti�onary��OR�DEAA V�is�� Mast�er���96 H���nalog I�/O���H551���uto Sof�tware Up�date  ��J���matic B�ackup��Pa�rt&�gro�und Edit���  8\apCamera��F��t\j6R�e�ll���LOADnR�omm��shq�ޝ�TI" ��co<��
! o����pane�� 
�!��tyle �select��H�59��nD���onoitor��48�����tr��Reli�ab���adin�Diagno�s"����2�2 ua�l Check �Safety UIF lg\a���hanced Rob Serv �q ct\��lU?ser FrU���DIF��Ext.� DIO ��fi�A d��end.r Err L@��KIF�r��  �����90��FCTN_ MenuZ v'���74� TP I�n��fac  SU (G=�}p��k Excn �g�3��High�-Sper Ski.+�  sO�H9 � �mmunic!�oknsg�teur� 4����V�����conn��2��E�N��Incrs�tru���5.f�dKAREL Cmd. L?�uaA� O�Ru�n-Ti� Env�����K� ��+%�sn#�S/W��74��LicenseT��  (Au* o�gBook(Sy���m)��"
�MACROs,~V/Offse��ap��MH� �����pfa5�Mech�Stop Pro�t��� d�b i��Shif���j545�!xr ��#�ޜ�,[�b od�e Switch.��m\e�!o4=.�& pro�4���g��Mult�i-T7G��net.Pos �Regi��z�P>��t Fun����3 Rz1��Numx �����9m�1� � Adjuj��1' J7�7�* ����6tatuq1EI�KRDMto}t��scove�� ��@By- }u'est1�$Go� � �U5\SNPX� b"���YA�"Libr����#��1 �$~@h�pd]0��Jts in V�CCM�����0� 8 �u!��2 R�0��/I�08��TM�ILIB�M J9u2�@P�Acc>��F�97�TPTXl�+�BRSQelZ0�M8 Rm��q%���692��Unex�ceptr mot}nT  CVV�P���KC����+-|��~K  II)�VSP CSXC�&�.c�� e�"�� t��@Wew�A3D Q�8bvr ngmen�@�iP� �a0y�0�pfGr�idAplay �!� nh�@*�3R�1M�-10iA(B2�01 �`2V"  �F���scii�l�oad��83 M��l����Guar��d J85�0�mP�'�L`���stuaPsat�&]$Cyc���|0ori_ x%D7ata'Pqu����ch�1��g`� j6� RLJam�5��|��IMI De-By(\A�cP" #^0�C  etkc>^0asswo%q�)650�ApU�Xsnt��Pven�C�TqH�5�0Y�ELLOW BO�?Y��� Arc�0v�is��Ch�We{ldQcial4Izt�Op� ��gs֛` 2@�a��pofG yRjT1 �NE�#HT� xy�Wb��! �p�`g�d`���p\� =P��JPN ARCP*�PR�A�� O�L�pSup̂fi�l�p��J�� ��cro�670�1C~E�d���SS�pe�teex�$ �P� So7 �t� ssagN5 D<Q�BP:� �9 "0F�QrtQC��P�l0dpn�笔�rpf��q�e�ppma�scbin4ps{yn�' ptx]0�8�HELNCL� VIS PKGsS �Z@MB �&��B J8@IP�E GET_VA�R FI?S (U�ni� LU�OOL�: ADD�@29�.FD�TCm���E�@DVp���`A�Т�NO WTWTE'ST �� f�!���c�FOR ��EC�T �a!� ALS�E ALA`�CP?MO-130��� �b D: HANG FROMg��2���R709 DR�AM AVAIL�CHECKS 5�49��m�VPCS� SU֐LIMC�HK��P�0x�FF� POS� F�� �q8-12 oCHARS�ER6��OGRA ��Z@A�VEH�AME��.#SV��Вאn$���9�m "y�TRC�v� SHADP�U_PDAT k�0���STATI��� �MUCH ���T�IMQ MOTN�-003��@O�BOGUIDE DAUGH���b��@$tou� �@C�y �0��PATH�_�MOVET�� �R64��VMXP�ACK MAY ?ASSERTjS��oCYCL`�TA���BE COR 7�1�1-�AN��RC� OPTIONS�  �`��APSH;-1�`fix��2�SO��B��XO򝡞�C_T��	�i��0j���du�byz p w1a��y�٠HI�����U�pb XSPD� TB/�F� \h�chΤB0���EN�D�CE�06\Q�p�{ smay n�@�pk��L ��tOraff#�	� ���~1from s�ysvar sc�r�0R� ��d�DJ�U���H�!A��/���SET ERR��D�P7����ND�ANT SCRE�EN UNREAO VM �PD�D���PA���R�IO� JNN�0�FI���B��GROUNנD Y�Т٠��h�SVIP 53� QS��DIGIT VERS��ká��NEW�� P06z�@C�1IMAG�hͱ���8� DI`<���pSSUE�5���EPLAN JO�N� DEL���15�7QאD��CAL�LI���Q��m���I�PND}�IMG oN9 PZ�19���MNT/��ES ܏��`LocR Ho�l߀=��2�Pn� P�G:��=�M��ca�n����С: 3�D mE2view� d X��eat1 �0b�pof Ǡ�"HCɰ�ANN�OT ACCESS M cpie�$Et.Qs a� l�oMdFlex)a:z��w$qmo G�s�A9�-'p~0��h0p�a��eJ AUTcO-�0��!ipu@�Т<ᡠIABLE�+� 7�a FPLNs: L�pl m6� MD<�VI�и�WIT HOC�;Jo~1Qui��":��N��USB�@�P�t & remo�v���D�vAxisO FT_7�PGɰ�CP:�OS-1�44 � h s s268QՐOST�p�  CRASH �DU��$P��WO�RD.$�LOG3IN�P��P:	�0��046 issu�eE�H�: Sl�ow st�cB�`6����໰IF��IMPR��SPO�T:Wh4���N1S�TY��0VMGR��b�N�CAT��4�oRRE�� � �58�1��:%�RT�U!Pe -M a�SE�:�@pp���AGpL���m@allء�*0a�OCB W�A���"3 CNTw0 T9DWroO0alarm�ˀm0d t�M�"0�2|�s o�Z@OME<�x� ��E%  #1-�gSRE��M�st}0g     5�KANJI5no� MNS@�IN�ISITALIZf'� E�f�we���6@� dr�@ fp� "��SCII �L�afails �w��SYSTE0[�i��  � Mq��1QGro8�m n�@vA����&���n�0q��RWRI� OF Lk��� �\ref"�
�up�� de-rela��Qd 03.�0S�Schőbetw�e4�IND exm ɰTPa�DO� �l� �ɰGig�E�soperab�il`p l,��H0cB��@]�le�Q0cflxz�Ð���OS {����v4pf;igi GLA�$��c2�7H� lapn�0ASB� If��=g�2 l\c�0���/�E�� EXCE 㰁�P���i�� o0��Gd`]Ц�yfq�l lxt��EFal��#0�i�xO�Y�n�CLOS��SRNq1NT^�F��U��FqKP�ANIOO V7/ॠ1�{8����DB �0���ᴥ�ED��DET�|�'� �bF�NLwINEb�BUG�Tt���C"RLIB���A��ABC JA�RKY@��� rk�ey�`IL���PRr��N��ITGAR� D$�R �Er *�T��a�U�0��h��[�ZE V� T�ASK p.vr��P2" .�XfJ�s�rn�S谥dIBP�	c���B/��BU]S��UNN� j0�-�{��cR'���L�OE�DIVS�CU�Ls$cb����BW !��R~�W`P�����IT(঱tʠ�O=F��UNEXڠ+�Ҧ�p�FtE��SV�EMG3`NML �505� D*�CC_SAFE�P*� �8ꐺ� PET��'P��`�F  !���IQR����c i S>�� K��K�H G_UNCHG��S�/MECH��M���T*�%p6u��tPORY LEAK�9J���SPEgD���2V 74\GR�I��Q�g��CTLN��TRe @�_�p l���EN'�IN�������$���r��T3\)�i�STO�A�s�L��͐X	���qb��Y� ��TO2�J m��0F<�K����SDU�S��O��3 9�J F�&��~�SSVGN-1#�I���RSRwQDAU��Cޱ� �T6�g��� �3�]���BRKCTqR/"� �q\j5�p�_�Q�S�qINVJ0D ZO�Pݲ���s ��г�Ui ɰ̒�a��DUAL� J5�0e�x�RVO117 AW�TH!Hr�%�N�247%�528��|�&aol ���RP���at�Sd�cU���P,�LER��iԗQ<0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�c�豓�{�U��ROP� 2�b�pB��IT�P4M��b !A�Ut c0< � pleste�N@� z1�^qR635 (AccuCal2kA=���I) "�ǰ�1a\�Ps��ǐ� �bЧ0P򶲊���i�g\cbacul "A3p_ �1��ն|���etaca��AT���PC�`����v�_p�.pc!�x���:�circB���5�tl��Bɵ�:�Cfm+�Ί�V�b�����r�upfrm.0����ⴊ�xed��Μ��~�pedA�D �|}b�ptlibB�� �_�rt��	��_\׊ۊ�6�fm �݊�oޢ�e��̆Ϙ�"��c�Ӳ�5�j>���F��tcȐ��	�r�����mm 1��T�sl^0��T�mѡ�#�rm3��ub Y�q�gstd}��pl;��&�ckv�=�r�vf0�䊰��9�vi�����ul�`�0fp�q ��.f��� da�q; i Data Acquisi���n�
��T`��1�89��22 �DMCM RRS�2Z�75��9 3� R710�o5�9p5\?��T ="��1 (D�T� nk@��������E �Ƒȵ��Ӹ�etdmm ��ER�����gE��1�q\mo ?۳�=(G���`[(

�2�` ! �|@JMACRO���Skip/OffCse:�a��V�4oy9� &qR662�H��s�H�
 6Bq�8����9Z�43� J77� 6�J783�o ��n��"v�R5IKC~Bq2 PTLC�vZg R�3 (�s, ��������03�	зJԷ\s�fmnmc "M�NMC����ҹ�%m;nf�FMC"Ѻ|0ª etmcr� ��8���� �,[�Df��   874\Oprdq>,jF0����axisHP�rocess A�xes e�rol�^PRA
�Dp� 5�6 J81j�59� 56o6� ���06w�690 98� [!GIDV�1��2(x2��2ont�0�
� ���m2���?C���etis "IS�D��9�� FpraxRAM�P� D�чdefB�,�G�i�sbasicHB��@޲{6�� 708*�6��(�Acw:� �����D
�/,��AMOX�� ��DvE��?;Td��>Pi� RAFM';�]�!PAM�V�W�E�e�U�Q'
bU�75��.�ceNe� nterface^4�1' 5&!54�K��b(Devam±�/@�#���/<�Tane`�"DNEWE���bt�pdnui �AI��_s2�d_rso!no���bAsfjN�>�bdv_arFvf�`xhpz�}w��hkH�9xstc��gApocnlGzv{�ff� �r���z�3{q�'Td>pcham�pr;e�p� ^59�77��	܀�4}0��m�Ɂ�/�����lf�!�p�cchmp]aMP�&B�� �mpevp�����pcs���YeS�� Macr%o�OD��16Q!)* �:$�2U"_,��Y�(PC ��$_;������o��J�gege=mQ@GEMSW�~Z>G�gesndy��OD�ndda��S��csyT�Kɓ�su^҈����n�m���L�� ' ���9:p'ѳ�޲��spotplusp���`-�W�l��J�s��t[�׷p�key�ɰ�$��s�-����m���\featu 0FEAWD�woolo�srn'!2 p���a�As3���tT.� (N. A.)��!e!�J# (j�,��oBLIB�oD -�.�n��k9�"K��u[-��_���p� "PS�EqW����wop "sEЅ�&�:�J� �����y�|��O8�� 5��Rɺ���ɰ[��X �������%�(
���q HL�0k�
�z�a!�B�Q�"( g�Q�����]�'�.� ����&���<�!ҝ_�#��tpJ�H�~Z��j� ����y������2�� e������Z����V�� !%���=�]�͂��^2n�@iRV� on�IQYq͋JF0� 8ހȖ`�	(^�dQueue���X\1�ʖ`��+F1tpvtsn���N&��ftpJ0v �RDV�	f��J1� Q���v�en���kvstk��m�p��btkclrqq���get�����r��`ka�ck�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�mc�N+v3�_� �����.v�/\=jF��� �`Q��΋ܒ�N50 (F�RA��+��͢fraparm��Ҁ�z} 6�J643p:~V�ELSE
#��VAR $SGSYSCFG.$�`�_UNITS 2��DG~°@�4Jgfr8��4A�@FRL-��0 ͅ�3ې���L�0NE �:�=�?@�8�v�9�~Qx304��;�BP�RSM~QA�5TX�.$VNUM_O�L��5��DJ507���l� Funct�ʂ"qwAP��琉�3# H�ƞ�kP9jQ�QA5ձ� ��@jLJzB J[�6N�kAP���|�S��"TPPR����QA�prnaS�V�ZS��AS8Dj5150U�-�`cr�`8 ���ʇ�DJR`jYȑH�  �Q ��PJ6�a21��4�8AAVM �5�Q�b0 lB�`T�UP xbJ5�45 `b�`616����0VCAM� 9�CLIOn b1�5 ����`MSC8�
rP �R`\sSTY�L MNIN�`J�628Q  �`N�REd�;@�`SCH� ��9pDCSU �Mete�`ORSsR Ԃ�a04 kREIOC �a]5�`542�b9vp�P<�nP�a�`�R�`7��`�MASKg Ho�.r7 �2��`OCO :��r3@��p�b�p���r0X�|�a�`13\mn�a39 HRM"�q��q��LCHK>�uOPLG B��a�03 �q.�pHC�R Ob�pCpPo�si�`fP6 is�[rJ554�òpDSW�bM�D�pqR�ag37 }Rjr0 �1��s4 �R6�7��5�2�r5 �2�r7 �1� P6���Reg�i�@T�uFRKDM�uSaq%�4�`�930�uSNBA��uSHLB̀\suf"pM�NPI��SPVC�J52�0��TC�`"MN�рTMIL�IF�V�PAC W�pT�PTXp6.%�T�ELN N Me��09m3UEsCK�b�`UFR�`ކ�VCOR��VI�PLpq89qSXC��S�`VVF�J�T�P �q��R626.l�u S�`Gސ�2?IGUI�C���PGSt�\ŀH8�63�S�q�����q3u4sŁ684��0�a�@b>�3 :B��s1 T��96 .��+E�51 y�q5�3�3�b1 ���b1� n�jr9 ���`V�AT ߲�q75 �s�F��`�sAWSM<��`TOP u�ŀ�R52p���a80 �
�ށXY q���0� ,b�`885�QXрOLp}�"pE࠱;tp�`LCMD���ETSS���6 |�V�CPE oZ1��VRCd3
�NL:H�h��001m2Epƌ�3 f��p��4 _/165C��6l�ꌰ7PR��008� tB��9 -20-0�`U0�pF�1޲1 ��޲2L"���p���޲4��5 \�hmp޲6 RBC�F�`ళ�fs�8 ��Ҋ��~�J�7 r'bcfA�L�8\PC����"�32m0u�n��K�Rٰn�5 5E7W
n�9 z��g40 kB��3 ���6ݲ�`00iB/���6�u��7�u��8` µ������sU0�`��t �1 05\rb��2 E���K�Ȇ�j���5˰��60 ��a�HУ`:�63�jA0F�_���F�7 ڱ݀�H�8�eHЋ��cU0$��7�p��1u��y8u��9 73��L����D7� ��5t󮊱97 ��8U�1(��2��1�1:���Eh��1np�"��8(�{U1��\pyl���,࿱v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6 B���цp��1�����1�`͵155�ض157 �2��6A2�S����1b�H�2����1Π"�2��&�B6`�1<c�34 7B�5 DR���8_�B/��187y uJ�8 06��90 rBn�1 (���202 0EWE,ѱ2^��2��90�cU2�p�2��2 b��4��2�a"RB4����9\�U2�`w�<l���4 60Mp��7������b�s
5� ��3����pB"9� 3 ����`ڰR,:7 �2��V�2��5���2^��a^	9���qr����n�A5����5᥁"�8a�$Ɂ}�5B���5���B�`UA���� ��86 V�6 S�0��5�px�2�#�529 �2P^�b1P�5~�A2`���&P5��E8��5��u�!�5���ٵ544��5��R��ąP nB^z�c �(�4�����U)5J�V�5��1�1^���%�����5 b�21��gA��58�W82� rb��5N�E�5890r� 1�95 �"���� ��c8"a��|�L ���!J"5|6��^!�6��B�"8�`#��j+�8%�6B�AME�޶"1 iC��62�2�Bu�6V��d� 4���84�`ANRS�P�e/S� C@�5� �6� ��� \� ��6� �V� 3t��� T20CA�R���8� Hf� 1DH�� �AOE� �� ;,[|�� �0\�,� �!64K��ԓrA|� �1 (M-7�!/50T�[PM��P�Th:1�C�#Pe�� �3�0� 5`M7�5T"� �D8p� ��0Gc� u�4��i1-O710i�1� Skd�7j�?6�:-HS,� �RN�@�UB�xf�X�=m75sA*A6an���!/CB�B2.6A �0;A�CIB@�A�2�QF1�UB2�21� /70�S� �4�����Aj1�3p�p��r#0 B2\m*A@C��;bi"i1K�u"�A~AAU� imm7c7��ZA@I�@�D�f�A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A �5*A�EA�5B�4>\77
B7=Q�D�2�Q�$B�E7�C�D/qAHEE�W7�_|`jz@�  2�0�Ejc7�`�E"l7�@7�A
1�EH�V~`�W2%Q�R9�.�@0L_�#����"�A���b��H3s=rA/2�R5nR4�74r�NUQ1ZU�A�s\m9
1M92L2�!F!^Y:�ps� 2ci��-?�qhimQ�t  w043 �C�p2�mQ�r�H_ �H20�Evr�QHsXBSt#62�q`s����� x��Pxq350_*AF3I)�2�d�u0�@�� '4TX�0�pa3i1A3sQ25�c&��st�r�VR1%e�q0
��j1��O2� ���A�UEiy�.�‐ ț0Ch20$CXB79�#A�ᓄM Q1]�~�� 9�Q��?PQ��qA !Pvs� 5	15aU����?PŅ���ဝQ9#A6�zS*�7�qb5��1����Q��00P(��V7]u�aitE1�� �ïp?7� !?�z��{rbUQRB1PM=��Qa9��H��QQ�25L�������Q��@�L��8ܰ��y00�\ry�"R2BL��tN  ���; �1Df��2�qeR�5���_b�3��X]1m1lcqP1�a�E�Q� 5F����!y5���@M-16Q� � f���r��Q�e� p��� PN�LT_�10��i1��9453��@8�e�|�b1l>F1@u*AY2�
��R8�Q0����RJ�J3�D}T� 85
Qg�/0��*A�!P�*A�Ð𫿽�2,ǿپ6t�6=Q��`�Pȓ��� AQ� g�*ASt]1^u�ajr I�B����~�|I�b�L�yI�\m�Qb�I�u�z�A�c3Apa9q� B6S��S��m���}��85`N�N�  �(M���f1��@�6����161��5�s`�SC��U��A�����5\set06�c����10�y�h8��a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��@���5�B��B��h`� F���X0���A:���C�M��AZ��@��4�6@i����� e�O�-	 ���f1��F �ᱦ��1F�Y	���T6HL3��U66~`���U�9dU�9D20Lf0�� Qv� ��fjq��N�� ����0v
� ��i	�\	��72lqQ2������� \chn?gmove.V���d���@2l_arf	�f~��6� �����9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�AX]��V�1\�Qn�BJ�2W�EM!`5���)�#:�64��F�e50S�\��0 �=�PV���e���逕��E�����mw7shqQSH"U��)��9�!A��(����� ,[�9�ॲTR1!��&,�60e=�4F���2��2��	 R-��� ��������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2�"�2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D��� 5V��@2cVE��p��dT��pt갖�1L~E��#�F�Q��9E�#De1/��RT��59���	��A�EiR������9o\m20�20��+�-u�19r4�`�E1 �=`O9`�1"ae���O�2��_$W}am�41�4�3�/d1c_std��1)Ķ!�`_T��r�_ 4\jdg�a�q�PJ %!~`-�r�+bgB���#c300�Y�5j�QpQb1�bq��vB��v25�U������qm43� �Q<W�" PsA��e��� �t�i�P�W.��c��FX.�e�kE14��44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2-a��2A;_2��QW�2�bF�(�V11�2�3�`��X5�Ra21B�J*9�a:88rJ9X�l5�m1a�0���*���(85�&� ������P6���RB,52&A����,fA�9IfI50\u�z�O@V
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq� &ŦP1��vB)e�m�x����1p� �1�Df��27�F�K�AREL Use{ S��FCTN��� J97�FA+�� (�Q޵�p%�)?��Vj9F?(�j�Rtk208 "Km�6Q�y�j��iæPr��9�s#��v�krcfp�RCFt3���Q~��kcctme�!�ME�g����6�ma�in�dV�� ��r!u��kDº�c���o�����J�dt�F �»�.vrT�f������E%�!��5�FRjK73B�K���UER��HJ�O  J�� (ڳF���F�q�Y��&T��p�F�z��19�tAkvBr���V�h�9p�E�y�<�k������8;�v���"CT��f ����)�
І��)�V 	�6���!��qFF�� �1q���=�����O�?� $"���$��je��TCP Aut�r~�<520 H5��J53E193��9V��96�!8��9���	 �B574��52��Je�(�� Se %!Y�����u��ma�Pqtool�ԕ�������conre�l�Ftrol Reliable�RrmvCU!��H51������ a551xe"�CNRE�I�c�&��it�l�\sfutst �"UTա��"X�\�u��g@�i�6Q]V0H�B,Eѝ6A� �Q �)C���X��Yf�Iȴ1|6s@6i��T�6IU��vR�d�
$e0%1��2�C58�E6���8�Pv�iV4OFH5�8SOeJ� mvBM6E~O58�I�0�E�# +@�&�F�0���F�P 6a���)/++�</N)0\tr1�����P� ,[�ɶ�rma;ski�msk�aA����ky'd�h	A	�P��sDisplay�Im�`v����J8�87 ("A��+He<ůצprds��I�T�ǅ�h�0pl�2�R�2��:�Gt�@��PRD�TɈ�r�C�@Fpm��D�Q�Asca��� V<Q&��bVvbrl�eې@��^S��8&5Uf�j8710��yl	��Uq���7 �&�p�p��P^@�P�firmQ����Pp� 2�=bk�6�r�3��6���tppl��PL ���O�p<b�ac�q	� �g1J�U�d�J��gait_9e��Y�&���Q���	�Shap���erationx�0��R67451tj9(`sGen� ms�42-f��r�p�50����2�rsgl�E���p�G���qF�205�p�5S���Ձ�ret�sap�BP�O�\s>� "GCR�ö?� �qngda�G ��V��st2axU�b�Aa]��bad�_|�btputl/��&�e���tplibB_��=�2.����5�Ό�cird�v�sl8p��x�hex��v��re?�Ɵx�key��v�pm��x�u9s$�6�gcr��F�������[�q27j92|�v�ollismq�Sk�9O�ݝ� (Gpl.���t��p!o���29$Fo8��cg7�no@�tptcls` CLS�o�b�\�#km�ai_
�s>�v�o	�t�b���ӿ�E��H��6�1en�u501�[m��u�tia|$calm�aUR��CalMa;teT;R51%�i=1]@-��/V� ��Z��� �fq1�9 "KA9E�L����2m��CLMTq�S#��et �LM3!} �:F�c�nspQ�cӞ��c_moq��� ���c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ����N�ve��C�clm��&Ao# �|$fin�de�0ST�D ter Fi?LANG���R��
��n3��z0gCen���r,�� ����J����� ��� K��Ú�=���_Ӛ����r� "FND�R�� 3��f��tguid�䙃N�."��J�tq�� ��������������J����_@������c��	m��Z��\fndr. ��n#>
B2p��Z�CP Ma�����C38A��� c��6� (���N�B����� �� 2�$�81��!m_���"ex�z 5�.Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$ �r*$��*$r*$%/s#�C�d/.,P�/0*ʲDPN��$���$�*�Gr�$k Ex�c�'IF�$MAS}K�%93 H5�%�H558�$548 H�$4-1�$��#21(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�4�9�0�4a�3�9j0"�M�49�4  �x�4�4tpsh��x�4�P�4- DQ� @�3�Q�4�R�4�pR%0 �2�r�4.b
E\���5�A�4��3adq\>�5K979":E�a~jO l "DQ^E^�3i�Dq ��4�R�O ?R�? ��q�5 ��T��3rAq�O�L#st�5~��7p�5��0REJ#�2�@av^Eͱ��F���4��.�5y �N� �2il(in8�4��31 JH1�2�Q4�251ݠ�4rmal� �3)�REo� Z_�æOx����4��^F�?onorTf��7_�ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4�REM���4yݱ"u@�RER5932fO��4�7Z��5lity,��U��e"Dil\��5��o ��798�7�?�25 �3hk9 10�3��FE�0=0|P_�Hl\mhm�5 ��qe�=$�^�
E���u�IAymptm`�U��BU��vste� y\�3��me�b�DvI� [�Qu�:F�Ub�*_��
E,�su��_ Er��ox���4�huse�E-�?�s�n�������FE��,�b#ox�����c݌," �������z��M�x�g��pdspw)� 	��9���b���(��1���c��Y� R�� �>�P���W��� �����'�0ɵ��[��͂���  ߤ ,[@� ��A�bum�pšf��B*�Bo!x%��7Aǰ60�BB�w���MC� (6�,�f�t I�s� ST��*��}B���z��w��"BBF
��>�`���)��\bbk968 "�X4�ω�bb�9vas69����etbŠb��X�����ed	��F��u�f� �seDa"������'�\��@,���b�ѽ�o6�$H�
�x�$�f���!�y���Q[�! tp�err�fd� T�Pl0o� Reco�v,��3D��R642 � 0��C@}s�� N@��(U�rr�o���yu2r���  �
  |����$$CLe�? �������������$z�_D�IGIT��������.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo�$j��+c:PRO�DUCTM�0\P_GSTKD��V&o�hozf99��D����$FEAT?_INDEX��xd���  �
�`ILECO_MP ;���#���`�cSETU�P2 <�e~�b�  N �a��c_AP2BCK� 1=�i  #�)wh0?{%&c����Q�xe%� I�m���8�� \�n����!���ȏW� �{��"���F�Տj� ��w���/�ğS���� �����B�T��x�� ����=�үa������ ,���P�߯t������ 9�ο�o�ϓ�(�:� ɿ^���Ϗϸ�G� ��k� �ߡ�6���Z� l��ϐ�ߴ���U��� y����D���h��� ���-���Q������ ���@�R���v���� )�����_�����* ��N��r��7 ��m�&�3�\�i
pP 2>#p*.VRc�*��� /���PC/1/OFR6:/].��/+T�`�/�/F%�/��,�`r/?�*.F�8?	H#&?e<��/�?;STM @�2�?�.K �?�=�iPendant Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OoO�O_:JPG  _J_�56_�O_�_��	PANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W �o�o�o)�Z4�o[��WI��
T�PEINS.XM)L��0\����qCustom Toolbar	���PASSWO�RDyFRS�:\L�� %P�assword ?Config��� ֏e�Ϗ�B0���T� f����������O�� s������>�͟b�� [���'���K��򯁯 ���:�L�ۯp����� #�5�ʿY��}��$� ��H�׿l�~�Ϣ�1� ����g��ϋ� ߯��� V���z�	�s߰�?��� c���
��.��R�d� �߈���;�M���q� �����<���`���� ��%���I������ ��8����n���! ��W�{"� F�j|�/� Se��/�/T/ �x//�/�/=/�/a/ �/?�/,?�/P?�/�/ �??�?9?�?�?o?O �?(O:O�?^O�?�O�O #O�OGO�OkO}O_�O 6_�O/_l_�O�__�_ �_U_�_y_o o�_Do �_ho�_	o�o-o�oQo �o�o�o�o@R�o v��;�_� ��*��N��G��� ���7�̏ޏm���� &�8�Ǐ\�돀��!� ��E�ڟi�ӟ���4� ßX�j��������į S��w������B�#���$FILE_D�GBCK 1=���/���� ( �)
�SUMMARY.�DGL���MD:����Dia�g Summar�y��Ϊ
CONSLOG�������D��ӱConsol�e logE�ͫ���MEMCHEC�K:�!ϯ���X�M�emory Da�ta��ѧ�{)}��HADOW���ϵ�J���Sha�dow Chan�gesM�'�-�?�)	FTP7Ϥ��3ߨ���Z�mme?nt TBD��ѧ�0=4)ETHERNET��������T�ӱEthe�rnet \�fi�guration�U�ؠ��DCSVR�F�߽߫�����%��� verif�y all��'�1�PY���DIFF������[���%��diff]�����1R�9�K��� ����X��CHGD������c��!r����2ZAS� ���GD���k��8z��FY3bI[� �/"�GD���s/�����/*&UPDA�TES.� �/���FRS:\�/�-�ԱUpdates� List�/��P�SRBWLD.C	M(?���"<?�/Y��PS_ROBOWEL��̯�?�?��? &�O-O�?QO�?uOO nO�O:O�O^O�O_�O )_�OM___�O�__�_ �_H_�_l_o�_�_7o �_[o�_lo�o o�oDo �o�ozo�o3E�o i�o���R� v���A��e�w� ���*���я`����� ����O�ޏs���� ��8�͟\�����'� ��K�]�쟁����4� ��ۯj������5�į Y��}������B�׿ �x�Ϝ�1���*�g� ����Ϝ���P���t� 	�ߪ�?���c�u�� ��(߽�L߶��߂�� ��(�M���q� ��� 6���Z������%��� I���B�����2������h����$FI�LE_� PR� ���������MDON�LY 1=.�� 
 ���q�� ��������~ %�I�m� 2��h��!/� ./W/�{/
/�/�/@/ �/d/�/?�//?�/S? e?�/�??�?<?�?�? r?O�?+O=O�?aO�? �O�O&O�OJO�O�O�O�_�O9_�OF_o_
VISBCKL6[*.VDv_�_.P�FR:\�_�^�.PVision� VD file �_�O4oFo\_joT_�o o�o�oSo�owo �oB�of�o�+ �������+� P��t������9�Ώ ]�򏁏��(���L�^� ������5���ܟk�  ���$�6�şZ��~������
MR_G�RP 1>.�L��C4  B���	 W������*u����RHB ��2� ��� ��� ���B�����Z� l���C���D��������Ŀ��K��L�57J�h�F��5UT+�QǱ�Ͳ��ֿ �G,�FI�/�E���.��9�:�]�@�'��A&�A}��_f�?��A}��r��E�� F@ ��������J��NJk��H9�Hu���F!��IP�s��?����(�9��<9�8�96C'6<�,6\b��B��Y%���A|��=�@�eߋ�^�A� �߲�v���r������ 
�C�.�@�y�d��� �����������?��Z�lϖ�BH�� y��R�?_��E�������
0�P=��P�H
��ܿ�� �B���/ ��@�33:��.�g&�/@UUU�U��q	�>u.�?! rX��	�-�=[z�=�̽�=V6<�=��=�=$q������@8�i�7G��8�D��8@9!�7��:����D��@ D�� C�,���C������Q� ,/������/M��/ q��/�/�/�??:? %?^?p?[?�??�?�? �?�? O�?�?6O!OZO EO~OiO�O�O�O�OW� �ߵ��O$_�OH_3_l_ W_�_{_�_�_�_�_�_ o�_2ooVohoSo�o wo�o�i��o�o�o ��);�o_J�j �������%� �5�[�F��j����� Ǐ���֏�!��E� 0�i�{�B/��f/�/�/ �/���/��/A�\�e� P���t��������ί ��+��O�:�s�^� p�����Ϳ���ܿ�  ��OH��o�
ϓ�~� �Ϣ����������5�  �Y�D�}�hߍ߳ߞ� �������o�1�C�U� y��߉������ ������-��Q�<�u� `��������������� ;&_J\� ���������ڟ �F�j4���� �����!//1/ W/B/{/f/�/�/�/�/ �/�/�/??A?,?e? ,φ?P�q?�?�?�?�? O�?+OOOO:OLO�O pO�O�O�O�O�O�O_ '__K_�o_�_�_�_ l��_0_�_�_�_#o
o Go.okoVoho�o�o�o �o�o�o�oC. gR�v���� �	���<�`�* <��`�����ޏ ��)��M�8�q�\��� ����˟���ڟ��� 7�"�[�F�X���|��� |?֯�?�����3�� W�B�{�f�����ÿ�� �������A�,�e� P�uϛ�b_�����Ϫ_ ��߀�=�(�a�s�Z� ��~߻ߦ��������  �9�$�]�H��l�� �����������#�� G�Y� �B�������z� ������
ԏ:�C. gRd����� �	�?*cN �r�����/ ̯&/�M/�q/\/�/ �/�/�/�/�/�/?�/ 7?"?4?m?X?�?|?�? �?�?�?��O!O3O�� WOiO�?�OxO�O�O�O �O�O_�O/__S_>_ P_�_t_�_�_�_�_�_ �_o+ooOo:oso^o �o�op��o�� �� $��o�o�~ �������5�  �Y�D�}�h������� ׏����
�C�.� /v�<���8������ П����?�*�c�N� ��r��������̯� �)��?9�_�q���JO �����ݿȿ��%� 7��[�F��jϣώ� �ϲ�������!��E� 0�i�T�yߟߊ��߮� �߮o�o��o>� t�>��b�������� ���+��O�:�L��� p������������� 'K6oZ�Z� |�~�����5  YDi�z�� ����/
//U/ @/y/@��/�/�/�/�� �/^/???Q?8?u? \?�?�?�?�?�?�?�? OO;O&O8OqO\O�O �O�O�O�O�O�O_�O�7_��$FNO ����VQ��
F0�fQ kP FLAG�8�(LRRM_C�HKTYP  rWP��^P�WP��{QOM�P_MI�N�P����P��  XNPSSB_CFG ?VU ���_���S ooIUTP�_DEF_OW � ��R&hIR�COM�P8o�$G�ENOVRD_D�O�V�6�flTH�R�V d�edkd_�ENBWo k`R�AVC_GRP s1@�WCa X"_ �o_1U<y �r�����	� �-��=�c�J���n� �������ȏ�����;�"�_�F�X���ibR�OU�`FVX�P��&�<b&�8�?��埘���|����  D?��јs���@@g�B��7�p�)�ԙ���`SMT�cG�mM����| �LQHOSTC�Rs1H���P��a�t�SM��f��\���	127�.0��1��  e��ٿ�����ǿ�@�R�d�vϙ�0�*�	�anonymou�s�����������.Q�[�� � ��� ��r����ߨߺ����� -���&�8�[�I�� �������1� C��W�y���`�r��� ���ߺ�������%� c�u�J\n���� �����M�"4 FX��i���� ��7//0/B/T/ ���m/��/�/ �/??,?�/P?b?t? �?�/�?��?�?�?O Oe/w/�/�/�?�O�/ �O�O�O�O�O=?_$_ 6_H_kOY_�?�_�_�_ �_�_'O9OKO]O__Do �Ohozo�o�o�o�O�o �o�o
?o}_Rd v���_�_oo! �Uo*�<�N�`�r��o ������̏ޏ�?Q�&�8�J�\���>�EN�T 1I�� P�!􏪟  �� ��՟ğ�������A� �M�(�v���^����� 㯦��ʯ+�� �a� $���H���l�Ϳ���� �ƿ'��K��o�2� hϥϔ��ό��ϰ�� �����F�k�.ߏ�R� ��v��ߚ��߾���1����U��y�<�QUICC0��b�t���1�����%���2�&���u�!ROUTERv�R�d���!PCJOG�����!192.�168.0.10���w�NAME �!��!ROBO�Tp�S_CFG� 1H�� ��Auto-started�t/FTP��� ���� 2D ��hz����U ��
//./�v�� �/���/�/�/�/ �/�!?3?E?W?i?�/ ?�?�?�?�?�?�?� ��AO�?eO�/�O�O �O�O�?�O�O__+_ NO�OJ_s_�_�_�_�_ 
OO.OoB_'ovOKo ]ooo�oP_>o�o�o�o �oo�o5GYk }�_�_�_��8o ��1�C�U�$y��� �����ӏf���	�� -�?�����Ə�� �ϟ�����;� M�_�q���.�(���˯ ݯ��P�b�t����� m���������ǿٿ�� ���!�3�E�h��{� �ϟϱ����$�6�H� J�/�~�S�e�w߉ߛ� jϿ��������*߬��=�O�a�s��YT_?ERR J5
�����PDUSIZ � ��^J�����>��WRD ?�t��  ?guest}���%�7�I�[�m�$SC�DMNGRP 2�Kt�������V$�K�� �	P01.14� 8��   �y����B  _  ;������ ���������
 �������������~�����C.gR|����  i  ��  
��������� +��������
����l .r���"B�l��� m
d�������_GROuU��L�� ��	����07EQU�PD  	պ��J�TYa �����TTP_AUT�H 1M�� <�!iPenda�ny��6�Y!�KAREL:*8��
-KC///�A/ VISION SETT�/v/�"�/�/�/#�/ �/
??Q?(?:?�?^?�p>�CTRL �N����5�
�.�FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������OYC�R.RDzVTA{��OGBOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G_BUFF 1X�]	��2	աϸ��� ���������!�N� E�W߄�{ߍߺ߱��� �������J����DCS Zr� =����^�+�ZE��������a�IO ;1[
{ ُ!�� �!�1�C�U�i�y� ��������������	 -AQcu��Ы����EfPTM  �d�2/A Sew����� ��//+/=/O/a/�s/�/�/��SEVt����TYP��/??y͒�R�S@"��×�FL 31\
������?��?�?�?�?�?�?/?T�P6��">�NGNAM�ե�U`�7UPS��GI}�����mA_LOAD��G %�%DF_MOTN����O�@MAXUALRM<��J��@sA�QD����WS ��@C �]m�-_���MP2�7�]^
{ ر�	�!+P�+ʠ�;_/�ƅRr�W�_�WU �W�_��R	o�_o?o "ocoNoso�o�o�o�o �o�o�o�o;&K q\�x���� ���#�I�4�m�P� ��|���Ǐ���֏�� !��E�(�i�T�f��� ��ß��ӟ���� � A�,�>�w�Z������� ѯ����د���O� 2�s�^�������Ϳ����ܿ�'��BD_L?DXDISAX@	���MEMO_AP�R@E ?�+
 � *�~ϐϢϴ�����������@ISCw 1_�+ �� IߨT��Q�c�Ϝ߇� �ߧ�����w����>� )�b�t�[����{� ���������:���I� [�/������������ o�����6!ZlS ��s��� �2�AS'�w ����g��./�/R/d/�_MST�R `�-w%SC/D 1am͠L/�/ H/�/�/?�/2??/? h?S?�?w?�?�?�?�? �?
O�?.OORO=OvO aO�O�O�O�O�O�O�O __<_'_L_r_]_�_ �_�_�_�_�_o�_�_ 8o#o\oGo�oko�o�o �o�o�o�o�o"F 1jUg���� �����B�-�f��Q���u�����ҏh/MKCFG b�-�㏕"LTARMu_��cL��� σQ�N�<�M�ETPUI�ǂ����)NDSP_CMNTh���|� ' d�.��ς��ҟܔ|�POSCF�����PSTOL� 1e'�4@�<#�
5�́5�E�S� 1�S�U�g�������߯ ��ӯ���	�K�-�?����c�u�����|�SI�NG_CHK  y��;�ODAQ,��f��Ç��DEV� 	L�	MC}:!�HSIZEh���-��TASK �%6�%$123456789 ������TRIG 1]g�+ l6�%܀��ǃ�����8�p�Y�P[� ��EM_I�NF 1h3�� `)AT&FV0E0"����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ������H�����A���AI�q�,��|����� ���ߵ��� ��J���n������W� ����������"���� X��/����e�� ����0�T; x�=�as�� /�,/c=/b/�/ A/�/�/�/�/��? ���^?p?#/�?�/ �?s?}/�?�?O�?6O HO�/lO?1?C?U?�O y?�O�O3O _�?D_�O�U_z_a_�_�ONIwTOR��G ?5��   	EX�EC1Ƀ�R2�X3��X4�X5�X���V7*�X8�X9Ƀ�RhB Ld�RLd�RLd�RLd
b LdbLd"bLd.bLd:b�LdFbLc2Sh2_h2�kh2wh2�h2�h2��h2�h2�h2�h3�Sh3_h3�R�R_�GRP_SV 1�in���(ͅ�
ߑ3�8��r�mۯ_MOx�_D=R�^��PL_NAM�E !6��p��!Defaul�t Person�ality (f�rom FD) ��RR2eq 1j�)TUX)TX��q��X dϏ8�J� \�n���������ȏڏ ����"�4�F�X�j�|������2'�П� ����*�<�N�`�r��<��������ү� ����,�>�P�b� ȝRdr 1o�y �=\�, �3����� @D�  &��?�����?䰺��A'�6�����;�	lʲ	 ��xJ������ �< �"��� �(pK��K ��K=*��J���J���JV���Z������rτ́p@j��@T;f���f���ұ]�l��I5��p������������b��3��´7  �
`�>�����bϸ�z��Ꝝ�r�Jm��
� B�H�˱]Ӂt�q��	� p�  �P�pQ�p��p|  Ъ�g���c�	'� � ���I� �  �����:�È~
�È=���"��s��	�ВI  ?�n @B�c���\��ۤ��tq�y��rN���  '������@2��@Ǔ����/�C���C�C�@ C�������
��A��  � @<�P�R�
h�B�b�A��j���a��������Dzۀ���߹�����j���( �� -��C���'�7��&����Y������ �?�ff ���gy ������q+q��
>N+�  PƱj�(�� ��7	���|�/?����xZ�p�<
6b<߈�;܍�<�ê�<� <�&Jσ�AI�ɳ+����?fff?I�?y&�k�@�.��J<?�`� q�.�˴fɺ�/�� 5/����j/U/�/y/ �/�/�/�/�/?�/0?q��F�?l??��?/�?+)�?�?�E��� E�I�G+� F��?)O�?�9O_OJO�OnO�Of�BL޳B�?_h�.��O �O��%_�OL_�?m_�?��__�_�_�_�_�
��h�Îg>��_Co�_goRodo�oF�GA�ds�q�C�op�o�o|�����$]Hq���D��fpC���pCHm�ZZ7t���6q�q�����N'�3A�A��AR1AO�^?�$�?�K��0±
=ç>�����3�W
�=�#�W��e��צ�@����{�����<���(�B�u���=B0��?����	L���H�F�G����G��H�U`�E���C�+����I#�I���HD�F���E��RC�j�=��
I���@H�!H�(� E<YD0 q�$��H�3�l�W� ��{��������՟� ��2��V�A�z���w� ����ԯ������� �R�=�v�a������� �����߿��<�'� `�Kτ�oρϺϥ��� �����&��J�\�G� ��kߤߏ��߳����� ��"��F�1�j�U�� y������������0��T�?�Q����(��1��3/E��<���5������M3�8�����M�4Mgs&I�B+2D�a���{�^^	�������uP2P7Q4_A��M0bt��R�������/   � /�b/P/�/t/�/ *�a)_3/�/�/�% 1a?�/?;?M?_?q?  �?�/�?�?�?��?O 2 F��$�vGb�/�A���@�a�`�qC��C@��o�O2���OF�� DzH@�� F?�P D���O�O�ys<O!_3_E_W_�i_s?���@@*pZ.t22!u2~
 p_ �_�_�_	oo-o?oQo couo�o�o�o�o��Q� ��+��1���$MSKCFM�AP  �5� �6�Q�Q�"~�cONREL  
q3�bEXCFENB?wq
s1uXqFNC_�QtJOGOVLI�M?wdIpMrd�bK�EY?w�u�bR�UN�|�u�bS?FSPDTY�av<Ju3sSIGN?Qt�T1MOT�Nq��b_CE_GRP� 1p�5s\ r���j�����T��� �������<��`�� U���M���̟��🧟 �&�ݟJ��C���7� ������گ��������4�V�`TCOM_�CFG 1q}иVp�����
P�_A�RC_\r
jyU?AP_CPL��nt�NOCHECK {?{ 	 r��1�C�U�g�y� �ϝϯ���������	���({NO_WAI�T_L�	uM�NT�X�r{�[m�_7ERRY�2sy3� &�������r��c� ��T_M�O��t��, ��C$�k�3�PARAuM��u{��V`[��!�u?�� =9@�345678901��&���E�W�3� c�����{������� �����=�U�M_RSPACE� �Vv��$OD�RDSP���jxO�FFSET_CAsRTܿ�DIS���PEN_FIL�E� �q��c֮�OPTION_IO���PWORK 5v_�ms �P(�R�@�6$j.j	 ��Hj(6$��p=�_DSBL  �5Js�\��RIENTTO>p9!C��PqfA� �UT_SIM_D�
r�b� V� LCT ww�bc���U)+$_PEXE�d&RATp �vju��p��2X�j)TU�X)TX�##X d-�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O?O�H2�/oO�O�O�O��O�O�O�O�O_]�< ^O;_M___q_�_�_�_ �_�_�_�_o���X��OU[�o(�꘯(���$o��, ��IpB` �@D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	l�mb�`�xJ�`�����a�< ��`��m�a, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�"���� �N	 W��  '!o�:q�pC	 C�@@sBq�|�:�� m�
�!�h@ߐ�n����Z��B	 �A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�����(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��� ��e ���Ӱ��ɆDT� Qy-����D � ��ӱ4�P :� L :�GP:�D :�@ :�U8�8�	8�
8�U8�8�8�8�Q8�X@:�8�8�8�8�8��:�E8�8�x�:�8�PP�:�d :�8�8�P��:�
�:�!8�"8�Q#8���:�%8�&8�U'8�(8�)8�*8�T��:�,8�-8�.8�/8�08�18�,�>� P�b�t���������Ο �����(�:�L�^� p���������L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�(�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_d��_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�_���*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p�������� //$)�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �" |"DEFSPD |�,�!!J �8 IN~ TRL }�-�" 8�(IPE__CONFI� ~g%��g!�$��$�"8 LID�#��-74GRP 1��7Q!�#!A ���&ff"!�A+33D�� �D]� CÀ SA@+6�!�" d�$�9�9*1*0� 	� +9�-+6�? ��	C�?�;B@3AO��?OIO3OmO"!>�?T?�
5�O�O��N�O =��=#�
�O_�O_J_ 5_n_Y_�O}_�_y_�_<�_�_  Dzco" 
oBo�_Roxoco �o�o�o�o�o�o�o�>)bM��;�
V7.10be�ta1�$  �A�E�rӻ�A " �p?!G���q>���r�܁0�q�ͻqBQ��qA\�p�q�4T�q�p�"�BȔ 2�D�V�h�w��p�?�?)2{ȏw�׏ ���4��1�j�U��� y�����֟������ 0��T�?�x�c����� ��ү����!o�,�ۯ P�;�M���q�����ο ���ݿ�(��L�7��p�+9��sF@  �ɣͷϥ�g%����� �+�!6I�[߆����� �ߵߠ���������!� �E�0�B�{�f��� ����������A� ,�e�P���t������� �����=(a L^������ �'9$]�Ϛ� �ϖ�������/ <�5/`�r߄ߖߏ/> �/�/�/�/�/?�/1? ?U?@?R?�?v?�?�? �?�?�?�?O-OOQO <OuO`O�O�O�O�O�� �O_�O)__M_8_q_ \_n_�_�_�_�_�_�_ o�_7oIot���o �o���o�o�o(/! L/^/p/�/{*o�� �������A� ,�e�P�b��������� �Ώ��+�=�(�a� L���p������Oߟ� ��� �9�$�]�H��� l�~�����ۯƯ��� #�No`oro�on��o�o �o�oԿ���8J \ng����vϯϚ� ������	���-��Q� <�u�`�r߫ߖ��ߺ� ������;�M�8�q� \��������z���� ��%��I�4�m�X��� |�����������:� L�^���Z������� ����$�6�H� Swb���� ���//=/(/a/ L/�/p/�/�/�/�/�/ ?�/'??K?]?H?�? ��?�?f?�?�?�?O �?5O OYODO}OhO�O �O�O�O�O�O&8J 4_F_����_�_� �_�_"4-o�O*o coNo�oro�o�o�o�o �o�o)M8q \������� ��7�"�[�m��?�� ��R�Ǐ���֏�!� �E�0�i�T���x��� �����_$_V_ �2��l_~_�_�����R�$�PLID_KNO�W_M  �T������SoV ��U͠�U��
�� .�ǟR�=�O�����m�ӣM_GRP 1���!`0u��T@Rٰo�ҵ�
�� �Pзj��`���!� J�_�W�i�{ύϟϱ����������߱�MR������T��s�w� s��ߠ޴߯߅��� �߻�����A���'� ���������� ����=���#����������}������S��S�T��1 1��U�# ���0�_ A .��,>Pb� �������3 (iL^p��P���2*N���<-/3/)/;/M/4f/x/�/�/5�/�/�/�/A6??(?:?7S?e?w?�?8�?�?�?��?MAD  �d#`PAR�NUM  �w�%OSCH?J �ME
�G`A�Iͣ�EUPD`OrE
a�OT_CMP_��B@�P�@'˥TER_wCHK'U��˪?R$_6[RSl�¯��G_MOA@�_�U_�_~RE_RES_G ��>�oo8o+o \oOo�oso�o�o�o�o��o�o�o�W �\ �_%�Ue Baf�S � ����S0�� ��SR0��#��S�0 >�]�b��S�0}������RV 1�����rB�@c]��t�(�@c\����D�@c[�$���RT?HR_INRl�DA���˥d,�MASS69� ZM�MN8�k��MON_QUEUE ���˦��x�� RDNPUbQN8{�P[��END���_�ڙEXE�ڕ�@B�E�ʟ��OPTI�OǗ�[��PROG�RAM %��%���ۏ�O��TAS�K_IAD0�OCFG ���tO��Š�DATA���Ϋ@��27�>�P�b� t���,�����ɿۿ������#�5�G���IN+FOUӌ������ �ϭϿ��������� +�=�O�a�s߅ߗߩ߀���������^�jč�� yġ?PDI�T �ίc���W�ERFL
��
RGADJ �n�A����?����@�~��IORITY{��QV���MPDSP(H�����Uz����oOTOEy�1�R� (!AF4��E�P]���!t�cph���!u�d��!icm���ݏ6�XY_ȡ�R��ۡ)� a*+/ ۠� W:F�j��� ���%7[�B�*��POR�T#�BC۠�����_CARTRE�P
�R� SKSTyAz��ZSSAV����n�	2500H863���r�$�!�R�����q�n�}/�/�'� UR�GE�B��rYWFF� DO{�rUVWV���$�A�WRUP_�DELAY �|R��$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?�3AQSKIP!�vn�l#x 	1/ +O+ OROdOvO9Hn� �O�G�O�O�O�O�O_ �O_D_V_h_._�_z_ �_�_�_�_�_
o�_.o @oRoovodo�o�o�o �o�o�o�o*<�Lr`���n��?$RCVTM������pDCR!��LЈqCl�f�C��C��>�?�A�>:���<l��4M�b�����O�
�n�������{�4Oi��O� <
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E0�kATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960�iW+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�Ml�P%aR  ��ϰ�P{_��P_INTVAL��@����JR_OPoTION�V �E�BpVAT_GR�P 2�����(y_Ho � e_vo�o�oYo�o�o�o �o�o*<�bOo NDpw����� �	���?�Q�c�u� ����/���ϏᏣ��� �)�;���_�q����� ����O�ɟ���՟ 7�I�[�m�/������� ǯٯ믁��!�3��� C�i�{���O���ÿտ ���ϡ�/�A�S�e� 'ωϛϭ�oρ����� ��+�=���a�s߅� Gߕ߻����ߡ��� '�9�K�]��߁��� ��y����������5��G�Y��E�$SCAN_TIM�AYue�w�R �(ӿ#((�<0.a�aPaP
Tq>��Q��oa�����OOE2/��:	d/"JaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>m�̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:P�_O�UT",REC 1�Z� d �  	 	�������
 �PJ��%6 (�&a�[w�,ݚ*  T J- �- �A�- c| �P�����/ /B/0/f/x/Z/�/�/ �/�/�/�/�/?�/? P?>?t?b?�?�?�?�? �?�?�?OOOLO:O pO�OdO�O�O�O�O�O �O�O$__H_6_X_~_ l_�_�_�_�_�_�_�_  ooDo2oTozo\o�o �o�o�o�o�o�o. R@vd��� �},����4� "�X�F�|���p����� ֏ď����0��@� f�T���x�����ҟ� Ɵ���,��<�b�P� ��h�z������ί� �(�:��^�L�n�p� ������ܿ�п� � 6�$�Z�H�jϐ�rϴ� �����������2�D� &�h�Vߌ�z߰ߞ��� ��������
�@�.�d��R��ZjV 1��w P�m��	�>   y��
TYPEV�FZN_CFGw ��d�7�GRP �1�A�c ,B� A� D;� �B���  B4~RB21/HELL:�(
�� X����%RSR����E 0iT�x��� ���/Se~w�  ��%w�����b#������犍2#�d����H�K 1���  �k/f/x/�/�/�/�/ �/�/�/??C?>?P?�b?�?�?�?�?��OM�M ����?��FTOV_ENB ����+�HOW_RE�G_UIO��IM/WAITB�JK�OUT;F��LIT�IM;E���OV�AL[OMC_UNI�TC�F+�MON_�ALIAS ?e~�9 ( he�� _&_8_J_\_��_�_ �_�_�_j_�_�_oo +o�_Ooaoso�o�oBo �o�o�o�o�o'9 K]n���� t���#�5��Y� k�}�����L�ŏ׏� �����1�C�U�g�� ��������ӟ~���	� �-�?��c�u����� ��V�ϯ������ ;�M�_�q�������� ˿ݿ����%�7�I� ��m�ϑϣϵ�`��� ����ߺ�3�E�W�i� {�&ߟ߱������ߒ� ��/�A�S���w�� ���X�������� ��=�O�a�s���0��� ����������'9 K]����b ���#�GY k}�:���� ��/1/C/U/ /f/ �/�/�/�/l/�/�/	? ?-?�/Q?c?u?�?�? D?�?�?�?�?O�?)O ;OMO_O
O�O�O�O�O �OvO�O__%_7_�C��$SMON_D�EFPRO ����`Q� *SYS�TEM*  d=�OURECALL� ?}`Y ( ��}.xcopy� fr:\*.*� virt:\t�mpback�Q=�>inspiron:6368 �R��_�_�_	o  }/�Ua�_�_�P�_aoso��od
xyzra?te 61 +o=o Oo�o�oe�g�X2112 �o�o] o��o�b+=O�p��)z400���\�n���i3�Ts�:orderfil.dat�l*�ӏ����	�`*�Rmdb:�o*�ˏ\�n��� i�_�o.�O����� o����7�Пa�s��� ����3�N�߯��� (�:�̯]�o������� 9�ʟۿ����$��� H�Y�k�}ϐ�����Ư ������� ���D�Uߘg�yߋ�}6�ϲ�e�mp��192.1�68.4��46:302R�����
��*.d������`�r��1 +�=�O������� ���0� ����c�u����4~ �:prgst�`.dg����U������
�ť�conslog���� ��ew�	io��<N����2��err?all.ls���p�fx� }9�����=S���/}0  ߻��b/t/�/����9R 8144  W/�/�/�/�/�)�/ `?r?�?���;?M?�? �?O�'��4�?�?cO uO�O��5/�'�O�O �O/"/�O�(�Ob_t_`�_����3�=_4 U_8�_�_
o }5 ϱ_ �_�_goyo�o�O�O9_ T_�o�o	_�oEo�o cu��_-o?o�_� ��o��No_�q� ���o�o1�oݏ�� &��J[�m������$SNPX_A�SG 1�������� �PT'%R[1]@1.1����?���%֟�� &�	��\�?�f���u� �������ϯ��"�� F�)�;�|�_������� ֿ��˿���B�%� f�I�[Ϝ�Ϧ��ϵ� ������,��6�b�E� ��i�{߼ߟ������� ����L�/�V��e� ������������ 6��+�l�O�v����� ����������2 V9K�o��� ����&R5 vYk����� /��<//F/r/U/ �/y/�/�/�/�/?�/ &?	??\???f?�?u? �?�?�?�?�?�?"OO FO)O;O|O_O�O�O�O �O�O�O_�O_B_%_ f_I_[_�__�_�_�_ �_�_�_,oo6oboEo �oio{o�o�o�o�o�o �oL/V�e �������� 6��+�l�O�v��������PARAM ���� ��	��P�����OFT_KB_?CFG  ヱ����PIN_SIM  ���C�U��g�����RVQST_P_DSB,���������SR ��/�� & MU�LTIROBOT�TASK������TOP_ON_�ERR  ����PTN z/�@�A	��RING_PRM�� ��VDT_?GRP 1�ˉ�  	�������� ����Я�����*� Q�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߣߠ߲��������� ��0�B�i�f�x�� ������������/� ,�>�P�b�t������� ��������(: L^p����� �� $6HZ �~������ �/ /G/D/V/h/z/ �/�/�/�/�/�/?
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8___�\_��VPRG_CoOUNT��@����RENBU��UM��S��__UPD �1�/�8  
 s_�oo*oSoNo`o ro�o�o�o�o�o�o�o +&8Jsn� �������� "�K�F�X�j������� ��ۏ֏���#��0� B�k�f�x��������� ҟ������C�>�P� b���������ӯί������UYSDE�BUG�P�P�)�d��YH�SP_PAS�S�UB?Z�LOoG ��U�S�)�#�0�  ���Q)�
MC:\x��6���_MPC����U���Qñ8� ��Q�SAV �b����ǲ&�η�SV;�TEM_T�IME 1��[k (m�0&�.:��}YT1SVGUNYS�P�U'�U����ASK_OPTICON�P�U�Q�Q���BCCFG Ì�[u� n�A�a�`a�gZo��߃ߕ� �߹�������:�%� ^�p�[������� �� �����6�!�Z�E��~�i���������&� ������&8��n Y�}�?��ԫ  ��(L:p ^������� / /6/$/F/l/Z/�/ ~/�/�/�/�/�/�/�/ 2?8 F?X?v?�?�? ?�?�?�?�?�?O*O <O
O`ONO�OrO�O�O �O�O�O_�O&__J_ 8_n_\_~_�_�_�_�_ �_�_o�_ o"o4ojo Xo�oD?�o�o�o�o�o xo.TBx� �j������ ��,�b�P���t��� ��Ώ��ޏ��(�� L�:�p�^�������ʟ ��o��6�H�Z� ؟~�l�������د� ��ʯ ��D�2�h�V� x�z���¿���Կ
� ��.��>�d�Rψ�v� �Ϛ��Ͼ�������*� �N��f�xߖߨߺ� 8���������8�J� \�*��n������ ������"��F�4�j� X���|����������� ��0@BT� x�d���� �>,Ntb�� ����/�(// 8/:/L/�/p/�/�/�/ �/�/�/�/$??H?6? l?Z?�?~?�?�?�?�? �?O�&O8OVOhOzO �?�O�O�O�O�O�O
_ _�O@_._d_R_�_v_ �_�_�_�_�_o�_*o oNo<o^o�oro�o�o �o�o�o�o J 8n$O����� X���4�"�X�B��v��$TBCSG_GRP 2�B���  ��v� 
 ?�  ������׏���� ���1��U�g�z����ƈ�d, ����?v�	 HC�=�d�>����e�?CL  B���П�ܘ�����\})��Y  A�ܟf$�B�g�B�Bl��i�X�ɼ���X��  D	J���r�����AC����үܬ���D�@v�=�W�j�}�H� Z���ſ���������v�	V3�.00��	m6;1c�	*X�PĘu�g�p�>���v�(�:�� ��p͟� ; O����p������z�JCFG -�B��� ����+������=��=�c�q�K�q� �߂߻ߦ�������� '��$�]�H��l�� �����������#�� G�2�k�V���z����� ���������p* <N���l��� ����#5GY }h����v� b��>�// /V/D/ z/h/�/�/�/�/�/�/ �/?
?@?.?d?R?t? v?�?�?�?�?�?O�? *OO:O`ONO�OrO�O �O��O�O�O_&__ J_8_n_\_�_�_�_�_ �_�_�_�_�_oFo4o jo|o�o�oZo�o�o�o �o�o�oB0fT �x������ �,��P�>�`�b�t� ����Ώ������� &�L��Od�v���2��� ��ȟʟܟ� �6�$� Z�l�~���N�����د Ư�� �2��B�h� V���z�����Կ¿� ���.��R�@�v�d� �ψϪ��Ͼ������ �<�*�L�N�`ߖ߄� �ߨ����ߚ����� ��\�J��n���� �������"���2�X� F�|�j����������� ����.TBx f������� >,bP�t �����/�(/ /8/:/L/�/�ߚ/�/ �/h/�/�/�/$??H? 6?l?Z?�?�?�?�?�? �?�?O�?ODOVOhO "O4O�O�O�O�O�O�O 
_�O_@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<oro`o�o�o �o�o�o�o�o&�/ >P�/���� �����4�F�X� �(���|�����֏� ���Ə0��@�B�T� ��x�����ҟ����� �,��P�>�t�b��� ������������ :�(�^�L�n������� 2d�����̿�$� Z�H�~�lϢϐ����� ���Ϻ� ��0�2�D� zߌߞ߰�j������� ���
�,�.�@�v�d� ������������ �<�*�`�N���r��� ����������& J\�t��B� �����F4 j|��^���8�/�  2 6#� 6&J/6"�$�TBJOP_GR�P 2����  ?��X,i#�p,� ��xJ� �6$�  �<� �� �6$� @2 �"	 ��C�� �&b  �Cق'�!�!>��1�
559>�0+1��33=�C�L� fff?+0?�ffB� J1�%Y?�d7�.��/>���2\)?0�5����;��hCY�� �  @� �!B�  A�P?�?�3~EC�  D�!8�,�0*BOߦ?�3�JB��
:���Bl�0��0�$�1�?�O6!Aə�A�̔C�1D�G6�=qq�E6O0�p��B��Q�;�A}�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH�1�ts�A@33@?1� C�� �@�_x�_&_8_>��D�U�V_0�LP�Q30<{�zR� @�0�V�P !o3o�_<oRifoPo^o �o�o�oRo�o�o�o�o M(�ol�p~(��p4�6&�q5	V3.00�#�m61c�$*�(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I�R�CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;S@;Q��|8�`rz@/&�8�6&<��1�w�^$�ESTPARS c *({ _#HR��ABLE 1�p+IZ�6#|�Q� � 1�|�|�|�5'=!*|�	|�
|�|�˕�6!|�|�|�N��RDI��z!ʟ@ܟ� ��$���O�������¯ԯ�����S��x# V���˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� U-����ĜP�9�K�]� o��-�?�Q�c�u���~6�NUM  ��z!� >  �Ȑ����_CFG ������!@b IMEBF_TT��p��x#��a�VER���b�w�a�R 1Ξp+
 (3�6"1 ��  6!������ ���� �9�$�:�H�Z� l�~����������������^$��_��@�x�
b MI_CH�ANm� x� kDOBGLV;0o�x��a!n ETHERA�D ?�� ��y�$"�\&n R�OUT��!p*!�*�SNMA�SK�x#�25�5.h�fx^$O�OLOFS_DI�[ՠ	ORQC?TRL �p+;/ ���/+/=/O/a/ s/�/�/�/�/�/��/��/�/!?��PE_D�ETAI��PON_SVOFF��33P_MON ��H�v�2-9STRTCHK ����42VTCOM�PATa8�24:0FPROG %��%MULTIROBOTTO!O06��PLAY��L:_�INST_MP 2GL7YDUS���?��2LCK�LPKQUICKMEt �O�2oSCRE�@�
tps��2�A�@�I��@_Y���9��	SR_GRP �1�� ���\�l_zZg_�_�_�_�_�_�^�^�oj �Q'ODo/ohoSe��o o�o�o�o�o�o�o !WE{i�������	1234567��!�ڎ�X�E1�V[
 ��}ipnl/�a�gen.htm�no��������ȏ~��Panel s/etup̌}�?�`�0�B�T�f� �� 񏞟��ԟ���o� ���@�R�d�v����� �#�Я�����*� ��ϯůr��������� ̿C��g��&�8�J� \�n�����϶����� ����uϣϙ�F�X�j� |ߎߠ����;��������0�B��*NUA�LRMb@G ?�� [������ ������ ��%�C�I��z�m�������v�SEoV  �����t�ECFG �Ё=]/BaA$  w B�/D
 �� /C�Wi{��� ���� PRց; �To\o�eI�6?K0(%�� ��0�����/ /;/&/L/q/\/�/�/�/l�D �Q�/�I_�@HIST �1ׁ9  (��0 ��(/S�OFTPART/�GENLINK?�current=�menupage,153,1 E�c0p?�?�?�?/C�'=?O>71n?�?	OO�-O�13�?O5edi�t[2MULTIR`f?O�O�O2O� FOP=962vO __$_06_�O�O�A36�O�_ �_�_�_IR�_�_�_o o+o=o�_aoso�o�o �o�oJo�o�o'9I|��a81�ou� �����o��� )�;�M��q������� ��ˏZ�l���%�7� I�[���������ǟ ٟh����!�3�E�W� ���������ïկ� v���/�A�S�e�P b������ѿ����� �+�=�O�a�s�ϗ� �ϻ�������ߒ�'� 9�K�]�o߁�ߥ߷� �������ߎ�#�5�G� Y�k�}�������� �������1�C�U�g� y���v����������� 	�?Qcu� �(���� )�M_q��� 6���//%/� I/[/m//�/�/�/D/ �/�/�/?!?3?�/W? i?{?�?�?�?�����? �?OO/OAOD?eOwO �O�O�O�ONO`O�O_ _+_=_O_�Os_�_�_ �_�_�_\_�_oo'o 9oKo�_�_�o�o�o�o �o�ojo�o#5G Y�o}�������?��$UI_P�ANEDATA �1������  	�}�0�B�T�f�x��� )�����4�ۏ� ���#�5���Y�@�}� ��v�����ן����� ��1��U�g�N������ �1��Ïȯ گ����"�u�F��� X�|�������Ŀֿ=� �����0�T�;�x� _ϜϮϕ��Ϲ������,ߟ�M��j�o� �ߓߥ߷������`� �#�5�G�Y�k��ߏ� ������������� �C�*�g�y�`����� ����F�X�	-? Qc����߫�� ��~;"_ F��|���� �/�7/I/0/m/�� ���/�/�/�/�/�/P/ !?3?�W?i?{?�?�? �??�?�?�?O�?/O OSOeOLO�OpO�O�O �O�O�O_z/�/J?O_ a_s_�_�_�_�O�_@? �_oo'o9oKo�_oo �oho�o�o�o�o�o�o �o#
GY@}d ��&_8_���� 1�C��g��_������ ��ӏ���^���?� &�c�u�\�������ϟ ���ڟ�)��M�� ���������˯ݯ0� ����7�I�[�m�� ��������ٿ�ҿ� ��3�E�,�i�Pύϟ�����Ϫ���Z�l�}����1�C�U�g�yߋ�) ߰�#������� �� $�6��Z�A�~�e�w� �����������2� �V�h�O����v�p���$UI_PAN�ELINK 1��v�  ��  ��}�1234567890����	-? G���o���� �a��#5GD�	����p&���  R����� Z��$/6/H/Z/l/ ~//�/�/�/�/�/�/ �/
?2?D?V?h?z?? $?�?�?�?�?�?
O�? .O@OROdOvO�O O�O �O�O�O�O_�O�O<_�N_`_r_�_�_�0, ���_��_�_�_ o2o oVohoKo�ooo�o�o �o�o�o�o��, >r}������� �����/�A�S� e�w��������я� ��tv�z����=� O�a�s�������0S�� ӟ���	��-���Q� c�u�������:�ϯ� ���)���M�_�q� ��������H�ݿ�� �%�7�ƿ[�m�ϑ� �ϵ�D��������!� 3�Eߴ_i�{�
�߂� ���߸������/�� S�e�H���~��R~ '�'�a��:�L�^� p���������������  ��6HZl~ ���#�5���  2D��hz�� ���c�
//./ @/R/�v/�/�/�/�/ �/_/�/??*?<?N? `?�/�?�?�?�?�?�? m?OO&O8OJO\O�? �O�O�O�O�O�O�O[� _��4_F_)_j_|___ �_�_�_�_�_�_o�_ 0ooTofo��o��o ��o�o�o,> 1bt����K ����(�:��� �{O������ʏ܏� uO�$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v�������� п���ϕ�*�<�N� `�rτ��O�Ϻ�Io�� �������8�J�-�n� ��cߤ߇����߽��� �o1�oX��o|�� ������������ 0�B�T�f�������� ������S�e�w�,> Pbt��'�� ���:L^ p��#����  //$/�H/Z/l/~/ �/�/1/�/�/�/�/?  ?�/D?V?h?z?�?�? �???�?�?�?
OO.O ��ROdO�߈OkO�O�O �O�O�O�O_�O<_N_ 1_r_�_g_�_7O�M�m�$UI_Q�UICKMEN � ���_AobRESTO�RE 1��  � |��Rto�o�im�o�o �o�o�o:L^ p�%����� �o����Z�l�~� ����E�Ə؏����  �ÏD�V�h�z���7� ������/���
��.� @��d�v�������O� Я�����ßͯ7� I���m�������̿޿ ����&�8�J��n� �ϒϤ϶�a������� Y�"�4�F�X�j�ߎ� �߲������ߋ����0�B�T�gSCRE�`?#muw1sco`u2��U3��4��5��6���7��8��bUSE�Rq�v��Tp���k�s����4��5��6���7��8��`ND�O_CFG ܶ#k  n` `P�DATE ���Noneb�SEUFRAME�  �TA�n�R�TOL_ABRT8y�l��ENB����?GRP 1�ci/aCz  A��� ��Q�� $6H!Rd��`U����~��MSK  ��4���Nv�%�U��%���bVISCAND_MAX��I��FAI�L_IMG� �P��P#��IMRE/GNUM�
,[gSIZ�n`�A��,VONTMOiU��@����2��a��a�����FR:�\ � �MC:\�\LO�G�B@F� !��'/!+/O/�Uz? MCV�8#oUD1r&EX{+�S�PPO64�_��0'fn66PO��LIb�*��#V���,f@��'�/� =	�(S�ZV�.����'W�AI�/STAT' ����P@/�?��?�:$�?�?��2�DWP  ���P G@+b=���� H�O_JMPERR 1�#k�
  �2345?678901dF�� �O{O�O�O�O�O�O_ �O*__N_A_S_�_
� MLOWc>
 ��_TI�=�'�MPHASE � ��F��PSoHIFT�1 9�]@<�\�Do�U #oIo�oYoko�o�o�o �o�o�o�o6l CU�y���� � ��	�V�-�e2�����	VSFT]1�2	VM��� �5�1G� ���~%A�  B8̀̀�@ pكӁ˂1�у��z�ME@��?�{��!c>&%�JaM1��k�0�{ ��$`0TDINE#ND��\�O� �z����S��w��P����ϜRELE��Q��Y���\�_ACTIV��:�R�A ��e���e��:�RD� ���YBOX �9�د�6���02���190.0.��83��25�4��QF�	 ��X�j��1��robot��� ?  p�૿�5pc��̿������7�����-�f�ZWABC�����,]@ U��2ʿ�eϢωϛ� �Ͽ����� ���V�@=�z�a�s߰�E�Z��1�Ѧ