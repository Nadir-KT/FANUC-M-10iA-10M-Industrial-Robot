��   ��A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���D�RYRUN_T   � $'�ENB  $�NUM_PORT�A ESU@$STATE P _TCOL_��PM�PMCmGRP_�MASKZE� O�TIONNLOG�_INFONiA�VcFLTR_E�MPTYd $P�ROD__ L �  � &J_  �4 $TYPE�NFST_IDX���_ICI�M_IX_BG-��� G_NAMc �%$MODc_U�SdCIFY_T�I<  $MK�R-  $�LINc   x_SIZc"� �.  $USE_FLGA�l�i�SIM�A�Q�QB�S�CANRAX�I�N�I��_COU�NrRO�_!_?TMR_VA�gyh>�i� p'` ���H�!^%��$$CLASS  ����!���5��5� VIRTUR �/� '/ �%_5�������8� �!2,�%I1�+�M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO���+6W?�%�! ���O�OV�O  10� �' 1�+ 4%zO*_��11_ ]_<_�_�_r_�_�_�_ �_�_�_#oooYo8o Jo�ono1�C���-54�� �b1�d,1�!�a�o. @Rdv���� ���?~c�a1&� 8�J�\�n��������� ȏڏ�����!�C��1�)  U�g�y��������� ӟ���	��-��G� `�r���������̯ޯ ���&�8�C�\�n� ��������ȿڿ��� �"�4�F�Q�j�|ώ� �ϲ����������� 0�B�M�_�xߊߜ߮� ����������,�>� P�[�t������� ������(�:�L�^� i��������������  $6HZe�w� �������  2DVh�F