��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  �(��ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1��  |UREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|~GRG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"�SB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5� UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COMW!2MO� 21� A�.	 \rVE��1$F�RA{�$O�UDcB]CTM�P1_FtE2}G1Q_�3�B�2�X�D�#
 d �$CARD_EX�IST4$FS?SB_TYP!A?HKBD_SNB�1�AGN Gn �$SLOT_NUyM�APREV4DEBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP��U0LETE_OK��BUS�P_CR��A$;4AV� 0LACIw1�R�@�k �1$@MEN�@$D�V�Q`PvVA�{G BL� OU&R ,A�0�!z� B� LM_O�z
eR�"CAM_;�1 xr$�ATTR4�@� A�NNN@5IMG_�HEIGH�AXcWoIDTH4VT� ��UU0F_ASP�EC�A$M�0E�XP�.@AX�f��CF�D X '$GR� � S�!.@=B�PNFLI�`�d� UIRE 3T!GOITCH+C�`N� MS�d_LZ`AC�"��`EDp�dL� J�4S�0� <za�!p�;G0 � 
?$WARNM�0f�!�@� -s�pNST�� CORN�"a1F�LTR{uTRAT�� T}p  $ACCa1�p��|{��rORI�P�C�kR�T0_S~BG CHuG,I1 [ �T�`�"3I�pTYP4D�@*2 3`#@�� �!�B*HDDcJ�* Cd�2_�3_�4�_�5_�6_�7_�8�_�94�ACO�$ <� �o�o�hK3 1�#`O_Mc@AC �t � E#6NGPvABA� �c1�@Q8��`,��@nr1�� d�P�0e���axnpUP&Pb26h���p�"J�p_R�r�PBC��J�rĘߜJV�@U� B��s}�g1��"YtP_*0OFS�&R @� RO_�K8T��aIT�3T�N'OM_�0�1p�384 >��D �� Ќd@��hPV��mEX�p�� �0g0ۤ�p�r
�$TF�2C$MDM3i�TO�3�0U� ^F� ��Hw2JtC1(�Ez�g0#E�{"F�"F�40CPh@�a2 �@$�P�PU�3N)�ύRևAX�!DU���AI�3BUFp�F=�@1 |pp����pPIT� PP�M�M�y��}F�SIMQSI��"ܢVAڤT���x T�`(zM��P�B^�qFACTb�@EW�P1�BTv?��MC� �$�*1JB`p�*1DE�C��F��Ž�Ԁ�� �H0CHNS�_EMP1�$G��8��@_4�3�p|@P��3�TCc�(r/� 0-sx��ܐ� MBi���!����JR� i�S/EGFR��Iv �a�R�TpN�C��P�VF4�+cw &��f{uJc!� Ja��� !28�ץ�AJ���SIZ�3S�c�B��TM���g��JaRSINFȑb���q�� ��н����L�3��B���CRC�e�3CCp����c��mc� �b�1J�cѿ�.����D$ICb�Cq�5r��`���@v�'���EV����zF��_��F,pN��ܫ�?�4�0A�! �r���h�� ���p�2�͕a�� ��دp�R�Dx Ϗ��o"27�!A�RV�O`C�$LG�pV�B�1�P��@�tB�aA�0'�|�+0Ro�� MEp`"1 CfRA 3 AZV�hg6p�O �FCCb�`�`F�`K������ADI��a�A�b A'�.p��p�`�c�`aS4PƑ�a�AMP�Ԓ-`Y�3P�M�]pUtR��QUA1  $@TITO1/S@S�!�����"0�DBPX�WO��B0!5�$�SK���28@DBdq�!"�"�PR�� 
� =����!#� S q1$2�)$z���L�)$�/�ä�� %�/�$C�!&�?�$ENE�q.1'*?�Ú RE�p2_(H ��O�0o#$L|3$$�#��B[�;���FO_9D��ROSr��#������3RIGGER�6PApS���ҟETURN�2�cM[R_8�TUw��0EWM��M�G1N�P���BLAH�<E��P��&$PD� �'P@T�3�CkD{��DQ���4�11���FGO_AWAY��BMO�ѱQ#!��DCS_�)  �PIS� I g�b {s�C��A��[  �B$�S��AbP�@�E9W-�TNTVճ�BV�Q.�C�(c`�UWr��P�J��P�$0��SAsFE���V_SV�b�EXCLU��NnONL<зSY��*a&�OT�a'�HI�_V�4��B���_G *P0� 9�_z���p ��ASG�� +nrr�@6A@cc*b��G�#@E�V.i|Hb?fANNUN$0,.$fdID�U�2�SC@�`�i�a��j�fQ��z��@I$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6r�!MS�W�E. 8Q�KE3YI5���TM�10s�qA�vIN��#�b���/ D��HOST_P!�rT��t�a��tn��tsp�pEMpӰV��� SBLc �ULI�0  p8	=ȳ�r�DTk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&Q�DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F��df�J� ���aC1+�6 H�bLL_DUs�~a3@{��3:���OTX"���s��r�0NOAUTO�!7�p$)�$�*�R�c4�(�C� 8��C, �""�L�� �8H *8�L H <6����c"�`,  `Ĭ�kª�q��q��Psq��~q��7��8���9��0����1��1�̺1ٺ1�1�1� �1�1�2(�2T����2̺2ٺ2�U2�2 �2�2ʕ3(�3��3��̺3�ٺ3�3�3 �3
�3�4(�ɢT�?��!9 <�9�&�z���I��1���M��QFqE@'@� : ,6���Q? �@P?Q9��5�9�E�@DA�- ��A� ;p�$TP�$V7ARI:��\���7UP2�P< ���TDe���K`Q��r��ፁBAC�"G= T�p��e$)_,p�bn�kp+ IFIG�kp�H  ��P���@`�!>t� ;E��sC�ST�D� D���c�<� 	C��{��_����l���R  ���F?ORCEUP?b���FLUS�`H�N�>�F ���RD_CM�@E������ ��@v\MP��REMr F�Q���1k@���7Q
Kr4	NJ�5EFFۓ�:�@IN2Q��OV�O�OVA�	TR3OV���DTՀ�DTMX� ��@ �
ے_PH"p��CL��_TpE�@�p2K	_(�Y_T��v*(��@A;QD� ������!0tܑ0RQ���_�a����M�7�CL�dρR�IV'�{��EAR6ۑIOHPC�@��2��B�B��CM9@����R �GCLF�e!DYk(M�ap#5TuDG��� :�%��`FSSD �s�? P�a�!�1����P_�!�(�!1��E��3�!3�+5�&�GSRA��7�@��;ᚔPW��ONn��EBUG_SD2H�P�{�_E A`|ꁣ��TERM`5�Bi5E��OR�I#e0C�9SM_h�P��e0D�9TA�9�Ei5aUP\�Fg� -�A{�AdP|w3S@B$SEG�:v� EL{UUSE�@NFIJ�B$�;1x젎4�4C$UFlP=�$,�|QR@��_G90Tk�D�~SwNST�PAT��<��APTHJ��E�p%B`�'EC����AR$P�I�aS�HFTy�A�A�H_�SHORР꣦6 ��0$�7PE��E�O#VR=��aPI�@��U�b �QAYLOW���IE"�r�A��?���ERV��XQ� Y��mG>@�BN��U�\��R2!P.uAScYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC���EaP;�uP;�6WOR>@�M`�!�GRSMT6�G3�GR��13�a�PAL@��p�q�uH� � ���T�OCA�`P	P�`$OP����p�ѡ��`0O��RE�`R4C�AO�p낎Be�`R�Eu�h�A���e$PWR�IMu�RR_�cN��q.=B I&2H���p�_ADDR��H_LENG�B�q�q�qVˠRR��S�JڢSS��SKN��u\�0�u̳�uٳSE�A��jrS��MN�!K������b����O�LX��p����`ACRO3pJ�@��X��+��Q��6�OUP3�b_�IX��a�a1��}򚃳���(�� H��D��ٰ��氋�VIO2S�D������	�7�L $xd��`Y!_OFFr��PRM_��ӾʠHTTP_+�H�:�M (|pOBJ�]"�p��$��LE�~Cd���N � ���֑AB_�T�qᶔS�`H�LV�h�KR"uHIT�COU��BG�LO�q���h�����`��`SS� ����HW�#A:�Oڠ�<`INCPU2VISIOW�͑��n���to��to�ٲ �IwOLN��P 8��yR��p$SLob� PUT_n�	$p��P& ¢��Y �F_AS�"Q���$L������Q  U�0	P4A��^���ZP#HY��-��y��sUOI �#R `� K����$�u�"pPpk���$�������2J5�S-���NE�6WJOGKG̲DI�S���Kp���#T� (�uAVF�+`�C�TR�C
�FLAG�2�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w�  m�_�{0a�^��cg��� 4�����Ǝ���{0��� SCH_���a7��N�9�VW���E �"����4��UM�A�r�`LJ�@�DAUfՃEAU�p��d|�r�GqH�b����BOO��WL ?�6 I�T��Y��REC���SCR ܓ�Dx
�\���MARGm� !��զ ��d%�����	S����W���U� ��JGM[�MNCH|J���FNKEY\��K��PRG��UF���7P��FWD��H]L��STP��V��=@��А�RS��HO`����C9T��b ��7�[�UL���6�(R�D� ����Gt��@P�O��������MD�F�OCU��RGEX.��TUI��I��4�@�L�����P����`��P��NE��CANA��Bj�oVAILI�CL !~�UDCS_HII4���s�O�(!�S���S��D����BUFF�!X�?PTH$m���vP`���1��AtrY��?P��j�3��`OS1Z2Z3Z8�>� Z � ��[apEȤ��ȤIDX�d	PSRrO���zA�+STL�R}�Y&��� Y$E�C ���K�&&���ѿ![ LQ��+00�	P ���`#qdt
�U�dw<�~��_ \ ?�@4Г�\��Ѩ#\0C4��] ��CLDP|L��UTRQLI��pdڰ�)�$FLG&�� 1�#�D���'B��LD�%�$�%ORG ڰ5�2�PVŇVY8�sp�T�r�$}d^ ��P�$6��$�%S�`T� ��B0�4�6RCLMC�4]?o?�9세�sMI�p}d_ d=�֚RQ��DS3TB�p� ;F�6HHAX�R JHdLEXCESr��B)M!p�a`��/B�T��b�B��`a�p=F_A7Ji��KbOtH:� K�db \Q��n�v$MBC�LI|�~)SREQUIR�R��a.\o�AXDEBUTZ�ALt M��c�b��{P����2ANDRѧ`�`d;�2��f�SDC��N�INl� K�x`��X� N&��apZ��D��RPST�w ezrLOC��RIrp�EX<fA�p�9AAODAQn��f XY�OND�rMF,Łf�s"���}%�e/� �1!FX�3@IGG�� g ��t"��ܓs#N�s$R�a%��iL���hL�v�@�DAT	A#?pE�%�tR���Y�Nh t W$MD`qI}�)nv� ytq�ytHP`�Pxux��(�zsANSW)�Pyt@��yuD+�)\b����0o�i �@C�Uw�V�p 0XeRR2��j Du�{Q��~7Bd$CALIA@���G��2��RI�N��"�<E�NTE��Ck�r^�آXb]���_N�qlk���9��D���Bm��DIVFFDH�@���qnI�$V,��S�$��$Z�X�o��*����oH ?�$BELT�u!_ACCEL�.�~�=�IRC�� ����D�T�8�$PS�@�"L���r��#�^�S�Eы T�PAT!H3���I���3x�p�A_W��ڐ���2n�C��4�_MG��$DD��T���$FW�Rp9��I�4���DE7�PPAB�N��ROTSPE!E�[g�� J��[��C@4���$US�E_+�VPi��S�YY���1 �aYNr!@A�ǦOFF�qnǡMOU��NGL����OL����INC �tMa6��HB��0HBENCS+�8q9Bp�X4�FDm�IN�Ix�0]��B��VE��#�>y�23_UP񕋳/LOWL���p� B���Du�9B#P`��x ���BCv�r�MO3SI��BMOU��@��7PERCH  ȳOV��â
ǝ� ���D�ScF�@MP����� Vݡ�@y�j��LUk��Gj�p�UPp=ó���ĶTRK�>�AYLOA�Qe� �A��x�����N`�F��RTI�A$��MO UІ�HB�BS0�p7D5����ë�Z�DU�M2ԓS_BCKLSH_Cx�k�� ��ϣ���=���ޡ< �	ACLAL"q�p�1м@��CHK� :�S�RTY���^�%E1Qq_�޴_�UM�@�C#��S�CL0�r�LMT_OJ1_L��9@H��qU�EO�p�b�_�e�k�e�SPC��u�L��N�PC�N�Hz �\P��C�0~"XT\��CN_:�N9�L�I�SF!�?�V����U�/���x�T���CB!�SH�:��E� E1T�T����y���T�f�PA ��_P��_� =������!����J6 L�@���OG�G�TORQU��ONֹ��E�R0��H�E�g_W2��ā_郅���I*�I�I��Ff`xaJ�1�~1�VC3�0BD:B�1�@SBJRKF9~�0DBL_SM�:�2M�P_DL2GRV�����fH_��d���CcOS���LNH ��������!*,�aZ���fcMY�_(�TH���)THET0��N�K23���"��C-B�&CB�CAA�B��"��!��!�&SB8� 2�%GTS�Ar�CIMa�����,4#<97#$DU���H�\1� �:Bk62�:AQ�(rSf$NE�D�`I ��B+5��$̀�!�A�%�5�7���LCPH�E�2���2S C%C%�2-&FC0JM&̀V�8V�8߀LUVJV!KV/KV=KUVKKVYKVgIH�8@FRM��#X!KH/KUH=KHKKHYKHgI�O�<O�8O�YNO�JO!KO/KO=KO*KKOYKOM&F�2�!�+i%0d�7SPBA?LANCE_o![c�LE0H_�%SP�c� &�b&�b&PFULC�h�b�g�b%�p�1k%�UTO_<��T1T2�i/�2N��"�{�t#�Ѡ�`�0�*�.�T��O�À<�v INSEG"�ͱREV4vͰl�gDIF�ŕ�1lzw6��1m��OBpq�ь�?�MI{���nL�CHWARY�_�A�B��!�$MEC�H�!o ��q�AX���P����7Ђ�`n� 
�d(�U�RO�B��CRr�H����(�MSK_f`��p P �`_���R/�k�z�����1 S�~�|�z�{���z��q�INUq�MTC�OM_C� �q � ���pO�$ONOREn����p�Ђr 8p GRle�uSDZ�AB��$XYZ_DAx�1a���DEBUUqX������s z`$��wCOD�� L����p�$BU�FINDX|� � <�MORm�t $فUA��֐�Р�r�<��rG��u� � $SIMUL  S�*�Y�̑a��OBJE�`̖AD�JUS�ݐAY_	IS�D�3���_FI�=��T u 7�~�6�'��p} =��C�}p�@b�D��FRiIr��T��RO@ �\�E}'�y�OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1���e��M��ED}�*�p ��N�PMֲ����c�w�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B�P2�G�B�_�M����q�E� x Hxw��p��ATUSWЅ��C�0o�s���BSTM�ǌ�I�k��4��x�԰q�y DBw�E&���@E�r���7��жЗ�EXE ��ἱ�����f q�gz @w���UP'�f�$�pQ�XN����������� �P�G΅{ h $GSUB����0_��|�!�MPWAIv�P7ã�LOR�٠F�\p˕$RCVF�AIL_C��٠B�WD΁�v�DEF�SP!p | L�w���Я�\���UCNI+�����H�R�,+�}_L\pP��x�t���p�}H�> �*��j�(�s`~�N�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��G���PLI��p� � $ˀP_S�WI�pq�J_PL~��AL_ ���J��A��B��� C���D�$E���.�C_�U�� � � ���*��J3K0����TIA�4��5��6��MOM��������ˀB��AD��������6��PU� NR��������m��?� A$PI�6q� �	�����K4��)6�U��w`��SPEEDgPG���� ����Ի�4T�� �� @��SAM�r`��\�]��MOV_�_$�npt5��5$���1���2���� ����'�S�Hp�IN�'�@�+�����4($4+T+GA�MMWf�1'�$G#ET`�p���Da���=

pLIBR>�I]I2�$HI=�_g�Ht��2�&E;��(A�.� �&LW�-6<�)@56�&]��v�p��V���$PDCK����q��_?���� �q�&���7��4����9+� �$I/M_SR�pD�s�r�F��r�rLE���O0m0H]��0�-�p�q��PJqUR_�SCRN�FA���S_SAVE_D��,dE@�NOa�CAA� b�d@�$q�Z�Iǡs	 �I� �J�K� ����H �L��>�"hq�� ����ɢ�� bWP^US�Aѩ��M4���a��)q`��3�W@W�I@v�_�=���MUA�o�� � $P9Y+�$W�P�vNG�{��P:��RA�0�RH��RO�PL������q� ��s'�X;�O�I�&�Zxe ���m��# p��ˀ�3s�O@�O�O�O�O�aa�_т� |��q�d@��.v ��.v��d@��[wFv��AE���%s�t;B�w��|�tP���PMvA�QUa ��qQ8��1٠QTH��HOLG�QHYSf��ES��qUE�ptZB��Oτ�  ـPܐ(�A����v�!�%t�O`�q��u�"�p��FA��IROG�����Q2���o�"���p��INFOҁ��׃V����R�H�OI� (�0SLEQ������Y�3���$�Á��P0Ow0�j��!E0NU���AUT�A�CO�PY�=�/�'��@Mg�N��=�}1������M ��RG��Á���3X_�P�$;ख�`��W��P��@��������EXT_CYC bHᝡRpÁ��r��_NAe1!А���ROv`	�?� � ��ЇPOR_�1�E2�S�RV �)_�I�DI��T_�k�}�'���PdЇ�����5��6��%7��8i�H�SdB��-�2�$��F�p���GPLeAdA
�TAR�Б@���P��2�裔d� ,�0F1L`�o@YN��K��M��Ck��PWR�+�9ᘐ��DELiA}�dY�pAD�a�� �QSKIPN4� �A�$�OB`�NT�} ��P_ $�M�ƷF@\br ݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q����TQ������ ���`�#�RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�dG�REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"�������2�Қ�߼��߸����� R��3�қ'�9�K�]�o��
�4�Ҝ�������(�����5�ҝ!�3��E�W�i�{��6�Ҟ��������������7�ҟ-?Qcu
�8�Ҡ����x���SMSKÁ%�l��a��EkA��oMOTE6������@�݂TQ�IO�}5�ISTP��PO9W@��� �pJ� ���p����E�"�$DSB_SIG!N�1UQ�x�C\��/S232���R�i�DEVICEUS��XRSRPARIT|��4!OPBIT�Q�I�OWCONT�R+�TQ��?SRCU�� MpSUXTAS�K�3N�p�0p$TA�TU�P�qRS��0�����p_XPC�)�$FREEF�ROMS	pna�GsET�0��UPD��A�2�#P� :���� !$US�AN�na&����ER1I�0�RpRYq5*"�_j@�Pm1�!�6WRK9KD���6��~QFRIEND�Q��RUFg�҃�0TO�OL�6MY�t$�LENGTH_VT\�FIR�pC�@�ˀE> +IUFINt-RM��RGI�1�ÐAITI�$GX�ñ3IvFG2v7G1`���p3�B�GPR�p�1F�O_n 0��!�RE��p�53҅U�T�C��3A�A�F �G((��":���e1n! ��J�8�%���%]���%�� 74�X TO0�L��T�3H&���8���%b453GE�W$�0�WsR�TD�����T��M����Q�T]�=$V 2����1��а91�8�02�;2
k3�;3�:ifa�9�-i�aQ��NS��ZR$)V��2BVwEV�2AQUQ�B;�����& �S�`��F�"�k�@�2�a�PS�E��$pr1C��_$Aܠ�6wPR��7vMU�cS��t '�/89�� 0�G�aV`��p�d`����50�@��-�
25S^�� ��aRW�����B�&�N�A)X�!�A:@LAh�^�rTHIC�1I�8��X�d1TFEj��q>�uIF_CH�3�qaI܇7�Q�pG1Rx�V���]��:�u�_�JF~�PRԀƱ��RVAT��� ���`���0RҦ�DO�fE��COUԱ��A�XI���OFFS=E׆TRIGNS����c����h�����Hx�Y��IGMA0�PA�pJ�E�ORG�_UNEV�J� ��S�����d ӎ$CА�J�GR3OU����TOށ�!DSP��JOG�Ӑ�#��_Pӱ�"O��q����@�&KEPF�IR��ܔ�@M}R&��AP�Q^�Eh0��K�SYS�q"K�;PG2�BRK�B��߄�pY�=�d�����`AD_�����BS�OC���N��DU�MMY14�p�0S}V�PDE_OP�#�SFSPD_OVR-���C��ˢΓ�OR٧3N]0ڦF��ڦ��OV��SF��p���F+�r!���CC��1q"LCHD}L��RECOVʤc0��Wq@M������#RO�#��Ȑ_+���� @0�e@VER��$OFSe@CV/ �2WD�}���Z2���TR�!|���E_FDO��MB_CM���B��BL�bܒ#��adt�VQR�$0p���G$�7�AM5��� e����_M;��"'����8$CA��'�E�>8�8$HBK(1���IO<�����QPPA������
���������DVC_DBhC;��#"<Ѝ�r!"S�1[ڤ�S�3[֪�/ATIOq 1q� �ʡU�3���CAB Ő�2�CvP��9P^�B��_� �SUBCPU�ƐS�P � M�)0NS�cM�"r�?$HW_C��U���S@��SA�A�pl$�UNITm�l_�A�T���e�ƐCYC=Lq�NECA����FLTR_2_F�IO�7(��)&B�LPxқ/�.�_SCT�CF_`�Fb�l���|��FS(!E�e�CHA��1��4�D°"3�RS�D��$"}����_Tb�PRO����� KEMi_��a�8!�a !�a��D�IR0�RAILAiCI���Mr�LO��C���Qq��#q��V��PR=�S�A�p�C/�c 	��FUsNCq�0rRINP`�Q�0��2�!RAC �B ��[���[gWARn���BL�A�q�A����D�Ak�\���LD@0���Q��qeq�TI"r��K�hPgRIA�!r"AF��Pz!=�;��?,`�R�K���MǀI�!�D�F_@B�%1n�LM��FAq@HRDY4�4_�P@RS�A�0|� �MULSE@x���a ���ưt��m�$�1-$�1$1o������ x*�EaGE ����!AR���Ӧ�09�2,%� 7�wAXE��ROB���WpA��_l-��SY�[�W!‎&S�'WR�U�/-1��@�STRП�����Eb� !	�%��J��AB� ����&9�����OTo0v 	$��ARY�s�#2��Ԓ�	ёFI�@��$LINK(|�qC1�a_�#����%kqj2XYZ@��t;rq�3�C1j2J^8'0B��'�40����+ �3FI���7`�q����'��_Jˑp���O3�QOP_�$2;5���ATBA�2QBC��&�DUβ�&=6��TURN߁"r��E11:�p��9GFL��`_���* �@�5�*7���Ʊ 1�� KŐM��&8���"r��ORQ��a �(@#p=�j�g�#qXUp�����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb��T {�, ��@;�uQ���P \�i��UuQ�We�eL�SERʑe	��!E� O���UdAas���4S�/7����AX��B�'q��E1�e ��i��irp�jJ@�j �@�j�@�jP�j@ �j �!�f��i��i��i ��i��i�y�y��'y�7yTqHyDEBU8�$32����qͲf2G + AB�����رnSVS�7� 
#�d��L�#�L� �1W��1W�JAW��AW� �AW�QW�@!E@?\D2�3LAB�29U�4�Aӏ��C  �o�ERf�5� �� $�@_ A��!�PO��à�0#��
�_MRAt�� �d � T��ٔEcRR����;TY&����I��V�0�cz�TOQ�d�PL[ �d�"ҍ�	��C! � pp`T)0���_V1Vr�aӔ�����2ٛ2�E����@�8H�E���$W���j��V!��$�P@��o�cI��aΣ	 �HELL_CFG�!� 5��Bo_BASq�SR3�\�� a#Sb�T��1�%��2��U3��4��5��6��e7��8���RO�����I0�0NL�\CAqB+�����ACK4� ����,�\@2@�&�?�7_PU�CO. U�OUG�P~ ����m�ذ�����TPհ_KcAR�l�_�RE*��P���7QUE����uP����CST?OPI_AL7�l��k0��h��]�l0SE�M�4�(�M4�6�T�YN�SO���DI�Z�~�A�����m_T}M�MANRQ���k0E����$KEYSWITCH��ص�m���HE��BE�AT��E- LE(~�����U��F!Ĳ�|��B�O_HOM=�OGREFUPPR�&��y!� [�C��O��-ECOC��Ԯ0_IOCMWD
�a��{(k��� �# Dh1���UX����M�βgPgCFOR�C�����OM.  �� @�5(�U��#P, 1��, 3���45��NPX_�ASt�� 0��A�DD���$SI}Z��$VAR��.�TIP/�.��A�ҹM�ǐ��/�1�$+ U"S�U!Cz���OFRIF��J�S���5Ԓ�NF�Ѝ�n � xp`SI���TE�C���CSGL��TQ2�@&����<� ��STMT��,�P �&BWuP��S�HOW4���SV|�$�� �Q�A00�@Ma}����@ �����&���5��U6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G��0 G���0G���@G���PG��1	1	1�	1+	18	1E	2���2��2��2��2���2��2��2��2���2��2	2	2�	2+	28	2E	3���3��3��3��3���3��3��3��3���3��3	3	3�	3+	38	3E	4��4��4��4��4���4��4��4��4���4��4	4	4�	4+	48	4E	5��5��5��5��5���5��5��5��5���5��5	5	5�	5+	58	5E	6��6��6��6��6���6��6��6��6���6��6	6	6�	6+	68	6E	7��7��7��7��7���7��7��7��7���7��7	7	7*	7+	78	7E�һVP��UPDs�  �`NЦ�5��YSLOt�� � L��d���A�a�TA�0d��|�AL1U:ed�~�CUѰjg=F!aID_L�Ñe�HI�jI��$FI�LE_���d��$�2�fSA>�� h�O��`E_BLCK���b$��hD_CPUyM�yA��c�o�d��Y����R ��Đ
PW��!� oqLA��S=�ts�q~tRUN�qst�q�~t���qst�q~t ��T��ACCs���X -$�qLEN;��tH��ph�_��I��ǀLOW_A�XI�F1�q�d2�*�MZ���ă��W�Ipm�ւ�aR�TOR���pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v�������GTCV��؁��T�� ي�����t�V�����V�Jj�R�MA�i�JH��m�u�b����q�2j�#�U�{�t�K�JK��VK;���H����3��J0����JJv��JJ��AAL��Pڐ��ڐԖ4Օ5���N1���ʋƀW�%LP�_(�g�,��p�r�� `�`GR�OUw`��B��N�FLIC��f�RE�QUIRE3�EB�U��qB���w�2�����p���q5�p��{ \��APPR��iC}�Y�
ްEN٨�CLO7��S_M���H���u�
�qu�7� ���MC������9�_MG��C�C�o��`M�в�N�BRKL�NOL|�N�[�R��_LINђ�|�=�J����Pܔ������������������6ɵ�̲8k�+��q���� ��
��q�)��7�PATH 3�L�B�L��H�wࡠm�J�CN�CA��ؒ�ڢB�IN�rUChV�4a��C!�UM��!Y,���aE�p�����ʴ���PAYL�OA��J2L`R'_AN�q�Lpp����$�M�R_F2�LSHR��N�LO�ԡ�Rׯ�`ׯ�ACRL_G�ŒЛ� �r�Hj`߂$HM�^��FLEXܣ�q}J�u� :� ������������1�F1�V�j�@�@R�d�v�������E�� ��ȏڏ����"�4� q���6�M���~��U��g�y�ယT��o�X ��H������藕?� ����ǟِݕ�ԕ�����%�7��P��J�� � V�h�z����`AT�採@�EL��� S��J|��v��JEy�CTR���~�TN��FQ��H�AND_VB-����v`�� $��Fa2M����ebSW�q��'��� $$	MF�:�Rg�(x�,4�%��0&A�`�=���aM)F�AW�Z`i�A�w�A��X X�'pi�D*w�D��Pf�G�p�)CSTk��!x��!N��DY�pנM�9$`%� ��H��H�c�׎���0� ��Pѵڵ�쵠�������J��� ���1��R�6���QASYMvř����v��J���cі�_SH>��ǺĤ�ED� ���������J�İ�%��C�IDِ�_VI�!X�2PV_UCNIX�FThP�J�� _R�5_Rc�cTz�pT�V ��@���İ�߷��U I�������Hqpfˢ��aEN�&3�DI����O4d`J�� x g"IJAA�az�aabp�coc��`a�pdq�a� �^�OMME��� h�b�RqT(`PT�@ � S��a7�;�Ƞ�@ȷh�a�iT�@<� �$DUMMY9�Q�$PS_��R�FC�  S�v �� ���Pa� XXƠ���STE����SBRY�M21_�VF�8$SV_E�RF�O��LsdsCLRJtA��Odb`�O�p � D ?$GLOBj�_LO���u�q�cAp�rܛ@aSYS�qADqR``�`TCH  � ,��ɩb�oW_NA����7���SR���l ���
*?� &Q�0"?�;'?�I)?� Y)��X���h���x��� ���)��Ռ�Ӷ�;�� Ív�?��O�O�O�D��XSCRE栘pњ���ST��s�}y`����/_:HA�q� TơgpTYP�b���G�aG���Od0I�S_䓀d�UE�Md� ����ppS<�qaRSM_�q*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCOUx��S�Ԕ 1�!��UE&��Ubwr��PoROGM�FL@o$CUgpPO�Q���5�I_�`H� �� 8�� �_H�E�PS�#��`RY ?�qp�b��d�p�OUS�� �� @6p�v$/BUTTp�RpR�COLUMq�e���SERV5�PA�NEH�q� � ��@GEU���F�y��)$HELP�õ)BETERv�) ෆ���A � ���0��0��0ҰI)N簪c�@N��I�H�1��_� �֪�LN�r� Ʉqpձ_ò=�$9H��TEXl��Ο�FLA@��RELV��D`������5��M��?,�ű��m����"�US�RVIEW�q� �<6p�`U�`�N�FI@;�FOCUܕ�;�PRI@mx�`�QY�TRIP�q�m�UN<`Md�� #@p�*eWAR�N)e6�SRTOLJ%��g��ᴰONCwORN��RAU��r��T���w�VIN�~Le� $ג�PATH9�גCA;CH��LOG�!�LIMKR����v����HOST��!�b�R��OBOYT�d�IM>� �� ���Zq�Zq�;�VCPU_AVgAIL�!�EX	�!AN���q��1r��1r��1 �ѡ�p��  #`C�����@$TOOL�$���_JMP� y���e$SS��|�ϑVSHIF��Nc�P�`ג�E��ȐR����OSURz��Wk`RADIL����_�a��:�9a���`a�r��LULQ$�OUTPUT_BM����IM�AB ��@�rTILSCO��C7��� ����&��3�� A���q���m�I�!2G�n�y@Md�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM���F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? �ϑZABC%��  $�"R���
ϐ�$$CLA}S������!�pϐ� � VIRT8]��/ 0ABS�����1 5�� <  �!F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o �$6HZi{0-�A�XL�p��"�63  �{tIN��qztGPRE�����v�p��uLARMRECOV 9�rwt�NG�� .;	 =#�
�.�0�PPLIC��?�5�p�H�andlingT�ool o� 
�V7.50P/2{3 �!�PB���
��_SWt� �UP�!� x�F�0��t���Aϐv�� 864�� �it�y� N�2 7D�A5�� j� �QB@��o�Ngoneisͅ˰ ��T�]�!�LAAxyrPE_l�V�uT��s9�UTO�"�Њt�y��?HGAPON
0g��1��Uh�D 1581����̟�ޟry����Q 1���p�,�蘦����;�@��q_��"{�" �c��.�H���D�HTTHKYX��"� -�?�Q���ɯۯ5��� �#�A�G�Y�k�}��� ����ſ׿1����� =�C�U�g�yϋϝϯ� ����-���	��9�?� Q�c�u߇ߙ߽߫��� )�����5�;�M�_� q�������%��� ��1�7�I�[�m�� ��������!���� -3EWi{�� ����)/ ASew���� /��/%/+/=/O/ a/s/�/�/�/�/?�/ �/?!?'?9?K?]?o? �?�?�?�?O�?�?�?0O#O]���TO�E��W�DO_CLEA�N��7��CNM  � �__�/_A_S_�DSPDgRYR�O��HIc��M@�O�_�_�_�_o o+o=oOoaoso�o�o0���pB��v �u����aX�t������9�PLUGG���G��U�WPRCvPB�@��_�orOr_7�/SEGF}�K[mw xq�O�O�����?rqLAP�_�~q� [�m��������Ǐُ�����!�3�x�TO�TAL�f yx�USWENU�p�� �H����B��RG_STRING 1u��
�Mn�S�5�
ȑ_ITE;M1Җ  n5��  ��$�6�H�Z�l�~� ������Ưد����� �2�D�I/O SIGNAL̕�Tryout� ModeӕI�np��Simul�atedבOu�t��OVER�R�P = 100�֒In cyc�l��בProg� Abor��ב~��StatusՓ�	Heartbe�atїMH F�aul��Aler'�W�E�W�i�{ύ���ϱ�������  �CΛ�A����8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|���WOR{pΛ��(� ������ ��$�6�H� Z�l�~���������������� 2PO ̛�X ��A{�� �����/ ASew�����SDEV[�o �#/5/G/Y/k/}/�/ �/�/�/�/�/�/??�1?C?U?g?y?PALTݠ1��z?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O_�?GRI�`ΛDQ �?_l_~_�_�_�_�_ �_�_�_o o2oDoVo�hozo�o�o�o2_l�R ��a\_�o"4F Xj|����� ����0�B�T��oPREG�>�� f� ��Ə؏���� �2� D�V�h�z��������ԟ���Z��$AR�G_��D ?	����;���  	$�Z�	[O�]O���Z�p�.�SBN_C�ONFIG �;�������CI�I_SAVE  �Z�����.�TC�ELLSETUP� ;�%HO�ME_IOZ�Z�%MOV_��
��REP�lU�(�UT�OBACKܠ���FRA:\z� \�z�Ǡ'`�z���ǡi�WINI�0z����n�MESSAG༠�ǡC���ODEC_D������%�O��4�n�PAUSX!��;� ((O >��ϞˈϾϬ����� �����*�`�N߄��rߨ߶�g�l TSK�  wͥ�_�q�UgPDT+��d!�~A�WSM_CF���;���'�-�G�RP 2:�?� �N�BŰA��%�XS�CRD1�1
7� �ĥĢ������ ����*�������r� ����������7���[� &8J\n��|*�t�GROUN�|UϩUP_NA��:�	t��_E�D�17�
 ��%-BCKED�T-�2�'K�`����-t�z��q�q�z���2 t1�����q�kp�(/��ED3/ ��/�.a/�/;/M/ED4�/t/)?�/.p?p?�/�/ED5`? ?�?<?.�?O�?�?ED6O�?qO�?.pMO�O'O9OED7�O `O_�O.�O\_�O�O�ED8L_,�_�^�-�_ oo_�_ED!9�_�_]o�_	-9o�oo%oCR_  9]�oF�o�k� � ?NO_DEL���GE_UNUSE���LAL_OU�T ����W?D_ABORﰨ~���pITR_RT�N��|NONS�k���˥CAM�_PARAM 1�;�!�
 8
�SONY XC-�56 23456�7890 �~��@���?��( А\�
����{����^�HR5pq�̹��ŏR57ڏ��Aff��K�OWA SC31�0M
�x�̆�d @<�
��� e�^��П\�����*�<��`�r�g�CE�_RIA_I�j!�=�F��}�vz� ��_LIU�Y]�����<���FB�GP 1��Ǯ�M�_�q��0�C*  ����CU1��9��@��G��Z�CR�C]��d��l��s��R�����U[Դm��v����}����� C���ő(�����=�HE�`ONFIǰ�B��G_PRI 1�{V���ߖϨϺ�����������CHK�PAUS�� 1K� ,!uD�V�@� z�dߞ߈ߚ��߾��� ���.��R�<�b���O��������_MOR�� }���BZ?����� 	 �����*��N�`�����H��?��q?;�;����R��K��9�P���>ça�-:���	�

��M���p U�ð��<��,~���DB���튒)
�mc:cpmidcbg�f�:���%B��C¥�p�/��  �9 :
9 ;� �s>+��p"�p#U��?�͋��bUg�/���p�Uf�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����g=L���'MC��1����?43���1��t�īCz�  BHH�CPU�eB��CF��;.<C����C5rY
K�D��nyDQ��D���>��D�;D���=�F��>F�$�G}RB�7Gz�0��Y	��Y!�&w�1����s���.�p���b���BDw�M@x8�b�1Ҩ�, fAD�p@�0EYK�EX��EQ�EJP� F�E�F�� G��>^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE ���F 
Q��;��(P  B_<_��Rb����	op6C4P)�Y
s@ ]AQ�2Js@C�0B3�MaC{@�@*cw��UT�pFPROG %�z�o�oigI�q���v���ldKEY_TBL�  �&S�#� �	�
�� !�"#$%&'()�*+,-./01�i�:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇���������������������9��p`LCK�l4�<p`�`STAT ��S�_AUTO_DO��5�INDTG_EN#���R�Q�?�1�T2}�^�STsOPb���TRLr`�LETE��Ċ_�SCREEN ��Zkcsc���U��MMENU� 1 �Y  <�l�oR�Y1�[� ��v�m���̟����� ٟ�8��!�G���W� i��������ïկ�� 4���j�A�S���w� ����迿�ѿ���� T�+�=�cϜ�sυ��� �ϻ�������P�'� 9߆�]�o߼ߓߥ��� �����:��#�p�G� Y����������� $����3�l�C�U��� y����������� ���	VY)�_MAN�UAL��t�DBC�O[�RIGڇ
�DOBNUM� ��B1� e
�PXWOR/K 1!�[�_�U/4FX�_A�WAY�i�GC�P  b=�Pj_A!L� #�j�Y��܅t `�_�  1"�[ , 
�mgP�&/~&lMZ�IdP�x@P@#ONTImMه� d�`&�
�e�MOTN�END�o�REC�ORD 1(�[8g2�/{�O��!�/ ky"?4?F?X?�(`? �?�/�??�?�?�?�? �?)O�?MO�?qO�O�O �OBO�O:O�O^O_%_ 7_I_�Om_�O�_ _�_ �_�_�_Z_o~_3o�_ Woio{o�o�_�o o�o Do�o/�oS�o L�o����@� ��+�yV,�c�u� �������Ϗ>�P�� ���;�&���q���� ����P�ȟ�^���� ��I�[����� ����$�6�������jTOLERENCwsB���L�͖ �CS_CFG �)�/'dMC�:\U�L%04dO.CSV�� c���/#A ��CH��z� //.ɿ��(S��RC_OUT �*��1/V�SG�N +��"���#�10-FEB�-20 18:2�4027-JAN�p�21:48+? P;��ɞ��/.��f�pa�m��PJPѲ���VERSION� Y�V2�.0.�ƲEFLOGIC 1,�/ 	:ޠ=��ޠL��PROG_�ENB��"p�UL�Sk' ����_WRSTJNK ��"�fEMO_OPT?_SL ?	�#�
 	R575/#=�����0�B�|���TO  ��صϗ��V_F EX�d�%��PAT�H AY�A\p�����5+ICT�-Fu-�j�#�egS�,�STBF_TTS�(@�	d���l#!w�� �MAU��z�^"MS%WX�.�<�4,#�
Y�/�
!J�6�%ZI~m��$SBL_FAUL(�y0�9'TDIA[��1<�<� ����1234567G890
��P�� HZl~���� ���/ /2/D/V/hh/�� P� ѩ�yƽ/��6�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�,�/�UMP���� �ATR���1OC@�PMEl�OOY_T�EMP?�È�3pF���G�|DUNI���.�YN_BRK �2_�/�EMGDI_STA��]��E�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�Q�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��QDzr�=#�דQXT_BWD��p��xf́t�_DIn�� 9�5�d��T�QsRֆSTEP���:P�OP_D�Ov�f�PFAC�TORY_TUN�wdM�EATUROE :�5̀rQ�Handl�ingTool ��� \sfm�English �Dictiona�ry��roduAA Vis�� Master��ީ�
EN̐nalog I/O��ީ�g.fd̐ut�o Softwa�re Update  F OR��matic Ba�ckup��H59�6,�ground Editޒ�  1 H5�Camera�F���OPLGX�elyl𜩐II) X�7ommՐshw���7com��co����\tp���pan}e��  opl���tyle sel�ect��al C�nJ�Ցonit;or��RDE���tr��Relia�b𠧒6U�Dia�gnos(�푥�5�528�u��he�ck Safet�y UIF��En�hanced Rob Serv%��q ) "S�r�U?ser Fr[������a��xt. D�IO �fiG� �sŢ��endx�Ekrr�LF� pȐ�ĳr됮� ���� � !��FCTN /Menu`�v-�ݡ|���TP Inې�fac�  ER_ JGC�pב_k Exct�g���H558��igh�-Spex�Ski~1�  2
P���?���mmunic�'�ons��&�l�uqr�ې��ST Ǡ���conn��2ި�TXPL��nc=r�stru�����"FATKA�REL Cmd.� LE�uaG�54�5\��Run-T�i��Env��d�
!���ؠ++�s�)�S/W��[�LicenseZ��� 4T�0�ogB�ook(Syڐm�)��H54O�MA�CROs,\�/O�ffse��Loa��MH������r,� k�MechStop Prot����� lic/�MiвShif����ɒ�Mixx��)���x�SPS�Mode �Switch�� �R5W�Mo�:�.�� 74 ����g��K�2h�ult�i-T=�M���LN (Pos�Regiڑ������|d�ݐt Fun��⩐.�����Numx~����� lne�|�ᝰ Adjup������  - W���tatuw᧒T��RDMz�o}t��scove U�9���3Ѓ�uest 492�b*�o�����62;�?SNPX b ����8 J7`���Li3br��J�48����"�� �Ԅ�
�6O��� Parts i�n VCCMt�3�2���	�{Ѥ�J9�90��/I� 2� P��TMILI�B��H���P�A�ccD�L�
TE�$TX�ۨ�ap1�S�Te����pke�y��wգ�d���Unexcep=tx�motnZ���������є�� qO���� 90J��єSP CSXC`<�f��Ҟ� Py�sWe}���PRI��>vr�t�menz�� ��iPɰ�a�����vGri=d�play��v���0�)�H1�M-�10iA(B20�1 �2\� 0\}k/�Ascii��l�Т�ɐ/�Col���ԑGuar� �
�� /P-�ޠ"Kv��st{Pat �:�!S�Cyc��΂�orie��IFn8�ata- quҐ��� ƶ��mH57m4��RL��am����Pb�HMI D�e3�(b����PC�Ϻ�Passwo�+!��"PE? Sp�$�[���tp��� vKen��Tw�N�p��YELLOW B�OE	k$Arc��v�is��3*�n0W�eldW�cialh�7�V#t�Op�����1y� 2F�a�portN�(�p�T1�T� �� �ѳxy]�&TX��t�w�igj�1� b� �ct\�JPN �ARCPSU P�R��oݲOL� S;up�2fil� &�PAɰאcro�� �"PM(����O$SuS� eвtex�ԣ r���=�t�s'sagT��P���P@�Ȱ�锱�rt�W��H'>r�dpn��n1
t�!�� z ��ascbi?n4psyn��+A}j�M HEL��NCL VIS �PKGS PLOA`�MB �,�4�VW�RIPE �GET_VAR {FIE 3\t���FL[�OOL: �ADD R729.FD \j8'�iCsQ�QE��DVvQ��sQNO WTW�TE��}PD  ��^��biRFOR ���ECTn�`��ALSE ALAfP�CPMO-130�  M" #h�D�: HANG F�ROMmP�AQfr���R709 DR�AM AVAIL?CHECKSO!���sQVPCS SU��@LIMCHK �Q +P~dFF PO�S��F�Q R59�38-12 �CHARY�0�PR�OGRA W�SwAVEN`AME�P�.SV��7��$E�n*��p?FU�{�TR}C|� SHADV0�UPDAT KC|JўRSTATI�`~�P MUCH y��1��IMQ MO?TN-003��}��ROBOGUIDE DAUGH�a8���*�tou�����I� Šhd�ATH|�PepMOVET��ǔVMXPACK� MAY ASS�ERT�D��YCL�fqTA�rBE C�OR vr*Q3rA�N�pRC OPToIONSJ1vr̐PSH-171Z@-x�tcǠSU1�1`Hp^9R!�Q�`_T�P���'�j�d{tb�y app wac 5I�~d�PHI����p�aTEL�MX?SPD TB5bLu� 1��UB6@�qEN�J`CE2�61��p���s	�may n��0� R6{�R� >�Rtraff)��� 40*�p��fr���sysvar ?scr J7��cNj`DJU��bH �V��Q/�PSET �ERR`J` 68���PNDANT �SCREEN U�NREA��'�J`D��pPA���pR`IgO 1���PFI�p}B�pGROUN�P�D��G��R�P�QnRS�VIP !p�a�PD�IGIT VER�S�r}BLo�UEW~ϕ P06  �!��MAGp�abZV��DI�`� SS�UE�ܰ�EPL�AN JOT` D�EL�pݡ#Z�@D�͐CALLOb�Q �ph��R�QIPN�D��IMG�R7{19��MNT/�PWES �pVL�c���Hol�0Cq���tP�G:�`C�M�caynΠ��pg.v�S�: 3D mK�v_iew d�` �p���ea7У�b� o�f �Py���ANN�OT ACCESGS M��Ɓ*�t47s a��lok��Flex/:�Rw�!mo?�PA?�-�����`n�pa S�NBPJ AUTO-�06f����TB���PIABLE1q �636��PLN:Y RG$�pl;pNW7FMDB�VI���t�WIT 9x�0@o���Qui#0�ҺPN� RRS?pUSB��� t & remov�@ )�_��&�AxEPFT_=� �7<`�pP:�OS�-144 ��h qs�g��@OST� �� CRASH �DU 9��$�P�pW� .$��L/OGIN��8&�J���6b046 issue 6 Jg���: Slow ��st��c (HCos`�c���`IL`�IMPRWtSPO�T:Wh:0�T�S�TYW ./�VMGqR�h�T0CAT��hos��E�q���� �O�S:+pRSTU' k�-S� ����E:��pv@�2�N� t\hߐ��m ���all��0�  �$�H� WA͐��3 CNT0 T��� WroU�alacrm���0s�d � @�0SE1���r R{�OMEBp���K� �55��REàSEs�t��g    } �KANJI��no���INIS?ITALIZ-p�d�n1weρ<��dr�� lx`�SCI�I L�fail�s w�� ��`�YSTEa���o��PvЧ IIH���1W�G�ro>Pm ol\�wpSh@�P��Ϡn� cflxL@АW{RI �OF Lq���p?�F�up��d�e-rela�d� "APo SY�c}h�Abetwe:0IND t0$gb#DO���r� `��GigE�#ope�rabilf  P�AbHi�H`��c�le{ad�\etf�P8s�r�OS 030��&: fig��GL�A )P ��i��7�Np tpswx�B��If�g�������5aE�a EXC�E#dU�_�tPCLO�S��"rob�NTdpFaU�c�!����PNIO V750�Q1��Qa��'DB ��P M�+Pv�QED�DET���-� \rk��ON�LINEhSBUG�IQ ߔĠi`Z�IB�S apABC �JARKYFq� ����0MIL�`� R��pNД �p0GAR��D*pR��P�"'! jK�0cT�P��Hl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P��`WIBPK05��!FȐB/��BUSY RUNN��C "�򁐈��R-p��LO�N�DIV�Y�CUL��fsfoaBW�p����30	V��ˠIT�`�a505.�@O=F�UNEX�P1bҬaf�@�E��SVwEMG� NMLq�� D0pCC_SA�FEX 0c�08"qD. �PET�`N@�#'J87����RsP�TA'�M�K�`K��H GUNCHG^۔MECH�pMcz� T�  y, g@��$ ORY LE�AKA�;�ޢSP�Em�Ja��V�tGR�Iܱ�@�CTLN�TRk�FpepR��j50�EN-`IN�����p �`�Ǒ�k!��T3/dqo�SKTO�0A�#�L�pA �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`D	U��aO�supk�t4� � P�F� Bnf��Q�PSVGN-18��V�SRSR)J�UP�a2�Q�#D�q� l O��QBRKCTR5Ұ�|"-��r�<pc�j!INVP�D ZO� ��T`�h#�Q�cHset,x|D��"DUAL� �w�2*BRVO117 A]�TNѫt�+bTa2473��q.?���sAUz�i�B�complete���604.� -^�`hanc�U�� F��e8��  ��npJtPd!q��`��w� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP��R�R(}\xPe� aʰ�I���E��1��p�� j  �� xSP�^P �A�AxP�q �5 sig��a��"AC;a��
�bCe�xPb_p��.pc�]l<bHbcb_cicrc~h<n�`tl1� ~`xP`o�dxP�b]o2�� �cb�c�ixP�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`�cptlibxzxP�l�cr�xrxP\�blpsazEdxP_fm�} gcxP�x���o|sp�or�mc(��ob_jzo"p�u6�wf��t���wms�1q��sld�)��jmc�o\�n�b�nuhЕ��|st�e���>�pl�qp�iwc1k���uvf0uߒ<��lvisn�CgoaculwQ
E �F  ! Fc.f9d�Qv�� qw����Data Acq/uisi��nF�|1��RR631`��TR��QDMCM �2֝P75H�1�P58�3xP1��71��559`�5�P57<PxP�Q����(���Q���o pxP!daq�\�oA��@�� �ge/�etdms�"�DMER"؟,�p#gdD���.�m���-��qaq.<᡾xP#mo��h���f{�u��`13��MACRO�s, SksaffP�@z����03�SR�QT(��Q6��1�Q9ӡ��R�ZSh��PxPJ6+43�@7ؠ6�P�@�PRS�@���e �Q��UС PIK�Q5?2 PTLC�W���xP3 (��p/O ��!�Pn �xP5���03\sfmn�mc "MNMCPq�<��Q��\$AcX�FM���ci,Ҥ�X�����cdpq+�
�sk��SK�xP�SH5�60,P��,�y�r�efp "REF�p�d�A�jxP	�of��OFc�<gy�to��TO_����ٺ����+je�u��caxis2�xPE�\�}e�q"ISDTc�|�]�prax ���MN��u�b�is�de܃h�\�w�xP!� isbasic���B� P]��QA7xes�R6�������.�(Ba�Q�ess��xP���2�pD�@�z�atis�� ��(�{�����~��m��FMc�u�{�
���MNIS��ݝ�� ��x����ٺ��x�� j75��Dev�ic�� Inte�rfac�RȔQJ�754��� xP�Ne`��xP�ϐ2��б����dn� "�DNE���
tpodnui5UI��ݝ	bd�bP�q_rsofOb
?dv_aro��u�����stchkc��z	 �(}�onl��G!ff L+H�J(��"l"/��n�b��z�haSmp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!2���xpc_2pcch=m��CHMP_�|8бpevws��2�ΌpcsF��#C �SenxPacro0�U·�-�R6�Pd�@xPk�����p��gT�L��1d M�2`��8��1c4ԡ�3 qem��GEM,\i(��Dgesnd�5���H0{�}Ha�@sy���c��Isu�xD��Fmd ��I��7�4���u���AccuCal�P��4� ��ɢ7ޠB0���6+6f�6��9!9\aFF q�S(�U��2�
X�p�!Bd�ѳcb_�SaUL�� � �� ?�ܖto���otplus\tsrnغ�qb�W�p��t���1��To�ol (N. A�.)�[K�7�Z�(P��m����bfclls� k94�"K4p���qtpap� �"PS9H�stpswo��p�L7��t\�q����D�yt5� 4�q��w�q��� �Mz�uk��rkey�����s��}t�sfe7atu6�EA��� cf)t\Xq�����df�h5���LRC0�md�!�587���a�R�(����2V��8lc?u3l\�pa3}@H�&r-�Xu���t,�� �q "�q�Ot��~ ,���{�/��1c�}����y�p�r��5����S�XAg�-�y���Wj�874�- iR�Vis���Queu�� Ƒ�-�6�1$���(����u����tӑ����
�tpv�tsn "VTS�N�3C�+�� v\pR�DV����*�prd�q\�Q�&�vst�k=P������nmx&_�դ�clrqν���get�TX��Bd���aoQϿ�0q�str�D[� ��t0�p'Z����npv��@�enlIP0��D!0x�'�|���sc ߸��tvo/��2�q���vb����q����!���h]��(� Control�PRAX�P5��5�56�A@59�P5-6.@56@5A��J69$@982 �J552 IDVR7�hqA���16�Hx���La�� ���Xe�frlparwm.f�FRL��am��C9�@(F �����w6{���A���QJ643�� 5}0�0LSE
_p�VAR $SGS�YSC��RS_UNITS �P�2�4�tA�TX.$VN�UM_OLD 5`�1�xP{�50+��"�` Funct ���5tA� }��`#@�`E3�a0�cڂ��9����@H5נ� �P���(�A����۶}�����ֻ}��bPR�b�߶~ppr4�TP�SPI�3�}�r�10�#;A� t�
`���1���96�����%C�� Aف��J�bIncr�	����\�`��1o5qni4�MNINp	xP�`����!��Hour_  � 2�21 �A�AVM���0 ���TUP ��?J545 ���6162�VC�AM  (��CLIO ���R6�N2�MSC� "P ��STYL�C�28�~ 13\�NRE� "FHRM S�CH^�DCS}U%ORSR {b��04 �E�IOC�1 j 5742 � os| �? egist��Ի��7�1�oMASK�934"�7 ��OCO ���"3�8��2���� 0 HB��ڢ 4�"39N� R�e�� �LCHK�
%OPLG%��3�"%MHCR.%MCd  ; 4? ��6 d�PI�54�s� D[SW%MD� pQ�K!637�0�0p"�Y1�Р"4 �6<2?7 CTN K � +5 ���"7��<2�5�%/�T�%FRD�M� �Sg!��9�30 FB( NBA��P� ( HLB  7Men�SM$@jB�( PVC ��290v��2HTC�C?TMIL��\@?PAC 16U�hA�J`SAI \@ELN���<29s�UE�CK �b�@FRM� �b�OR���I�PL��Rk0CSXsC ���VVFna}Tg@HTTP �N!26 ��G�@~obIGUI"%�IPGS�r� H863 qb�!�07r�!�34 �r�84 �\so`! Qx`CC3� Fb�21�!969 rb!51 ���!S53R% 1!s3!���~�.p"9js V{ATFUJ775"���pLR6^RP�WS�MjUCTO�@xT5�8 F!80���1X�Y ta3!770 ���885�UOL�  GTSo
�{` L�CM �r| TSS��EfP6 W�\@CPgE `��0VR� �l�QNL"��@00�1 imrb�c3� =�b�0���0�`6� w�b-P- R-��b8n@5EW�b9 �Ґa� ���b�`ׁ~�b2 2000���`3��`4*5�`5 !�c�#$�`7.%�`�8 h605? U�0�@B6E"aRp76� !Pr8 t�a�@�tr2 iB/d�1vp3�vp5 ȂRtr9Σ�a4@-pN�r3 F��r5&0�re`u��r7 ��r�8�U�p9 \h7�38�a�R2D7�"�1f��2&�7<� �3 7iC���4>w5Ip�Or60� C�L�1bEN�4 I�pyL�uP��@N�&-PJ8�N�8NeN�C9 H�r`�E�b7]�|���8�ВࠂG9 2��a`0�q�Ђ5�%U097 �0��@1�0���1� (�q�3 5R ���0���mpU���0�0�7*�H@(q��\P"RB6�q124�b;��@���@�06� x�3 pB�/x�u ��x�6 H606�a1� ��7 6 ���p��b155 ����7>jUU162 ��3 g��4*�65 2e "_��P�4#U1`���B1���`=0'�174 �q���P�E186 R L��P�7 ��P�8&��3 (�90 B�/�s191����@2s02��6 3���A�RU2� d��O2 b2h`��4��b��2�4���19v RQ�2��u2d�Tpt)2� ��H�a2hP�$2�5���!U2�p�p"
�2�p��@5�0-�@��8 @�9��T�X@�� �e5�`rb	26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0@�gqGA���a�52ѐ�Ḳ6�6�0ہ5� ׁ2��84�E��9�EU5@ٰE\�q5hQ`S�2ޖ5�p\w�۲�pJ �4-P��5�p1\t�H�-4��PCH�7j��phiw�@��P�x��?559 ldu� P �D���Q�@�������A �`.��P>��8�g581�"�q58�!�AM۲T�A iC�a589��@�x���F�5 �a��12׀ 0.�1���,�2�����,�!P\h8��Lp ���,�7��6�084�0\��ANRS 0C}A��p��{��sran��FRA�� �Д�е���A%�� �ѹ�Ҍ�����(�� ��Ќ���З���������ь����$�G��1��ը��������� xS�`�q�  �����`6�4��M��iC/50T-H������*��)p46��� C��xN����m75s֐�� Sp��b46���v����ГM-7�1?�7�З����4A2������C��-��F��70�r�E��/h����O$��rlD���c7c7C� q��Ѕ���L��/���2\imm7c7�g������`���(��e�����"� �������a r��&c�T,�Ѿ�"��,��� ��x�Ex�m7�7t����k���5������)�iC��-HS-� B
_� >���+�Т�7U�]P���Mh7�s��a7������-9?�?/260L_������Q�������]�9pA/@���q�S�х��^�h621��c��92������.�)92c0�g$�@������)$��5$���pcylH"O"
�21�8��t?�350� ���p��$�
�� F�350!���0�x�9�U/0\m9��M9A3��4%�� s��3M$��X%u<���"him98J3����� i d�"m4~��103p�� ����h�794̂�&R���H �0����\���g�5A U��՜��0���*2� �00��#06�а�Ճ�է!07{r  ��������kЙ@�����EP�#�������?��#!�;&0s7\;!�B1P��@�A��/ЁCBׂ2�!��:/��?�ҽCD25�L����0�"l�2BL
#��B��\20�2_�r�re� ��X��1��N����A@��z��`C�pU��`��04��Dy	A�\�`fQ��s�U���\�5  ��� p�^P��<$85���+P=�ab1l��1LT��lA8�!uDnE(�.20T��J�1 e�bH85���b�Ռ�5[�16Bs��������d2��x��m6t!`Q����b�ˀ���b#�(�6iB ;S�p�!��3� ���b�s��-`�_�W80�_����6I	$�X5�1�U85��R�p6S����/�/+q�!@�q��`�6o��5m[o)�m6sW��Q�|�?��set06p h��3%H�5��10p$@����g/�JrH��?  ��A��856����F�� ���p/2��h�܅�✐)�5��̑v�𘜐(��m6��Y�H�ѝ̑m�6�Ҝ��ae6�DM����-S�+��H2�����Ҽ� � �r̑��✐��l���p1���F����2�\t6h T6H����Ҝ�'Vl ���ᜐ�V7ᜐ/�(���;3A7��p ~S��������4�`堜��V���!3��2��PM[��%ܖO�chn��vel5���8�Vq���_arp#���̑�.���2l_h�emq$�.�'�6415���5���?����F�����5g�L�ј�[���1��𙋹1<����M7NU�Р���eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h������ u���㜐��ZS0�!ܑ4���M-����S�$̑�ք �� 0���<�����07shJ�H�v�À�sF� �S*󜐳���̑���vl�3�A�T�#��Q�0��Te��q�pr����T@75j�5�dd�̑ 1�(UL�&�(�,���0��\�?���̑�a�� xSP���a�eD�w�2��(�	�2�C��A/���\�+p�<����21 (ܱ�CL S����B̺@��7F���?�<�lơ1L����c� ���u19�0����e/q���O���9�K��r9 (��,�Rs�ז�5�<G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O���M1!41w���2T@� _std��G�y�� �ң�H� jdgm����w0\� �1L� ��	�P�~�W*�b���t 5������3�,���E{���d���L��5\L��3�L�|#~���~!���4�#��O����h�L6A�������a2璥���44������[6\j4s ��·���#��ol�E"w�8Pk�����?0x j�H1�1Rr�>��]�2a�2Aw�P ��	2��|41�8��ˡ��@{� �%�A<��� +� ?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R�� ˑb�W���Fs���) �ѐ�!���a�1�����5��16�16C���C����0\imBQ��d����b��\Be5�-���DiL����O�_�<ѠPEtL �E�RH�ZǠPgω�am1l��u���̑�b@�<����<�$�T� ̑�F����Ȋ�DpbĜ�X"��hr��pĻ ���^P��9��0\� j971\�kckrcfJ�F�s�����c��e "CTME�r���ɛ�|�a�`main.[�8�g�`run}�_vc�#0�w�1Oܕ�_u����bctme���Ӧ�`ܑ�j73�5�- KARE�L Use {�U���J��1���p� Ȗ�9�B@���L�9��7j[�atk208 "K��(Kя��\��9��a���̹����cKRC4�a�o ��kc�qJ� &s�����Grſ�fs�D��:y��s�ˑ1X\�j|хrdtB�, L��`.v�q�� �spǑIf�Wfj52��TKQuto Seut��J� H5K7536(�932���-91�58(�9�BA��1(�74O,A$�(TCP Ak���/�)Y� �\tpqtool.v���v���! con�re;a#�Cont�rol Re�b{le��CNRE(� T�<�4�2���D�)���NS�552��q(g�� (򭂯4X�cOux~�\sfuts�UTS`�i�栜���At�棂��? 6�T�!�SA OO+D6���������,!��6c+� igt�t6i��I0�T�W8 ���la��vo58�o�bFå򬡯i��Xh��!Xk�0Y!8�\m6e�!6EC���v��6���������<16�A���A�6s����U�g�T|�,����r1�qR����Z4�T�����,#�eZp)g����<ONO0���uJ��tCR;��F<�a� xSP�f���prdsuchk� �1��2&&?���t��*D%$�r(�✑ �娟:r��'�s�qO��<scrc�C�\At�trldJ"o��\�V����Pay�lo�nfirm�l�!�87��7��A�3ad�! �?@ވI�?plQ��3���3"�q��x pl��`���d7��l�calC�uDu���;���mov�����initX�:s8O��a8�r4 ��r67A4|��e Genera#tiڲ���7g2q$g R� (S�h��c ,|�bE��$Ԓ\�:�"���4��4�4�. sg��5�F$d6"�e;Qp "SHA�P�TQ ngcr pGC�a(�&"� ���"GDA¶��r�6�"aW�/�$d�ataX:s�"tp�ad��[q�%tput;a__O7;a�o8�1�yl+s�r�?�:�#$�?�5x�?�:c O�:Ay O�:�IO�s`O%g�qǒ�?�@0\ۜ�"o�j92;!�Pp�l.Collis�QSkip#��@5� �@J��D��@\ވ�C(@X�7��7�|s}2��ptcls�#LS�DU�k?�\_� ets�`�< �\�Q��@���`dcKLqQ�FC;��J,όn��` (��4eN����T�{���' j(�c�����/IӸaȁ<��̠H������зa�e\mcc�lmt "CLM��/��� mate\v��lmpALM�?>p7qmc?�����2vm�q��%�3s��_�sv90�_x_msu�2L^v_� K�o��{in�8(3r<�c_logr��r�trcW� �v_3�~yc��d�<�ste��der$c;Ce� Fiρ��R��Q�?�l�enter߄|��(�Sd��1�TX�+fZK�r�a99sQ9+��5�r\tq\� _"FNDR����STDn$�LANG�Pgui��D⠓�S������csp�!ğ֙uf䟀ҝ�s����$�����e +�=����������������w�H�r\fn�_�ϣ��$`x�tcp�ma��- TCP������R638 aR�Ҡ��38��M7p,���Ӡ�$Ӡ��8p0Р�VS,�>�tk��99�a��B3���P�զԠ��D�2�����UI��t���hqB���8���������p���re8�ȿ��exe@4π��B���e38�ԡG�r�mpWXφ�var @�φ�3N�����v�x�!ҡ��q�R�BT $cOP�TN ask E�0��1�R MAS�0�H593/�96g H50�i�480ԅ5�H0��m�Q�K(��7�0�g�Pl�h�0ԧ�2�ORDP���@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`am��b��7�.f���u�d��r��splayD�E���1wПUPDT Ub��8o87 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60�q��B����qs�can��B���aAd@�������q`� �䗣�#��К�`2�� vlv��Ù�$�0>�b���! S���Easy/К�Ut�il��룙�511# J�����R7 ���Nor֠��inc�),<6Q�� �`c��"4�[���986(FVRx So����q�nd6����P��4� a\ (��
  ������"�d��K�bdZ����men7���- Me`tyFњ�Fb��0�TUa�577?i3R��\�5�au?��!� n����f������l\m�h�Ц�űE|h#mn�	��<\O�$��e�1�� l!���y��Ù�\|p�����B���Ћmh �@��:.aG!�� �/�t�55�6�!X��l�.us��Y/k)eOnsubL���eK�h�� �B\1;5g?�y?�?�?D��?*rmx�p�?Ktbox O�2K|?�G��C?A%das���?1ӛ#� � TR��/��P�4B�`�U@�P�V�P"�Q�P0�U �PO��P�"�T3�U�P �f�Pk"�2}�4�T�P �f�P2�"�Q5�S�Q@���R?Ă�Q3t.�PF׀al��P+O�n�P517��IN0a���Q(}g��PES	Tf3ua�PB�l�i�g�h�6�aq��P �� xS��` � n�0mbump�P�Q969g�69�Qq��P0�baAp�@>Q� BOX��,�>vche�s�>ve�tu㒣=wffse�3���]�;u`aW��:zol�sm<u�b�a-��]D�K�ib�Q�c����Q<twaǂ �tp�Q҄Taror Recov�br�O�P�642�����a�q��a⁠QErǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>��pjot��PXc��C��1�adb -�ail���nag���b�QR629�a�Q��b�P�  �
 � �P��$$CL~[q ����������$�PS?_DIGIT���"�!�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��������*璬1:P�RODUCT�Q0�\PGSTK�bV�,n�99�\����$FEAT_INDEX���~�� �搠ILECOM�P ;��)���"��SETUPo2 <��?�  N !��_AP2BCK �1=�  �)}6/E+%,/i/��W/�/~+/�/O/ �/s/�/?�/>?�/b? t??�?'?�?�?]?�? �?O(O�?LO�?pO�? }O�O5O�OYO�O _�O $_�OH_Z_�O~__�_ �_C_�_g_�_�_	o2o �_Vo�_zo�oo�o?o �o�ouo
�o.@�o d�o���M� q���<��`�r� ���%���̏[���� ���!�J�ُn����� ��3�ȟW������"� ��F�X��|����/� ��֯e������0��� T��x������=�ҿ �s�ϗ�,ϻ�9�b�t� P/ 2) *.VRiϳ�!�*���������Ɲ�PC�7�!�F'R6:"�c��χ��T��߽�Lը����x���*.F���>� �	N�,�k�x�ߏ��STM �⠸���Qа���!��iPendant? Panel���H��F���4������GIF�������pu����JPG&�P��<����	�PANEL1.D	T��������2�Y�G��
3w�����//�
4�a/��O///�/�
TP�EINS.XML�/���\�/�/�!�Custom T?oolbar?��PASSWOR�D/�FRS:�\R?? %Pa�ssword Config�?��? k?�?OH�6O�?ZOlO �?�OO�O�OUO�OyO _�O�OD_�Oh_�Oa_ �_-_�_Q_�_�_�_o �_@oRo�_voo�o)o ;o�o_o�o�o�o*�o N�or��7� �m��&���\� ����y���E�ڏi� �����4�ÏX�j��� �����A�S��w�� ���B�џf������� +���O��������� >�ͯ߯t����'��� ο]�򿁿�(Ϸ�L� ۿpς�Ϧ�5���Y� k� ߏ�$߳��Z��� ~�ߢߴ�C���g��� ��2���V����ߌ� ��?����u�
��� .�@���d������)� ��M���q�����< ��5r�%�� [�&�J� n��3�W� ��"/�F/X/�|/ /�/�/A/�/e/�/�/ �/0?�/T?�/M?�?? �?=?�?�?s?O�?,O >O�?bO�?�OO'O�O KO�OoO�O_�O:_�O ^_p_�O�_#_�_�_Y_��_}_o�_�_Ho)f��$FILE_DG�BCK 1=���5`��� ( �)
S�UMMARY.DyGRo�\MD:�o��o
`Diag� Summary��o�Z
CONSLOG�o�o�a
J�a�ConsoleO logK�[�`�MEMCHECK�@'�o�^qMe�mory Dat�a��W�)>�qHADOW����P��sShad�ow Chang�esS�-c-��)	FTP=��9�����w`qmmen�t TBD׏�W0�<�)ETHERNET̏�^�q��Z��aEther�net bpfiguration[���P��DCSVRF�ˏ��Ïܟ�q%��� verify� allߟ-c1P{Y���DIFFԟp��̟a��p%��diffc���q���1X�?�Q�� �����X��CH�GD��¯ԯi��px��� ���2`�G�Y��� ��� �GAD��ʿܿq��p���Ϥ�FY3h�O�aώ�� ��(�GAD������y��p�����0�UPDAT�ES.�Ц��[FORS:\�����a�Updates �List���kPS�RBWLD.CM�.��\��B��_pP�S_ROBOWEL���_����o��,o !�3���W���{�
�t� ��@���d�����/ ��Se����� N�r� =� a�r�&�J� ��/�9/K/�o/ ��/"/�/�/X/�/|/ �/#?�/G?�/k?}?? �?0?�?�?f?�?�?O �?OUO�?yOO�O�O >O�ObO�O	_�O-_�O Q_c_�O�__�_:_�_ �_p_o�_o;o�__o �_�o�o$o�oHo�o�o ~o�o7�o0m�o � ��V�z� !��E��i�{�
��� .�ÏR���������� .�S��w������<� џ`������+���O� ޟH������8���߯�n����$FIL�E_��PR����������� �MDONL�Y 1=4�� 
 ���w�į�� 诨�ѿ�������+� ��O�޿sυ�ϩ�8� ����n�ߒ�'߶�4� ]��ρ�ߥ߷�F��� j�����5���Y�k� �ߏ���B�����x� ���1�C���g���� ��,���P����������?��Lu�VI�SBCKR�<�a��*.VD|�4 OFR:\��4 �Vision VD file�  :LbpZ�# ��Y�}/$/� H/�l/�/�/1/�/ �/�/�/�/ ?�/1?V? �/z?	?�?�???�?c? �?�?�?.O�?ROdOO �OO�O;O�O�OqO_ �O*_<_�O`_�O�__�%_�_�MR_GR�P 1>4�L~�UC4  B�P�	 ]�ol`��*u����RHB ��2 ���� ��� ���He�Y�Q`ork bIh�oJd�o�Sc�o��oLp��M��e�K3MF�{5U�aS����o��o D���D��D�U��-��p9%���>C�}@��"A�_�lq?4?�ZA�[Dxq}�E�� F@ �r�d�a}J��N�Jk�H9��Hu��F!��/IP�s}?�`��.9�<9���896C'�6<,6\b��}B��B���C{��B���>B�B��� �"7�A����B��A���VA�SA��#���, A�PA�����|�ݏx����%���p�A6Β@U��{ �v�a�������П�� ��ߟ��<�'�hz;BH�P �a`�Q��QAK�@������ǯ�P
6�PJ��PJ�N˯�o�o�B��P5���@�3�3@���4�m�T�U�UU��U�~w�>u?.�?!x�^���ֿ���3��=[�z�=�̽=�V6<�=�=��=$q��~���@8�i7G���8�D�8?@9!�7ϥ��@Ϣ���:t�@ D��� Cϫo��C��P��P'�6��_ V� m�o��To��xo�� �o������A�,�e� P�b��������� ����=�(�a�L��� p��������������� ��*��N9r]� ������� 8#\nY�}� ������/ԭ// A/�e/P/�/p/�/�/ �/�/�/?�/+??;? a?L?�?p?�?�?�?�? �?�?�?'OOKO6OoO �OHߢOl��ߐߢ��O �� _��G_bOk_V_�_ z_�_�_�_�_�_o�_ 1ooUo@oyodovo�o �o�o�o�o�o Nu���� �����;�&�_� J���n�������ݏȏ ��%�7�I�[�"/� 描�����ٟ����� ��3��W�B�{�f��� ����կ������� A�,�e�P�b������� �O�O�O��O�OL� _p�:_�����Ϧ��� �����'��7�]�H� ��lߥߐ��ߴ����� ��#��G�2�k�2�� Vw����������� 1��U�@�R���v��� ����������- Q�u���r�� 6��)M4 q\n����� �/�#/I/4/m/X/ �/|/�/�/�/�/�/? ֿ�B?�f?0�BϜ? f��?���/�?�?�?/O OSO>OwObO�O�O�O �O�O�O�O__=_(_ a_L_^_�_�_�_���_ ��o�_o9o$o]oHo �olo�o�o�o�o�o�o �o#G2kV{ �h������ �C�.�g�y�`����� �����Џ���?� *�c�N���r������� �̟��)��M�_� &?H?���?���?�?�? ����?@�I�4�m�X� j�����ǿ���ֿ� ���E�0�i�Tύ�x� �Ϝ���������_,� �_S���w�b߇߭ߘ� �߼�������=�(� :�s�^������� ���'�9� �]�o� ���~����������� ��5 YDV� z������ 1U@yd�� v�����/Я*/�� 
/�u/��/�/�/�/ �/�/�/??;?&?_? J?�?n?�?�?�?�?�? O�?%OOIO4O"�|O BO�O>O�O�O�O�O�O !__E_0_i_T_�_x_ �_�_�_�_�_o�_/o ��?oeowo�oP��oo �o�o�o�o+=$ aL�p���� ���'��K�6�o� Z������ɏ��폴 � ��D�/ /z�D/ ��h/ş���ԟ��� 1��U�@�R���v��� ��ӯ������-�� Q�<�u�`���`O�O�O ���޿��;�&�_� J�oϕπϹϤ����� ���%��"�[�F�� Fo�ߵ����ߠo��d� !���W�>�{�b�� ������������� A�,�>�w�b������� ��������=���$FNO ����\��
F0l �q  FLAG>�(�RRM_CHK�TYP  ] �\�d �] ��{OM� _MIN� �	���� �  �XT SSB_C�FG ?\ �����OTP_D�EF_OW  �	��,IRCO�M� >�$GENOVRD_DO�s�<�lTHR�� d�dq_EN�B] qRAV�C_GRP 1@�I X(/  %/7//[/B//�/x/ �/�/�/�/�/?�/3? ?C?i?P?�?t?�?�? �?�?�?OOOAO(O�eOLO^O�OoROUr�F\� ��,�B,�8��?���O�O�O	__  D�UPE_�Hy_6�\@@m_B�=�vRp/��I�O�SMT�G���
�oo�+l�$HOSTC��1H�I� �\�zMSM�l[�bo�	12�7.0�`1�o  e�o�o�o#z �oFXj|�l60s�	anonymous��������ao�&�&� �o�x��o������ҏ �3��,�>�a�O� ���������Ο�U%� 7�I��]����f�x� �������ү���� +�i�{�P�b�t����� �������S�(� :�L�^ϭ�oϔϦϸ� �����=��$�6�H� Zߩ���Ϳs������ ����� �2���V�h� z��߰��������� 
��k�}ߏߡߣ�� �߬���������C� *<Nq�_��� ���-�?�Q�c�e J��n���� ���/"/E�X/ j/|/�/�/�% '/?[0?B?T?f?x? ��?�?�?�?�??E/�W/,O>OPObO�KDaE�NT 1I�K sP!�?�O  �P�O�O�O�O�O#_�O G_
_S_._|_�_d_�_ �_�_�_o�_1o�_o go*o�oNo�oro�o�o �o	�o-�oQu 8n������ ��#��L�q�4��� X���|�ݏ���ď֏�7���[���B�QUICC0��h�z�۟��1ܟ��ʟ+����2,���{�!ROUTER|�X�j��˯!PCJOG�̯��!192�.168.0.1�0��}GNAME �!�J!ROB�OT�vNS_CF�G 1H�I ��Auto�-started^�$FTP�/�� �/�?޿#?��&�8� JϏ?nπϒϤ�ǿ�π[������"�4�G�#�������������� ���������&�8�J� \�n��������� ����/�/�/F���j� �ߎ������������� 0S�T��x� ����!�3��G ,{�Pbt��C ����/�:/ L/^/p/�/��� 	/�/=?$?6?H?Z? )/~?�?�?�?�/�?k? �?O O2ODO�/�/�/ �/�?�O�/�O�O�O
_ _�?@_R_d_v_�_�O -_�_�_�_�_oUOgO yO�O�_ro�O�o�o�o �o�o�_&8J mo�o�����o )o;oMoO!��oX�j� |�����oď֏��� �/���B�T�f�x����^�ST_ERR �J;�����PDU�SIZ  ��^�P����>ٕWR�D ?z��� � guest���+�=�O�a��s�*�SCDMNG�RP 2Kz�Ð��۠\���K�� 	P0�1.14 8�q _  y���B    �;����{ �����������������������~ �ǟI�4��m�X�|��  �i  �  k
���� �����+�������_
���l�.x�+���"�l�ڲ۰s�d�������__GROU��L��� ��	��۠0�7K�QUPD  ����PČ�TY�g�����TTP�_AUTH 1M��� <!iP�endan����<�_�!KAR�EL:*������KC%�5�G��V�ISION SE!TZ���|��Ҽ� ����������
�W��.�@��d�v���CTRL N��������
�FFF�9E3���FR�S:DEFAUL�T�FANU�C Web Se/rver�
��� ���q��������������WR_CONF�IG O�� ����IDL_C_PU_PC"��sB��= �BH#�MIN.�BGNR_IO��� ����% NPT_SIM�_DOs}TPMODNTOLs} �_PRTY��=!OLNK 1P���'9�K]o�MAST�Er �����O_C3FG��UO���>�CYCLE����_ASG 1Q���
 q2/D/ V/h/z/�/�/�/�/�/��/�/
??y"NU�M���Q�IP�CH��£RTRY_CN"�u����SCRN����b�� ���R�����?��$J23_DSP_EN������0OBPR�OC�3��JOG�V�1S_�@��8��?�';ZO'??>0CPOSREO�?KANJI_�Ϡ�u�A#��3T ��x�E�O�ECL_LM �B2e?�@EYLOGWGIN��������LANGUAGgE _�=�Y }Q��LG�2U��V��� �x����j�PC � �'0������MC:�\RSCH\00�\˝LN_DISP V��������TOC�4Dz�\=#�Q�?PBOOK W+��o�0��o�o���Xi�o@�o�o�o�o~}	x(y��	ne�i�e�kElG_BUFF� 1X���}2 ����Ӣ���� ��'�T�K�]����� ������ɏۏ����#�P��ËqDCS �Zxm =��� %|d1h`���ʟܟg�IO 1[+# �?'����'�7� I�[�o��������ǯ ٯ����!�3�G�W� i�{�������ÿ׿��El TM  ��d ��#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߈tN�SEV�0m�TYP�� ��$�}�ARS"�(_�s>�2FL 1\��0��������������5�TP<P����DmNGNAMp�4�U�f�UPS`�GI�5�A�5s�_�LOAD@G �%j%@_MO�V�u����MAXUALRMB7�P8��y���3�0]&q��Ca]s�3�~�� t8@=@^+ طv�	��V0+�P�A5d�r���U������ E(iTy�� �����/ /A/ ,/Q/w/b/�/~/�/�/ �/�/�/??)?O?:? s?V?�?�?�?�?�?�? �?O'OOKO.OoOZO lO�O�O�O�O�O�O�O #__G_2_D_}_`_�_ �_�_�_�_�_�_o
o oUo8oyodo�o�o�o��o�o�o�o�o-��D�_LDXDISA�^�� �MEMO_{APX�E ?��
 �0y�����������I�SC 1_�� �O����W�i� ����Ə�����}�� ߏD�/�h�z�a���� ����������@� ��O�a�5��������� ���u��ׯ<�'�`� r�Y������y�޿� ۿ���8Ϲ�G�Y�-� ��}϶ϝ�����m������4��X�j�#�_M?STR `��}տSCD 1as}� R���N��������8� #�5�n�Y��}��� ���������4��X� C�|�g����������� ����	B-Rx c������ �>)bM�q �����/�(/ /L/7/p/[/m/�/�/ �/�/�/�/?�/"?H? 3?l?W?�?{?�?�?�?�n�MKCFG �b���?��LTA�RM_�2cRuB �3WpTN>BpMETPUOp�2�����NDSP_CMNTnE@F��E�� d���N��2A�O�D�EPOS�CF�G�NPST�OL 1e-�4@�<#�
;Q�1;U K_YW7_Y_[_m_�_�_ �_�_�_�_o�_oQo 3oEo�oio{o�o�a�A�SING_CHK�  �MAqODA�Q2CfO�7J�eD�EV 	Rz	�MC:'|HSIZ�En@����eTAS�K %<z%$1�23456789� ��u�gTRIGw 1g�� l<u%���3���>s�vvYPaq��kEM_INF 1h9G� `)�AT&FV0E�0(���)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ���ڄH������G�ֈAO�w�2�������џ ������ ��͏ߏP��t����� ��]�ί�����(� ۟�^��#�5����� k�ܿ� ϻ�ů6�� Z�A�~ϐ�C���g�y� �������2�i�C�h� ό�G߰��ߩ��ߙ� ���������d�v�)� ���߾�y������ ��<�N��r�%�7�I� [������9�&��J[�g��>O�NITOR�@G �?;{   	�EXEC1�3�2*�3�4�5��p��7�8�9�3 �n�R�R�R RRR(R4�R@RLR2Y2�e2q2}2�2��2�2�2�2*�3Y3e3��a�R_GRP_SV� 1it��q(�5��
��5���6�MO~q_DCd~��1PL_NAME� !<u� �!�Default� Persona�lity (from FD) �4�RR2k! 1j)TEX)TH��!�AX d�?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O�O�Ox2-?�O�O�O __0_B_T_f_x_�b<�O�_�_�_�_�_�_�o o2oDoVoho&xR�j" 1o�)&0\��b, �9��b~�a @D�  �a?��c�a?�`�a�a�A'�6�ew;��	l�b	 �xJp��`�`	p ��< �(p� ��.r� K�K� ��K=*�J����J���J�V��kq`q�P�x�|� @j��@T;f�r�f��q�acrs�I�� ��p���p�r�p�h}�3��´  ��>��ph��`z���Ζ"�Jm�q�  H�N��ac��$�dw���  �  �P� Q� �� | � а�m�Əi}	�'� � ��I� �  {����:�È�?È=���(��#��a	���I  �n @H�i~�ab�Ӌ�b�$w���"yN0��  'Ж��q�p@2��@�c���r�q5�C�p}C0C�@ C�����`
�A�1q   U@B�V~X�
nw�B0h�A��p�ӊ0�p�`���aDz����֏���Я	�pv��( �� -��I��-�=��A�a��we_q�`�p �?�ff ���m��� ��@��Ƽ�!@ݿ�>1�'  P�apv(�`ŀ�� �=�qst��?����`x`�� <�
6b<߈;�܍�<�ê<� <�&P�ό�AO��c1��ƍ��?fff?O�?&���qt@�.�?J<?�`��wi 4����dly�e߾g;� ��t��p�[ߔ�߸� ������ ����6�wh�F0%�r�!���߷�1ى����E��� E�O�G+� F�!���/���?��e�P���t���lyBL�cB��Enw4����� ��+��R��s����������h��Ô�>� �I�mXj���#A�y�weC��8������#/*/hc/N/wi�����v/3C�`� CHs/`
D=$�p�<!�!��ܼ��'�3A�A�A�R1AO�^??�$�?����±
=ç>�����3�W
=�#�]�;e����a@����{����<�>�(�B�u�����=B0�������	R��zH��F�G���G���H�U`E���C�+��}�I#�I���HD�F���E��RC�j=��>
I��@�H�!H�( E<YD0w/ O*OONO9OrO]O�O �O�O�O�O�O�O_�O 8_#_\_G_�_�_}_�_ �_�_�_�_�_"ooo XoCo|ogo�o�o�o�o �o�o�o	B-f Q�u����� ��,��P�b�M��� q�����Ώ���ݏ� (��L�7�p�[���� ��ʟ���ٟ���6�@!�Z�E�W���#1( �g��9�K���ĥ �����Ư!�3�8���!4�Mgs��,�IB�+8�J��a���{�d�d�����ȿP���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ�����X�����  %�� � �h�Vߌ�z߰�&�g�@/9�$�������7�����A�S�e�w�  ��������������2 F�$N�&Gb������X���!C���@���8�����F� �DzN�� F�P D�������)#B�'9K]o~#?���@@v
�4$8�8��:8�.
 v� ��!3EWi�{����:� ���ۨ�1���$MSKCFMA�P  ��� ���(.��ONREL  ��!9��E�XCFENBE'
8#7%^!FNCe/W$�JOGOVLIM�E'dO S"d�KE�YE'�%�RU�N�,�%�SFSPDTY0g&P%�9#SIGNE/W$TO1MOT�/T!��_CE_GRP [1p��#\x� �?p��?�?�?�?�? O�?OBO�?fOO[O �OSO�O�O�O�O�O_ ,_�OP__I_�_=_�_ �_�_�_�_oo�_:o��TCOM_C_FG 1q	-��vo�o�o
Va_AR�C_b"�p)UA�P_CPL�ot$N�OCHECK ?=	+ �x� %7I[m� �������!��.+NO_WAITc_L 7%S2NT^a�r	+�s�_E�RR_12s	)9��� ,ȍޏ��x����&��dT_MO���t��, �A�*oq�9�PARAM:��u	+��a��ß'g{�� =?�3�45678901 ��,��K�]�9�i��������ɯۯ��&g������C��cUM_RSPACE/��|����$ODR�DSP�c#6p(OF�FSET_CAR9T�o��DISƿ���PEN_FILE�尨!�ai��`OPT?ION_IO�/���PWORK ve7s# ��V������p�4�p�	 ����p��<���R�G_DSBL  ���P#��ϸ�R�IENTTOD �?�C�� !=#���UT_SIM_ED$�"���V��?LCT w}�h��iĜa[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ���� ��2�H(���H3k7HS�M5G�22G�?��Gp
͜��'f�/-,2�CR�>�D!�M#{Z/���3�����4y H "�c/u/�/�0B_����=jc��t�!�/ �/�"t32���~�/6  ��UP%�Q%��%�|T���S62�q?'e	'�� � �2I�� �  ��+==��ͳ?�;	��h	�0�I  �n @�2�.���Ov;��ٟ?&gN	 [OaA''�uD@!� Cb@C�@F#H!�/�O�O sb
�ATb@�@�@��@$�e`0Bb@QA�0Y�v: �13Uwz $oV_�/z_e_�_�_	���( �� -�2�1�1ta�UDa�c���:A-���~.  �?�ff���[o"o�_U�`oXâ�Q8���o�j>�1  Po�V(���eF0��f�Y���L�?˙���xb�P<
�6b<߈;����<�ê<�? <�&�,�/aA�;r�@Ov0P?offf?�0?&ipޘT@�.{r�J<?�`�u#	�B dqt�Yc�a�Mw �Bo��7�"�[�F� �j�������ُ� ���3����,���~(�E�� E��3?G+� F��a�� ҟ�����,��P�(;���B�pAZ�>� �B��6�<OίD���P� �t�=���a�s������6j�h��7o��>�S��O�����Fϑ�A�a�_���C3Ϙ�/�%?��?Ƀ��������#	���P �N||CH����Ŀ������@�I�_�'�3A��A�AR1A�O�^?�$�?���� �±
=�ç>����3�W
=�#� U���e���B��@���{����<����(�B��u��=B0�������	��b�H�F�G����G��H��U`E���C��+��I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻�������� � �9�$�]�H�Z��� ~�������������# 5 YD}h�� �����
C .gR����� ��	/�-//*/c/ N/�/r/�/�/�/�/�/ ?�/)??M?8?q?\? �?�?�?�?�?�?�?O �?7O"O[OmOXO�O|O �O�O�O�O�O�O�O3_:Q(������b���gUU��xW_i_2�3�8��_<�_2�4Mgs�_�_��RIB+�_�_�a?���{�mi�Go5okoYo�o}l��P'rP�nܡݯ�o=_`�o�_�[R?�Q�u���  �p���o��/�� S��z
uүܠ�������ڱ�����������  /�M�w��e��������l2 wF�$��Gb���t��a�`�p�S�C��y�@p�5�G�Y�۠F�� Dz��� F�P D��]����پ��ʯܯ�� ��~�?��ͫ@@�?�K��K���K���
 �|�������Ŀֿ �����0�B�T�f�ܽ�V� ���{���1��$PARA�M_MENU ?�3�� � DEF�PULSEr�	�WAITTMOU�T��RCV�� �SHELL_�WRK.$CUR�_STYL���	�OPT��PT�B4�.�C�R_DECSN���e��� �ߣ����������� !�3�\�W�i�{����USE_PROG %��%�����CCR���e�����_HOST !F��!��:���T�`�V��/�X����_TIME��^���  ��GDEB�UG\�˴�GINP_FLMSK�����Tfp����PGA�  ����)CH�����TYPE���������� � -?hcu �������/ /@/;/M/_/�/�/�/ �/�/�/�/�/??%?�7?`?��WORD �?	=	RS�fu	PNSU�Ԝ2JOK�DRT�Ey�]TRACE�CTL 1x3���� �`: ;&�`�`�>�6_DT Qy3�%@��0D � [ `2@,6DU-6D.6D/6D06D16A�c2@�`8B V�8BR�8BM 8BJ�8BTF�8B6D6D	6DU
6D6D6D6DE6D6D^�8B6DU6D6D6D6D�8B6D6D~P8BA6DV�8Bj�8B6DA6DҀ8B�8B!6DE"6D#6D�8B%6DU&6D'6D(6D)6D*6D5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m�� ������Ǐن.A�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� r�����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ����������� �*��$PGT�RACELEN � )�  ���(��>�_�UP z��e�m�u�Y�n��>�_CFG {�m�W�(�n����PКӂ�DEFS_PD |���a�P��>�IN��T_RL }��(��8����PE_CO�NFI��~m�'�mњ��ղ�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�p�ح֚��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P;t _��������  Dz (�
 H�X~i�� ����/�/D/�//h/S/�/��
V�7.10beta�1��  A��E�"ӻ�Ay (�� ?!G��!/>���"����!����!BQ��!A\� �!���!2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?OO :O%O7OpO[O�OO�O �O�O�O�O_�O6_!_ Z_E_~_i_�_�_�_�_ �_�_'o2o�_VoAo So�owo�o�o�o�o�o �o.R=v1�<�/�#F@ �y�} ��{m��y=��1� '�O�a��?�?�?���� ��ߏʏ��'��K� 6�H���l�����ɟ�� �؟�#��G�2�k� V���z��������o ��ίC�.�g�R�d� ���������п	��� -�?�*�cώ���� �������B�;� f�x�������DϹ��� ���������7�"�[� F�X��|������� ����!�3��W�B�{� f��������� ��� ��/S>wbt ������ =OzόϾψ��� �ϼ� /.�'/R�d� v߈߁/0�/�/�/�/ �/�/�/#??G?2?k? V?h?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O���O�O�O_ _?_*_c_N_�_r_�_ �_�_�_�_o�_)oT fx�to���/ �o/>/P/b/t/ mo�|���� ���3��W�B�{� f�x�����Տ����� ��A�S�>�w�b��� �O��џ������+� �O�:�s�^������� ͯ���ܯ�@oRodo �o`��o�o�o��ƿ�o ���*<N�Y�� }�hϡό��ϰ����� ���
�C�.�g�Rߋ� v߈��߬�����	��� -��Q�c�N�ﲟ�� ��l��������;� &�_�J���n������� ����,�>�P�:L ����������� �(�:�3��0iT �x�����/ �///S/>/w/b/�/ �/�/�/�/�/�/?? =?(?a?s?��?�?X? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O*\&_8_r���_�_��$PL�ID_KNOW_�M  ��� Q�TSV ����P��?o"o4o�O�XoCoUo�o R�SM_GRP 1��Z�'0{`�@�`uf�e�`
�5� �g pk'Pe ]o�����������SMR�c�b�mT�EyQ}? yR ����������폯��� ӏ�G�!��-����� ������韫���ϟ� C���)���������`��寧���QST�a�1 1��)��v�P0� A 4� �E2�D�V�h������� ߿¿Կ���9��.� o�R�d�vψ��ϬϾϔ���2�0� Q�<3��3�/�A�S��4l�~ߐߢ��A5���������6
��.�@��7Y�k�}����8���������MAD  �)��PARNU/M  !�}o+���SCHE� S�
���f���S��UPD�f�x��_C�MP_�`H�� �'��UER_CHK-���ZE*�<RSr��_�Q_M�OG���_�X�__RES_G��!� ��D�>1bU �y�����/ �	/����+/ �k�H/g/l/��Ї/ �/�/�	��/�/�/� X�?$?)?���D?c?�h?����?�?�?�V� 1��U�ax�@c�]�@t@(@c�\�@�@D@c�[�*@��THR_INRr�J�b�U�d2FMASS?O �ZSGMN>OqCMO�N_QUEUE ���U�V P~P *X�N$ UhN�FV��@END�A��IEcXE�O�E��BE�@|�O�COPTIO�G���@PROGRAoM %�J%�@��?���BTASK_�IG�6^OCFG ���Oz��_�PDA�TA�c��[@Ц2=�DoVohozo�j 2o�o�o�o�o�o�);M jINFO
[��m��D�� ������1�C� U�g�y���������ӏ����	�dwpt�l �)�QE DIT ���_i��^WER�FLX	C�RGA�DJ �tZAЄ����?נʕFA��I�ORITY�GW�>��MPDSPNQ�����U�GD��OT�OE@1�X� _(!AF:@E� �c�Ч!tcp|n���!ud��>��!icm���?n<�XY_�Q�X�{��Q)� *�1�5��P��]�@� L���p��������ʿ ��+�=�$�a�Hυ�z��*��PORT)Q�H��P�E��_CARTREPP|X��SKSTA�H^�
SSAV�@�tZ�	2500H8�63���_x�
�'��*X�@�swPtS��ߕߧ���URGE��@B��x	WF��DO�F"[W\��������WRUP_DE?LAY �X��ԟR_HOTqX	B%��c���R_NOR�MALq^R��v�S�EMI�����9�Q�SKIP'��tUr�x 	7�1�1� �X�j�|�?�tU���� ����������$ J\n4���� ����4FX |j����� ��/0/B//R/x/�f/�/�/�/tU�$R�CVTM$��D��� DCR'����Ў!C`N�C��d�C��o?���>��L<|��{:��g�&���/���%��t����|���}'�:�o?�� �<
6b<߈�;܍�>u.��?!<�& �?h?�?�?�@>��?O  O2ODOVOhOzO�O�O �O�O�O�?�O�O__ @_+_=_v_Y_�_�_�? �_�_�_oo*o<oNo `oro�o�o�o�_�o�o �o�o�o8J-n ��_������ �"�4�F�X�j�U�� ����ď���ӏ�� �B�T��x������� ��ҟ�����,�>� )�b�M����������� �ïկ�Y�:�L�^� p���������ʿܿ�  ����6�!�Z�E�~� ��{ϴϗ�����-��  �2�D�V�h�zߌߞ� ����������
���.� �R�=�v��k��� �������*�<�N� `�r������������ ����&J\? �������� "4FXj|���!GN_ATC �1�	; �AT&FV0E0��ATDP/6/9/2/9��ATA�,�AT%G1%B�960�++U+�,�H/,�!�IO_TYPE � �%�#t�R�EFPOS1 1}�V+ x�u/�n�/j�/
=�/ �/�/Q?<?u??�?4?�?X?�?�?�+2 1�V+�/�?�?\O�?x�O�?�!3 1�O�*O<OvO�O�O_�OS4 1��O�O�O_��_t_�_+_S5 1�B_T_f_�_o	oBo>�_S6 1��_�_��_5o�o�o�oUoS7 1�lo~o�o�oH�3l�oS8 1� %_����SMASK 1��V/  
?�M��XNOS/�r�����~�!MOTE  n���$��_CFG ᢫��q���"PL_�RANG�����POWER ������SM_DRYPRG %o��%�P��TART� ��^�UME_PRO-�?����$�_EXEC_EN�B  ���GS�PD��Րݘ��T3DB��
�RM�
��MT_'�T�����OBOT_NA_ME o�����OB_ORD_�NUM ?��b!H863�  �կ����PC_TIMoEOUT�� x�oS232Ă1��� LTEA�CH PENDA1N��w��-���Mainte�nance Co#ns���s�"���?KCL/Cm��
�
���t�ҿ ?No Use-��8Ϝ�0�NPO�򁮋���.�C7H_L������q�	��s�MAVA#IL�����糅���SPACE1 2��, j�߂�D��s�߂� �{S�?8�?�k�v� k�Z߬��ߤ��ߚ�  �2�D���hߊ�|�� `����������  �2�D��h��|����`���������y���2����0�B���f� ����{���3);M_ ������/� /44FXj| */���/�/�/?(??=?5Q/c/u/�/ �/G?�/�/�?O�?$OEO,OZO6n?�?�? �?�?dO�?�?_,_�O A_b_I_w_7�O�O �O�O�O�_�O_(oIo@o^oofo�o8�_ �_�_�_�_�oo6oE�f){���Gw �o� �:��
M� ��� *�<�N�`�r������� w���o�収���d.��%�S�e�w��� ��������Ǐَ��� Θ8�+�=�k�}����� ��ůׯ͟����%� '�X�K�]��������� ӿ������#�E��W� `� @ �������x�����\�e����������� R�d߂�8�j߬߾߈� �ߤ����������0� r���X�������@������8����
�����_MODE � �{��S �"�{|�2�0��ψ��3�	S|)CWORK_AD���X9(+R  ��{�`� �� _?INTVAL���d����R_OPTI[ON� ��H �VAT_GRP �2��up#(N�k| ��_����� /0/B/��h�u/T�  }/�/�/�/�/�/�/? !?�/E?W?i?{?�?�? 5?�?�?�?�?�?O/O AOOeOwO�O�O�O�O UO�O�O__�O=_O_ a_s_5_�_�_�_�_�_ �_�_o'o9o�_Iooo �o�oUo�o�o�o�o�o �o5GYk-� ��u����� 1�C��g�y���M��� ��ӏ叧�	��-�?� Q�c������������ ���ǟ�;�M�_�����$SCAN_GTIM��_%}��R �(�#(�(�<04+d d 
!AD�ʣ��u�/X�����U��25�����dA�8�H�g��]	����������dd�x�  P~���� ��  8� ҿ�!���D��$�M�_�q� �ϕϧϹ��������8ƿv��F��X��/� ;�o�b��pm��t�_DiQ̡  � l�|�̡ ĥ�������!�3�E� W�i�{�������� ������/�A�S�e� ]�Ӈ����������� ��);M_q ������� r���j�Tfx� ������// ,/>/P/b/t/�/�/�/p�/�/�%�/  0�� 6��!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O *�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo �O�OJ�o�o�o�o�o �o�o 2DVh z�������
�7?  ;�>�P� b�t���������Ǐُ ����!�3�E�W�i��{�������ß � ş3�ܟ��&�8�J��\�n�������������ɯ����,�� �+�	12�345678��W 	� =5���@f�x���������� ���
��.�@�R�d� vψϚ�៾������� ��*�<�N�`�r߄� �Ϩߺ��������� &�8�J�\�n�ߒ�� �����������"�4� F�u�j�|��������� ������0_�T fx������ �I>Pbt �������! /(/:/L/^/p/�/�/ �/�/�/�/�2�/�?�#/9?K?]?�i�Cz  Bp˚ /  ��h2��*��$SCR_GR�P 1�(�U8�(�\x�d�@ � ��'�	 ?�3�1 �2�4(1*�&�I3�Fp1OOXO}m��CD�@�0ʛ)���H�UK�LM-10�iA 890?�9�0;��F;�M61�C D�:�CP��1

\&V�1	�6F� �CW�9)A7Y	(R�_��_�_�_�_�\���0i^�oOUO>o Po#G�/���o'o�o��o�o�oB�0ƐrtAA�0* C @�Bu&Xw?���ju�bH0{UzAF?@ F�`�r� �o�����+�� O�:�s��mBqrr����������B�͏b�� ��7�"�[�F�X���|� ����ٟğ���N��� AO�0�B�CU
L���xE�jqBq>HE����$G@�@pϯ BȆ��G�I
E�0E�L_DEFAUL�T  �T���E��MI�POWERFL � 
E*��7�WF�DO� *��1E�RVENT 1����`(�� L�!DUM_EI�P��>��j!AF_INE�¿C�O!FT�����r�!o:� ���a�!RPC_M'AINb�DȺPϭ�Nt�VIS}�Cɻ�����!TP��PU��ϫ�d��E�!
P�MON_PROX	YF߮�e4ߑ��_��f����!RD�M_SRV�߫�g��)�!R�IﰴYh�u�!
v�M���id���!RL�SYNC��>�8|���!ROS��4��4��Y�(�}��� J�\����������� ��7��["4F� j|����!��Eio�ICE_�KL ?%� �(%SVCPRG1n>���3��3���4//�5./3/�6V/[/��7~/�/��D�/�9�/�+�@��/�� #?��K?��s?�  /�?�H/�?�p/�? ��/O��/;O��/ cO�?�O�9?�O� a?�O��?_��?+_ ��?S_�O{_�)O �_�QO�_�yO�_� �Os����>o�o }1�o�o�o�o�o�o�o ;M8q\� �������� 7�"�[�F��j����� ��ُď���!��E� 0�W�{�f�����ß�� �ҟ���A�,�e� P���t��������ί��y_DEV ���MC:��@`!�OU�T��2��RE�C 1�`e�j�{ �� 	 � ����˿���ڿ��
 �`e���6�N� <�r�`ϖτϦ��Ϯ� ������&��J�8�n� ��bߤߒ��߶����� ��"��2�X�F�|�j� ������������� �.�T�B�x�Z�l��� ����������, P>`bt��� ���(L: \�d�����  /�$/6//Z/H/~/ l/�/�/�/�/.��/? �/2? ?V?D?f?�?n? �?�?�?�?�?
O�?.O @O"OdORO�OvO�O�O �O�O�O�O__<_*_ `_N_�_�_x_�_�_�_ �_�_oo8oo,ono \o�o�o�o�o�o�o�o �o "4jX� �������� �B�$�f�T�v����� �������؏��>��,�b�P�r���p�V [1�}� P
�6!����� �#<��TYPE\���HELL_CFG� �.��� � 	�����RSR������ӯ���� ���?�*�<�u�`�������������� ����%�3�E�(�Q���ӐM�o¦p��d��2Ӑd�]�K�:�HK 1�H� u������ �A�<�N�`߉߄ߖ� ������������&��8��=�OMM �H���9�FTOV�_ENB&���1�O�W_REG_UI����IMWAITr��a���OUT������TIM��;���VAL����_UNIT��K�1��MON_ALIA�S ?ew� ( he�#�������� ��Ӕ��);M�� q����d�� %�I[m �<������ !/3/E/W//{/�/�/ �/�/n/�/�/??/? �/S?e?w?�?�?F?�? �?�?�?�?O+O=OOO aOO�O�O�O�O�OxO �O__'_9_�O]_o_ �_�_>_�_�_�_�_�_ �_#o5oGoYokoo�o �o�o�o�o�o�o 1C�ogy��H ����	��-�?� Q�c�u� �������Ϗ Ꮜ���)�;��L� q�������R�˟ݟ� ����7�I�[�m�� *�����ǯٯ믖�� !�3�E��i�{����� ��\�տ�����ȿ A�S�e�wω�4ϭϿ� ���ώ����+�=�O� ��s߅ߗߩ߻�f��� ����'���K�]�o� ���>��������� �#�5�G�Y��}���������n��$SM�ON_DEFPR�O ������ �*SYSTEM*�  d=��RECALL ?}��� ( �}/x�copy fr:�\*.* vir�t:\tmpba�ck7=>ins�piron:12732 Ybt�.� }0.a6H@Z_��4/�s:orderf?il.dat�Mpbt�� }+/mdb:�MZ� �/�-�Qb/t/ �/�/�</�a/�/? ?);��/p?�?�? ���]?�? OO%/ �/�/[/lO~O�O�/�/ FO�/�O�O_!?3?�? W?h_z_�_�?�?L_�? �_�_
oO/O�OSOdo vo�oo�O>o�O�o�o +_=_�_�or� ��_D�__��� 'o�o�o]on������o�6�H��o������
�xyzrate 61 ��ˏݏn���䒟��.�M�4804 H�Z�������3.@��a�s�������*�I���Y�������..�A���ݯn� ����%���G�đ^�� ��&�8���ܯm�� �Ϥ���ȯZ������ "�4�ǿX�i�{ߍߠ� ��C�ֿ������0� B�T�e�w��Ϯ�I� ��������,߿�P� a�s�������;���`� ��(�������o0����M�28ǟY ��!�3��a s����E�Y� �/!�3�F��n/ �/�/��6/H/� ^/�/ ??&8��m?? �?���Z?�?�?O�!w�$SNPX_�ASG 1�����9A�� P 0 '�%R[1]@1�.1O y?�#s% dO�OsO�O�O�O�O�O �O __D_'_9_z_]_ �_�_�_�_�_�_
o�_ o@o#odoGoYo�o}o �o�o�o�o�o�o* 4`C�gy�� �����	�J�-� T���c�������ڏ�� ���4��)�j�M� t�����ğ������ݟ �0��T�7�I���m� �������ǯٯ��� $�P�3�t�W�i����� ���ÿ����:�� D�p�Sϔ�wω��ϭ� �� ���$���Z�=� dߐ�sߴߗߩ����� �� ��D�'�9�z�]� ���������
��� �@�#�d�G�Y���}� ������������* 4`C�gy�� ����	J- T�c����� �/�4//)/j/M/ t/�/�/�/�/�/�/�/�?0?4,DPARAoM �9ECA_ �	��:P�4��0$HOFT_�KB_CFG  �p3?E�4PIN_�SIM  9K��6�?�?�?�0,@RV�QSTP_DSBº>�21On8J0SR� ��;� & �MULTIROBOTTASK=O�p3�6TOP_�ON_ERR  ��F�8�APTN ��5�@�A�BRING_P�RM�O J0VD�T_GRP 1�<Y9�@  	�7n8 _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D khz����� ��
�1�.�@�R�d� v���������Џ��� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\��������� ��ȯگ����"�I� F�X�j�|�������Ŀ ֿ����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�a�^�p��� ��������� �'�$� 6�H�Z�l�~���������������3VPRG�_COUNT�6q��A�5ENB�O�M=�4J_UP�D 1��;8  
p2���� �� )$6Hq l~�����/ �/ /I/D/V/h/�/ �/�/�/�/�/�/�/!? ?.?@?i?d?v?�?�? �?�?�?�?�?OOAO <ONO`O�O�O�O�O�O �O�O�O__&_8_a_�\_n_�_�_�_YS�DEBUG" � ��Pdk	�PSP_PwASS"B?�[�LOG ���m�P�X�_ � �g�Q
MC�:\d�_b_MPACm��o�o�Qa��o �vfSAV ��m:dUb�U�\gSV�\TEM�_TIME 1��� (�`ųS��2o	T1SVGgUNS} #'k��spASK_OPTION" �go�spBCCFG 3��| �b�{�}`����a&� �#�\�G���k����� ȏ������"��F� 1�j�U���y���ğ�� �ӟ���0��T�f��UR���S���ƯA� ����� ��D��nd� �t9�l���������ڿ ȿ�����"�X�F� |�jϠώ��ϲ����� ����B�0�f�T�v� xߊ��ߦؑ������ �(��L�:�\��p� ����������� � 6�$�F�H�Z���~��� ����������2  VDzh���� �����4Fd v������ //*/�N/</r/`/ �/�/�/�/�/�/�/? ?8?&?\?J?l?�?�? �?�?�?�?�?�?OO "OXOFO|O2�O�O�O �O�OfO_�O_B_0_ f_x_�_X_�_�_�_�_ �_�_oooPo>oto bo�o�o�o�o�o�o�o :(^Lnp �����O��$� 6�H��l�Z�|����� Ə؏ꏸ����2� � V�D�f�h�z�����ԟ ����
�,�R�@� v�d���������ίЯ ���<��T�f��� ����&�̿��ܿ�� &�8�J��n�\ϒπ� �Ϥ����������4� "�X�F�|�jߌ߲ߠ� ����������.�0� B�x�f��R������� �����,��<�b�P� ������x��������� &(:p^� ������  6$ZH~l�� ������/&/D/ V/h/��/z/�/�/�/��/�&0�$TBC�SG_GRP 2���%� � �1 
 ?�  /?A?+?e? O?�?s?�?�?�?�?�;�23�<d,� �$A?1	 H�C���6>���@E�5CL  B�p'2^OjH4J��B�\)LFY  A��jO�MB��?�IBl�O�O�@�JG_�@�  D	�15_ __$YC-P{_F_`_j\	��_�]@0�>�X�U o�_�_6oSoo0o~o�o�k�h�0	�V3.00'2	�m61c�c	*`�`�d2�o�e>�JC20(�a�i ,p�m�-  �0�����omvu1JCFG� ��% 1 �#0vz��rBrv�x����z � �%��I�4�m�X� ��|��������֏� ��3��W�B�g���x� ����՟������� �S�>�w�b�����'2 A ��ʯܯ������ E�0�i�T���x���ÿ տ翢����/��?� e�1�/���/�ϜϮ� �������,��P�>� `߆�tߪߘ��߼��� �����L�:�p�^� ������������  �6�H�>/`�r���� ������������  0Vhz8��� ���
.�R @vd����� ��//</*/L/r/ `/�/�/�/�/�/�/�/ �/?8?&?\?J?�?n? �?�?�?�?���?OO �?FO4OVOXOjO�O�O �O�O�O�O__�OB_ 0_f_T_v_�_�_�_z_ �_�_�_oo>o,obo Poroto�o�o�o�o�o �o(8^L� p������� $��H�6�l�~�(O�� ��f�d��؏���2�  �B�D�V�������n� ���ԟ
���.�@�R� d����v�������� Я���*��N�<�^� `�r�����̿���޿ ��$�J�8�n�\ϒ� �϶Ϥ�������ߊ� (�:�L���|�jߌ߲� �����������0�B� T��x�f������ �������,��P�>� t�b������������� ��:(JL^ ������ � 6$ZH~l� �^���dߚ // D/2/h/V/x/�/�/�/ �/�/�/�/?
?@?.? d?v?�?�?T?�?�?�? �?�?OO<O*O`ONO �OrO�O�O�O�O�O_ �O&__6_8_J_�_n_ �_�_�_�_�_�_�_"o oFo��po�o,oZo �o�o�o�o�o0 Tfx�H��� ����,�>��b� P���t���������Ώ ��(��L�:�p�^� ������ʟ���ܟ�  �"�$�6�l�Z���~� ����دꯔo��&� ЯV�D�z�h������� Կ¿��
��.��R��@�v�dϚτ�  ���� ��������$TBJOP_�GRP 2ǌ���  �?�������������x�JBЌ��9� �< �X�ƞ�� @���	� �C�� t�b�  C����>ǌ�͘Րդ�>���йѳ33=��CLj�fff?>��?�ffBG���Ќ�����t�ц�>;�(�\)�ߖ��E噙�;��h{CYj��  @h�~�B�  A�����f��C�  D�hъ�1��O��4�N����
:�/��Bl^��j�i��l�l����Aə�3A�"��D���Ǌ=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������<$�6�>B�\��T����Q�tsx�@g33@���C����y�1����>��Dh����������O<{�h�@i�  ��t��	� ��K&�j� n|���p�/��/:/k/�ԇ����!��	V3.0}0J�m61cIԃ*� IԿ��/�'� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�I�!CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;��;Q�UT,8�4` *���?�2���3\�X/�O��ESTPAR�S  ��	���H�R@ABLE 1%����0��
H�7Q 8��9
G
H
H�����
G	
H

H�
HYE��
H
H:
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_�^:BS _� �JGoYo ko}o�o�o�o�o�o�o �o1CUgy ����`#oRL�y�_ �_�_�_�O�O�O�O�O�X:B�rNUM  ����P���� V@P:B_CF�G ˭�Z�h�@���IMEBF_T�T%AU��2@�VE�RS�q��R {1���
 (�/����b� ����J� \���j�|���ǟ��ȟ ֟�����0�B�T�@��x�������2�_����@�
��MI_�CHAN�� � >��DBGLV����������ETHE�RAD ?��
O�������h������ROUT�!���!������SN�MASKD��U�255.���#������OOLOFS_�DI%@�u.�OR�QCTRL � ����}ϛ3rϧϹ��� ������%�7�I�[��:���h�z߯�APE?_DETAI"�G��PON_SVOF�F=���P_MON� �֍�2��S�TRTCHK ��^�����VTCOMPAT��O������FPROG �%^�%MULTIROBOTTݱx���9�PLAY&H���_INST_M�ް ������US8�q��LCK���QUICKME��=���SCREZ�}G�tps� @���u�z����_���@@n�.�SR_GR�P 1�^� �O����
��@+O=sa�� ��
m������ L/C1gU� y�����	/��-//Q/?/a/�/	1234567�0h�/�/@Xt�1����
 �}ipn�l/� gen.htm�? ?2?D?V?�`Panel� setupZ<}�P�?�?�?�?�?�? �??,O>OPObOtO �O�?�O!O�O�O�O_ _(_�O�O^_p_�_�_ �_�_/_]_S_ oo$o 6oHoZo�_~o�_�o�o �o�o�o�oso�o2D Vhz�1'� ��
��.��R�� v���������ЏG����UALRM��G ?9� �1�#� 5�f�Y���}������� џן���,��P���SEV  �����ECFG C��롽�A���   BȽ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �(�� ��3�/SOFTPAR�T/GENLIN�K?curren�t=editpa7ge,��,1���8!�3��� �����menu��962 �߆����K�]�o�36u�
��.�@��� W�i�{���������R� ����/A��e w����N�� +=O�s� �������f�� f//'/9/K/]/` �/�/�/�/�/�/j/�/ ?#?5?G?Y?�/�/�? �?�?�?�?�?x?OO 1OCOUOgO�?�O�O�O �O�O�OtO�O_-_?_ Q_c_u__�_�_�_�_ �_�_��)o;oMo_o qo�o�_�o�o�o�o�o �o%7I[m � ������ �3�E�W�i�{���� ��ÏՏ������� A�S�e�w�����*��� џ�����ooO� a�s���������ͯ߯ ���'���K�]�o� ��������F�ۿ��� �#�5�ĿY�k�}Ϗ� �ϳ�B��������� 1�C���g�yߋߝ߯� ��P�����	��-�?� *�<�u������� ������)�;�M��� �������������l� %7I[�� �����hz !3EWi��� ����v////�A/S/e/P���$U�I_PANEDA�TA 1������!  	�}w/�/�/�/�/?? )?>?� �/i?{?�?�?�?�?*? �?�?OOOAO(OeO LO�O�O�O�O�O�O�O��O_&Y� b� >RQ?V_h_z_�_�_�_ _�_G?�_
oo.o@o Rodo�_�ooo�o�o�o �o�o�o*<#`@G��}�-\�v �#�_��!�3�E�W� �{��_����ÏՏ� ��`��/��S�:�w� ��p�����џ����� �+��O�a����� ����ͯ߯�D���� 9�K�]�o�������� ɿ���Կ�#�
�G� .�k�}�dϡψ����� ����n���1�C�U�g� yߋ��ϯ���4����� 	��-�?��c�J�� ������������ ��;�M�4�q�X���� �������%7 ��[������ �@��3W iP�t���� �/�//A/����w/ �/�/�/�/�/$/�/h ?+?=?O?a?s?�?�/ �?�?�?�?�?O�?'O OKO]ODO�OhO�O�O �O�ON/`/_#_5_G_ Y_k_�O�_�_?�_�_ �_�_oo�_Co*ogo yo`o�o�o�o�o�o�o �o-Q8u�O�O}��������)�>��U-�j� |�������ď+��Ϗ ���B�)�f�M��� �����������ݟ��&�S�K�$UI_�PANELINK� 1�U�  �  ���}1234567890s����� ����ͯդ�Rq���� !�3�E�W��{����� ��ÿտm�m�&����Qo�  �0�B� T�f�x��v�&ϲ��� ������ߤ�0�B�T� f�xߊ�"ߘ������� ���߲�>�P�b�t� ���0��������� ���$�L�^�p����� ,�>������� $�0,&�[gI� m������ �>P3t�i� �Ϻ� -n��'/ 9/K/]/o/�/t�/�/ �/�/�/�/?�/)?;? M?_?q?�?�UQ�= �2"��?�?�?OO%O 7O��OOaOsO�O�O�O �OJO�O�O__'_9_ �O]_o_�_�_�_�_F_ �_�_�_o#o5oGo�_ ko}o�o�o�o�oTo�o �o1C�ogy �����B�	� �-��Q�c�F����� |�������֏�)� �M���=�?��?/ ȟڟ����"�?F� X�j�|�����/�į֯ �����0��?�?�? x���������ҿY�� ��,�>�P�b��� �Ϫϼ�����o��� (�:�L�^��ςߔߦ� ��������}��$�6� H�Z�l��ߐ����� ����y�� �2�D�V� h�z����-������� ��
��.RdG ��}����c� ��<��`r�� ������//&/ 8/J/�n/�/�/�/�/ �/7�I�[�	�"?4?F? X?j?|?��?�?�?�? �?�?�?O0OBOTOfO xO�OO�O�O�O�O�O _�O,_>_P_b_t_�_ _�_�_�_�_�_oo �_:oLo^opo�o�o#o �o�o�o�o ��6 H�l~a��� �����2��V� h�K�������1� U
��.�@�R�d�W/ ��������П����� �*�<�N�`�r��/�/ ?��̯ޯ���&� ��J�\�n�������3� ȿڿ����"ϱ�F� X�j�|ώϠϲ�A��� ������0߿�T�f� xߊߜ߮�=������� ��,�>���b�t�� ����+���� ��:�L�/�p���e��� �������� ��6����ۏ��$U�I_QUICKM�EN  ����}��RE�STORE 1����  �
�8m3\n���G ����/�4/F/ X/j/|/'�/�/�// �/�/??0?�/T?f? x?�?�?�?Q?�?�?�? OO�/'O9OKO�?�O �O�O�O�OqO�O__ (_:_�O^_p_�_�_�_ QO[_�_�_I_�_$o6o HoZoloo�o�o�o�o �o{o�o 2D�_ Qcu�o���� ���.�@�R�d�v���������Џ⏜S�CRE� ?��u1sc� �u2�3�4�5*�6�7�8���USER����TL���ks'���4��U5��6��7��8���� NDO_CFG� ڱ  �  �� PDATE �h��No�ne�SEUFR�AME  �ϖ��RTOL_A�BRT����EN�B(��GRP 1���	�Cz  A�~�|�%|�������į֦��X�� �UH�X�7�MSK � K�S�7�N��%uT�%�����V�ISCAND_M;AXI�I�3����FAIL_IMG�I�z �% #S���IMREGNUMI�9
���SIZI�� ��ϔ,�ONOTMOU'�K�Ε��&����a���a��s��FR:\�� � MC:\(��\LOGh�B@Ԕ !{��Ϡ������z MCyV����UD1 ֓EX	�z ��POO64_�Q���n6��PO!�L!I�Oڞ�e�V�N��f@`�I�� =�	_�SZVmޘ���`�WAImߠ�S?TAT �k�% !@��4�F�T�$#�x���� �2DWP  ?��P G��=��͎����_JMPERR �1ޱ
  �p2�345678901���	�:�-�?� ]�c������������������$�MLOWp�ޘ�����_TI/��˘'��MPHA�SE  k�ԓ|� ��SHIFT%�k1 Ǚ��< z��_���� F/|Se�� �����0/// ?/x/O/a/�/�/�/�/�/����k�	V�SFT1\�	V:��M+3 �5�Ք� p����A�  �B8[0[0�Πp�g3a1Y2�_3Y�7ME��K�͗	6e���W&%��M����b��	��$��TDINEND3�4��4AOH�+�G1�OS2O�IV I���]LRELEvI��4.�@�~�1_ACTIV�IxT��B��A �m�0�/_��BRDBГO�Z�YBOX �Xǝf_\��b�2�T�I190.�0.�P83p\N�V254p^�Ԓ�	 �S�_�[b���robot�84q_   �p�9o\�pc �PZoMh�]Hm�_Jk@1��o�ZABCd��k�,���P\�Xo}�o 0);M�q� �������>��aZ�b��_V