��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG(�ET�H_FLTR.�  $� �  �FTP�_CTRL. �@ $LOG_�8	�CMO>$�DNLD_FIL�TE� � SUBD�IRCAP� o �HO��NT.� 4� H_NA�ME !A?DDRTYPA �H_LENGTH�' �z +L�S D $?ROBOTIG �PEER^� MA�SKMRU~O�MGDEV#����RDM*�DI�SABL&�T�CPIG/ 3 $ARPSIZ&�_IPF'W_�MC��F_IN�� FA~LASS�s�HO_� IN{FO��TELKG PV�b�	 WORD  �$ACCESS�_LVL?TIM�EOUTuORT� � �ICEUS�= ��$#  ����!�� � �� VIRTUAL��/�!'0 �%�
���F����l�$�%���+g �����$�� �-2%;�SHA�RED 1�)  P!�!�?���!|?�?�?�?�?O �?%O�?1OOZOOBO �OfO�O�O�O�O_�O �OE__i_,_�_P_�_ t_�_�_�_o�_/o�_ SooLo�oxo�opo�o �o�o�o�o*O s6�Z�~�� ���9��]� ��� D�V���z�ۏ���� #���Y�H�}�@����)7z _LIST �1=x!1."ܒ0��d�ە1�d�255.$������%ړ2��X� ��+�=�O�3Y��@Р�������O�4ѯ��H���	��-�O�5 I����o�������O�6���8������ �$���-� � ��-��%�%��&!Òu�)�0H!� ����rj3_'tpd���! � �!!KC� e�0�x���&W�!Cm ��w߉�S�!C�ON� ��1�=�s'mon��W�