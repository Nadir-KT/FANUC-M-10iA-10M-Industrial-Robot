��   ��A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����DRYRUN�_T   � �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L � &&J_ � 4 $T�YPENFST_�IDX��_IC�I �MIX�_BG-�� G�_NAMc %$gMODc_USd~CIFY_TI<� #MKR-�  $LIN�c   x_S�IZa#� . � $USE_FLGA�l�i�SIMA�Q��QB�SCAN�RAX�IN�I���_COUNrR�O�_!_TMR�_VA�gy h>�i�p'` ���H�!^%�$$�CLASS  O����!��5��}5� VIRTUR �/� '/ �%�5��������8� �!2�%I1�+�M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmO��+6W�?�%�! ����O�O�O  �10� ' 1=�+ 4%zO*_��11_]_<_�_ �_r_�_�_�_�_�_�_ #oooYo8oJo�ono�1�C���-54`�� �b1�d,1 �!�a�o.@Rd v������� ?~c�a1&�8�J�\� n���������ȏڏ�`����!�C�1�) U�g� y���������ӟ��� 	��-��G�`�r��� ������̯ޯ��� &�8�C�\�n������� ��ȿڿ����"�4� F�Q�j�|ώϠϲ��� ��������0�B�M� _�xߊߜ߮������� ����,�>�P�[�t� ������������ �(�:�L�^�i���� ���������� $ 6HZe�w���� ���� 2D Vh�F