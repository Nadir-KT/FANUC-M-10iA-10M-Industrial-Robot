��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ����ALRM_�RECOV1   $ALMO�ENB��]ON�i�APCOUPwLED1 $[�PP_PROCE�S0  �1�� GPCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y12 � u3�|4|GRG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WAx�471�:OFF_ �N�3DELHLO�Gn25Aa2?i1@N?�� -M���AW+0�$�Y $DB� 6CkOMW!2MO� �21H _A.	 \vrVE�1$F��A{$O��D�B~�CTMP1_F�E�2�G1_�3�B�2��GXD�#
 �d $CARD�_EXIST4�$FSSB_TY�PuAHKBD_YS�B�1AGN Gn� $SLOT�_NUMJQPREV,DBU� g1G �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��AETE_OK�RUS�P_CR�Q$;4�V� 0LACIw1�RAP�k �1x@ME@$D�V�Q�Pv�Ah{oQL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa�!ip;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I�9�TY�D,P*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6��U7��8��94�qO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS�`�}Aw��"�tP_*0wOFSzR @� �RO_K8���aIT<�3��NOM_�0�1�ĥ34 ��T !�� $���AxP��K}EX�� �0g0I01�<�p�
$TFa��Co$MD3��TO�3��0U� �� R�Hw2�C1|�EΡg0wE{vF�vF�C��p@�a2 
P$A`PU�3N�)#�dR*�AX��!sDETAI�3B�UFV��p@1 �|�p۶�pPIdTV� PP[�MZ�Mg��Ͱj�F[�SIMQ�SI�"0��A.������lw Tp|zM��P�B�FACTrbHPEW7�P1Ӡؖ�v��MCd�5 �$*1JB�p<�*1DECHښ�H��|(�c� � +P�NS_EMP��#$GP���,P_��3d�p�@Pܤ��TC�� |r��0�s��b�0�� `�B���!
���JR� ���SEGFR��ITv �aR�TkpN&S�,�PVF4��� &k�Bv�u�c u��aE�� !2��+�MQ��E�SIZ�3��䂖�T��P�����aRSINF�����kq@��������LX�8����F�CRCMu�3CClpG��p���O} ���b�1�������2�*V�DxIC��C���r�����P��{� EVT �zF_��F�p)NB0�?������A�! �r�Rx ����V�lp�2��aR��t�,�g��RTx #�5�5"2���uAR���`CX�$L	G�p��B�1 `s�P��t�aA�0{�У+0R���tME�`!Bu�pCrRA 3tAZЪл�pc�OT�FC�b�`�`FNp���1��ADI+�a%� �b�{��p$�pSp�c��`S�P��a,QMP$6�`Y�3��M'�p�U��aU  $.>�TITO1�S�S��!��$�"0�DBP�XWO��!���$SK��2�DBd�"�"@�PR8� 
� ���#� >�q1$��)$��+�L9$?(ӤV�%@?R4C&�_?R4ENE��1'~?(�� RE�pY2�(H �OSn��#$L�3$$3�R��;3�MVOk_9D@!V�ROScrr��w�S���CRIGGER2FPA�S��7�ETURN0B�cM[R_��TUː[��0EWM%���G1N>`��RLA���E�ݡ�P�&$PD�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWAY�RMO#�aw!��DCS_)  `IS#� ��� �s3S�AQ汯  4Rx�ZSW�AQ�p�@1U9W��cTNTV)�5RV
a���|c�éWƃ¤�JB��x0��SAsFEۥ�V_SV�b�EXCLUU�;�N�ONL��cYg��~az�OT�a{�HI�_V? ��R, M�_G *�0� ��_z��2� �CdSGO  +�rƐm@�A@�c~b���w@��V�i|�b�fANNUNx0,�$�dIDY�UABc�@Sp�i�a+ �j�fs�'P�pOGIx2,��$F�b�$ѐ�OT�@A $DUMMY��Ft���Ft±� 6U- 7` !�HE�|s��~bc�B@ SUF�FI��4PCA*�Gs5Cw6Cq�DMSWU. 8���KEYI��5�T�M�1�s�qoA�vIN�ޱw�ib, / D���HOST�P! 4���<���<�°<��p�<�EM'���Z�� S�BL� UL��0  �	��E�� �T�01 � �$��9USAMPL�о�/���決�$ I�@갯 $SUB ӄ��w0QS�����#��SAV�����c�S�< 9�`�fP$�0E�!� YN_B�#2� 0��DI�d�pO�|�m��#$F�R_�IC� �ENC�2_Sd3  ��< 3�9���� cgp����4�"��2�rA��ޖ5�� �`ǻ�@Q@K&D-!<�a�AVER�q�����DSP
���PC_�q��"�|�ܣ�oVALU3�HE��(�M�IP)���OkPPm �THЈ*��S" T�/�Fb�;�d����d D�pѼ�16 H(rLL_DUǀ�a�@��0k���֠OT�"U��/���"@@NOAUkTO70�$}�Hx�~�@s��|�C� ���C� 2v�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3*T�3a�3n�4|�q8���9 <���z�ΓKI����H硵�BaFEq@{@: y,��&a? PF_P?��>�����E�@���!QQ��;�fp$TP�$�VARI����,�U�P2Q`< W�߃TD��g���`����������BAC�"= T2����$)�,+r³�p IFI��p��� q M�P"�l@``>>t ;��6����ST����@T��M ����0	�� i���F���������kR�t ����FORCE�UP�b܂FLUS

pH(N��� ��6b/D_CM�@E�7�N� (�v�P��REM� Fa��@(j���
K�	N����EFF/���@IN̆QOV��OV=A�	TROV �DT)��DTMX :e �P:/��Pq��vXpCLN _ �p��@ ��	_|���_T: �|�&PA�QDI���10��0�Y0RQm��_+qH���M���C9L�d#�RIV{�ϓnN"EAR/�IO�#PCP��BR��cCM�@N 1b 3�GCLF��!DY��(�q�#5T�D�G���� �%r�S9S� )�? P(q1�1�`_1"81�1�EC13D;5�D6�GRA���@������PW�ON<2EBUG�S�2�C`gϐ_E �A ��?����T�ERM�5B�5���'ORIw�0C�5���SM_-`���0D��6 �TA�9Eܽ5GP�UP��Fg� -QϒA�P|�3�@B$SEGGJv� EL�UUSEPNFI��pBx��1x@��4>DC$UF�P��$���Q�@C���G�0T�����SwNSTj�PATۡ<g��APTHJq�A�E*�Z%qB\`F�{E���F�q�pARxPY�aS�HFT͢qA�AX_�SHOR$�>��6 �@$GqPE���O#VR���aZPI@P@$�U?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi� [Y)��G�@R��i�e԰�i�R�!P�uAScYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UaP���P���WOR�@�M��u�GRSMT��G��GR��3�a�PA�@���p5�'�H� � j�A�T�OCjA7pP]Pp$OPd�O��C�%��p�O!��RE.pR�C�AO�?��Be5pR�EruIx'Q�G�e$PWR) IMdu�RR_$s��5�.�B Iz2H8�=��_ADDRH�H_LENG�B�q�q:��x�R��So�J.�SS��SK������ ��-�SE*���rmSN�MN1K	��j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ���p�Q� ��OUPW3��b_>�I��!q�a1 ��������|��� �����-���:���i+IOX2S=�D�e���^���L $x��p�!_OFF[r�_�PRM_�^�aTTP_�H��wM (�pOBJ�"l�pG�$H�LE�C���ٰN � \9�*�AB_�T��b
�S�`�S��LV���KRW"duHITC�OU?BGi�LO�q����d� Fp�k�GpSS� ���HQWh�wA��O.��`�INCPUX2VISIO��!��¢.��á<�á-� �IO�LN)�P 87�R�'�[p$SL�b�d PUT_��$�dp�Pz �� F�_AS2Q/�$ALD���D�aQT U�0�]P�A������PH�YG灱Z�̱5�UO� 3R `F���H�@Yq�Yx�ɱvpP�S�dp���x��ٷZ ��UJ��S����N�E�WJOG�G �DIS��r�KĠ��3T |��AV��`_��CTR!S^�FLA�Gf2r�LG�dU ��n�:��3LG_SIZ��ň��,=���FD��I���� Z �ǳ��0�Ʋ�@s�� -ֈ�-�=�-���-��0<-�ISCH_��DqR��N?���V��EAE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��OGB�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S S�n���_BUFF�1XY��PT�$�� �v��fĵ�1�A�rYY��P ���\��pOS1�2��3���_�0Z �  ��aiE�*�.�IDX�dP�RhraO�+��A&ST���R��Yz�<! Y$EK&CK+����Z&m&KF�1[ L ��o�0��]PL�6pwq��t^����w��7�_ \ �`��瀰��7��#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3b�DM�R7��LDR5<4R5ORG.���e2�(`���V�8.��T<�3�d^ �q�<4��-4R5S�`T00m��0�DFRCLMC�!D�?�?3I@��MI�C��d_ d���R�Qm�q�DSTB�	�  �Fg�HA�X;b �H�LEXGCESZrKrBMup
�a`��B;d��rB�`��`a��F_A@�J��$[�O�H0K�d�b \��ӂS�$M�B��LIБ}SREQUIR�R>q�\Á��XDEBU��oAL
� MP�c�ba��P؃4ӂ!BoAND���`��`d�҆�c�cDC1��IN�����`@��(h?Nz�@q��o���UPST8� en�rLOC�RI�p�EX�fA�p��A�oAODAQP�f �X��ON��[rMF �����f)�"I��%�e|��T�$�FX�@�IGG� g �q��"E�0��#���$R�a%;#7y��Gx�VvCPi�DATAw�pE:�y��RFЭ��NVh t $+MD�qIё)�v+�tń�tH�`�P�u�<|��sANSW}��t�?�uD�)DAp�`�	@Ði �@�CU��V�T0�A'��0RR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2N�RIN��v�<��'NTE���kE����,��b����_Nl@��ڂ��kDׄRm�7DIViFDH�@ـ:n�$V��'c!$���������~�0R�o�H �$BEL�Tb��!ACCEL�+��ҡ��IRC��t����T/!���$PS�@#2LP q�Ɣ83������� ��PATH��������3̒Vp�A_�Q�.��4�B�Cᐈ�_M=G�$DDQ���G�$FWh��p���m�����b�DE��P�PABNԗROTSPEED����00�J�Я8��@��P�$USE_��P���s�SY��c�A �>qYNu@Ag��OsFF�q�MOUN�3NGg�K�OL�H�INC*��a��q��Bxj�L@�BENCS���q�Bđ���D��IN�#"I̒��4�\BݠV�EO�w�Ͳ23_UyPE�߳LOWLA���00����D��@�BwP��� �1RCʀ�ƶMOSIV�JRM�O���@GPERC7H  �OV�� ^��i�<!�ZD<!�c@��d@�P��V1�#P͑��L���EW�ĆĸUP������T�RKr�"AYLOA'a�� Q-�̒<�1�8�`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H�����b�DUM2(�S_�BCKLSH_C ̒��>�=�q�#�U��������2�t�]ACLA�LvŲ�1n�P�C�HK00'%SD�RT�Y4�k��y�1�q_�6#2�_UM$Pj�C�w�_�SCL��ƠLMT_J1_LO�"�@���q��E������๕�幘SPC`��7������PCo�B��H� �PU�m�C/@��"XT_�c�CN_b��N��e���SFu���V�&#����9�̒d��=�C�u�SH6# ��c����1�Ѩ�o�0�0͑
��_�PAt�h�_Ps�W�_10��4֠R�01D�VG�J� L��@J�OGW���ToORQU��ON*ɀMٙ�sRHљ��_	W��-�_=��C��TI��I�I�II�	F�`�JLA.�1[��VC��0�D�BO1�U�@i�B\JRK�U��	@DBL_�SMd�BM%`_D9LC�BGRV��0C��I��H_� �*COS+\�(LN�7+X>$C�9)�I�9)u*c,)�Z2 HƺMY@!�( "�TH&-�)THET=0�NK23I��"l=�A CB6CB=�C�A�B(261C�61�6SBC�T25GT	S QơC��aS$�" �4c#�7r#$DUD�EX�1s�t��B�6䆱�AQ|r�f$NE�DpIB U�\B5��	$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2��&�C�J�&!�VAHV�6H3�YLVhJVuKV��KV�KV�KV�KV�IHAHZF`RXM��wX�uKH�KH�KH�KH��KH�IO2LOAHOT�YWNOhJOuKO�KUO�KO�KO�KO�&�F�2#1ic%�d4GS�PBALANCE�_�!�cLEk0H_�%SP��T&�bc&�b>r&PFULC�hr��grr%Ċ1ky�U�TO_?�jT1T2Cy��2N&�v�ϰ ctw�g�p�0Ӓ~����T��O���� IN�SEGv�!�REV8�v!���DIF�鉳1l�w�1m�0OaB�q
����MIϰ�1��LCHWAR̭���AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|�n��ROBR�CR�����N�'�MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD�0�ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDX�Р  ��MOR^��t $-�U�� )��r�B���͓��Gؒu � $SIMULT ��~�x�� ���OBJE�`> �ADJUS>�1�OAY_Ik��D_�����C�_FIF�=�T� ��Ұ��{���p� �����p�@��DN�FRI��ӥT�ՓRO� ��E����͐OPWO�ŀv�0��SYSBU<�@ʐ$SOP�����#�U"��pPRUYN�I�PA�DH��D����_OU��=��qn�$}�IMKAG��ˀ�0P�q3IM����IN�q�~��RGOVRDȡ:���|�P~���Р�0�L_6p���i��R)B���0��M���SEDѐF� ��N`�M*������˱SL��`ŀw x $�OVSL�vSDI��DEXm�g�e�9Hw�����V� ~�N����w����Ûǖȳ�M��͐�q<��� �x HˁE�F�AWTUS���C�08àǒ��BTM����If���4����(�.ŀy DˀEz�g���PE�r�����
���EXE��V��E�pY�$Ժ ŀz @ˁf��UP{�h�$�p��XN���9�H�� �PG"�{ h $SUB���c�@_��01\�MP�WAI��P����L�O��-�F�p�$�RCVFAIL_9C�-�BWD"�F����DEFSPup | Lˀ`�D��8� U�UNI���S���R`���_L*�pP���P�ā}��� B�~���|��`:ҲN�`KET��y����P� $�~���0SIZE�ଠ�{���S<�OR��FORMAT/p � XF���rEMR���y�UX�����P�LI7�ā  �$�P_SWI������_PL~7�AL_ �ސJR�A��B�(0C���Df�$Eh��ւ�C_=�U� � � ���~��J3�0����TIA�4��5��6��MOM������ �B�AD��*��*6 PU70NRW���W ��V����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�!O�0\H��6@���U�� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�Hӱt@�W�UpS��ћ�L;@���O㵐.'}q��C�g���@ʣ���тM��AÂ� � $sPY��$WH`'�NGp���H`��Fb`��Fb��Fb��PLM�@��	� 0h�H�{�X��	O��z�Z�eT�M���G� pS��C���O__0_B_�a��_%�� |S����@	 �v��v �@���w�v2��EM��% �frJ�B�ː��ftP��PM��QU� ��U�Q��A-�Q�TH=�HOL��Q7HYS�ES�,��UE��B��O#��  -�P0�|�gAQ�(��ʠu���O��ŀ��ɂv�-�A;ӝR#OG��a2D�E��Âv�_�ĀZ�INF�O&��+����b�v��OI킍 (��SLEQ/�#� �����o���S`c0QO�0�01EZ0sNUe�_�AUT�Ab�COPY��Ѓ�{��@M��N�����1h�P�
� ��RGI������X_�Pl��$�����`�W��P���j@�G���EX_T_CYCtb����p����h�_N�A�!$�\�<�R�O�`]�� � 9m��POR�ㅣ\���SRVt�)��6��DI �T_l����Ѥ{�ۧ��ۧ �ۧ5*٩6٩7٩8��A��PS�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#q���Q�SKIP�� Ĵ��x�O�`NT!���P_x���ǚ@ �b�p1�1�1Ǹ� ?� �?��>��>�&��>�3�>�9�J2�R;쐖 4��EX� TQ����ށ�Q����[�KFд���R;DCIf� �U`�X}�R�#%M!*�0��)��$RGEAR_�0IO�TJBFLG��igpERa��TC�݃������2TH2�N��� 1� ��Gq T�0 �����M���`I�b���AREF�1��� l�h��ENsAB��lcTPE?@ ���!(ᭀ����Q �#�~�+2 H�W���2�Қ���"�4�F�X�j�3�қ{���P������j�4�Ҝ��@
��.�@�R�j�5���u�����������j�6�Ҟ��(:Lj�7�ҟo�������P��8�Ҡ���"4Fj�SwMSK��  ��+@��E�A����M�OTE�����`�@ "1��Q�IO�5�"%I��P���PO9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C�ШP^�S232%�Sb��iDEVICEU�S#�R�RPARI�T�!OPBIT��Q��OWCON�TR��Qⱓ�RC�U� M�SUXTA�SK�3NB��0�$TwATU�P�8��RS@@쐦F�6�_��PC}�$FRE?EFROMS]p�a�i�GETN@S�UPeDl�ARB��SP%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG �G|�.2���F��1�!d�9Z�8+5K��+5��E�y�L0�4��X �0m�LN�T�3Hz��89��%�4�3%G��W�0�W�RdD�Z��Tܳ��K�a�3d��$cV 2!���1��I1H�0U2K2sk3K3J ci�aI�i�a�L��SLL��R$Vؠ�BV�E�Vk��AbQ*R��� �,6Lc���9V2�F{/P:B��PS_�E���$rr�C�ѳ3$A0��wPR���v�U�cSk�� {�@#�2���� 0���VX`�!�tX`��0P��ꁂ
�5SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V����S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD��<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C���:c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQ�pfC��30=	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�q� �X��ȑ� �p.A$�1$�c1 Ē���7� x~�EG� ݓ��q!AR����0�9>B�%��AXE.��ROB��W�A4�_�-֣SY���!6���&S�'WR���-1���STR��5�:9�E�� 	5B��=QB90�@6�������OT�0o 	$�ARY8�w20�Ԛ�	%�FI��;�$LINK�H��1%�a_63�5�q�2XYZ"��;�qH�3@��1�2�8{0	B�{D��� CFI��6G��
�{�_J��6��3NaOP_O4Y;5�FQTBmA"�BC
�z�DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ �@�5<:7�� W1�?0K�Mc��68Cb�vrb�4�ORQ��X�>8�#op ������wq�Uf����N�TOVE�Q��M;����E#�UK#�UQ"�VW �ZQ�W���Tυ� ;� ����QH�!`�ҽ��U��Q�WkeK#kecXE)R��	GE	0��S�dAWaǢ:D���0�7!�!AX�rB !{q��1uy-! y�pz�@z�@z6P z\Pz� z1v� y�y�+y�;y� Ky�[y�ky�{y�x�y�q�yDEBU��$����L�!º2WG`  AB!�,�r�SV���� 
w� ��m���w����1���1 ���A���A��6Q��\Q����!�m@��2CLAB3B�U������S  V ER|���� � $@ڳ Aؑ!p�PO���Z�q0w�^�_M�RAȑ� d r T�-�ERR�L�TYz�B�I�qV3@�cΑTOQ�d:`L� �d2�p ��|˰[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	�SFZ�N_CFG_!� 4��?º�|�ų����8@�ȲW ]���\$� �n���Ѵ��09c�Q��(�FA�He�,�XEDM�(���H��!s�Q�g�P{R�V HELLĥ�� 56�B_BAS!�RSR��ԣo E�#S��[��1r�U%��2ݺ3ݺ4ݺU5ݺ6ݺ7ݺ8ݷ��ROOI䰝0�03NLK!�CAB� n��ACK��IN��T:�1�@�@ z�m�7_PU!�CO� ��OU��P� Ҧ) ���޶��TPFWD�_KARӑ��R�E~��P��(�Q�UE�����P
��C�STOPI_AL �����0&���㰑�0GSEMl�b�|�M��6d�TY|�SOK�}�DI�����(����_TM\�MANR�Q�ֿ0E+�|�$�KEYSWITCaH&	���HE
�OBEAT��cE� �LEҒ���U��F�O�����O_HOuM�O�REF�P�PRz��!&0��Cr+�OA�ECO��xB�rIOCM�D8׵��]���8�` G� D�1����U���&�MH�»P�CFO3RC��� ����OM�  � @�V��|�U,3P� 1(-�`� 3-�4���NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F��V ��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7s|'��VP��UPD�� � ��|�԰
��Y�SLOǢ� � z��и���o�E��`p>�^t��АALUץL����CU���wFOq�ID_L�ӿuHI��zI�$FILE1_���t��$`�^�vMsSA��� h��~�E_BLCK��#�C,�D_CPU <�{�<�o����t����R ��
�PW O� ��L�A��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ� �T�BCu�C� ��X -$�LEN@i��v������I���G�LOW_AXI��F1��t2X�M�����D�
 ��I�� 9��}�TOR��"��Dh��� L=�������s���#�_MA�`�ޕ��ޑTCV����T���&��@ݡ����J�����J����Mo���J�Ǜ ��)�����2��� �v�����F�JK��V�Ki�Ρv�Ρ3��J�0�ңJJڣJJ�AALң�ڣ���4�5z�&�N1�-�9���␅�L~�_�Vj�*q���� =` �GROU�pD���B�NFLIC���REQUIREa�EBUA��p����2¯������c�� \��A�PPR��C���
v�EN�CLOe��S_M v�,ɣ�y
���� ����MC�&���g�_M	G�q�C� �{�9����|�BRKz�NO�L��|ĉ R��_L!I|��Ǫ�k�J����P
���ڣ�����&����/���6��6��8���������# ��8�%�W�2�e�PATHa�z�pӠz�=�vӥ�ϰ�x�CN=�CA�����p�IN�UC��bq��-CO�UM��YZ������qE%���2����~��PAYLOA���J2L3pR_AN��<�L��F�B�6�R��{�R_F2LSHR��|�LOG��р���ӎ���ACRL_@u�������.���H�p��$H{���FL�EX
��J�� :�/�����6�2�����;�M�_�F16����n���������ȟ��Eҟ���� �,�>�P�b���d� {������������5���T��X��v��� EťmFѯ��� ����&�/�A�S��e�D�Jx�� � �������j�4pATر���n�EL  ԁ%øJ���ʰJEΧ�CTR�Ѭ�TN���F&��HAND_VB[
�pK�7� $F2{�6Ì �rSW$#�U��?� $$Mt�h�R��08��@<b 35��^6A�p3�k��q{9t�QA�̈p��A��A��P�0��U���D��D��eP��G��IST��h$A��$AN��DYˀ �{�g4�5D���v�6� v��5缧�^�@��P�����#�,�5�t>�r�J�� &0��_�ER!V9�SQAS�YM��] �����px��ݑ���_SHl� ������sT�(����(�:�JA���S�ci\r��_VI�#Oh|9�``V_UNI��td�~�J���b�E�b ��d��d�f��n��� ������uN����vr��H�������"CqEN� a�DI���>�Obt2Dpx�S� ��2IxQA�� ��q��-��s �� �ܒ��� ��OMME��rr�QTVpPT�P ���qe�i����P�x ��y�T�Pj� $D�UMMY9�$7PS_��RFq�0;$:� ����!~q� X����K��STs�ʰSBR���M21_Vt�8�$SV_ERt�O���z���CLRx�A�  O�r?p? Oր �� D $GgLOB���#LO�ЀՅ$�o��P�!S;YSADR�!?p��pTCHM0 �� ,����W_N�A��/�e�$%S�R��l  (:]8:m�K6�^2m� i7m�w9m��9���ǳ� �ǳ���ŕߝ�9ŕ� ��i�L���m��_��_�_�TD�XSCR�E�ƀ�� ��STF���}�pТ6��1] _v AŁ�s T����TYP�r��K��u�!u��Z�O�@IS�!��uD�UE{t� �Ȯ��H�S���!RS�M_�XuUNEX�CEPWv��CpS_ ��{ᦵ�ӕ���÷�ӎ�COU ��� �1�O�UET����r���PROGM�� FLn!$CUƕ�PO*q��c�I_��pH;� � 8\��N�_HE
p���Q��pRY ?����,�J�*��;�O�US�� � @�d���$BUTT��R@���COLU�M�íu�SERV<c#=�PANEv Ł�� � �PGE�U�!�F��9�)$�HELP��WRETER��)״���Q ������@� P��P �IN��s��PNߠw v�1������ ���L�N�� ����_���k�$H��M T�EX�#����FLA�n +RELV��DP4p�������M��?,��ӛ$����P�=�USRVIE�WŁ� <d��pU:�p0NFIn i��FOCU��i�PR�ILPm+�q��T�RIP)�m�U9Njp{t� QP��XuWARNWud�S�RTOLS�ݕ�t����O|SORN��'RAUư��T��%���VI|�zu�� $�PATH�g��CACHLsOG6�O�LIMyb�M���'��"�HOS�T6�!�r1�R��OBOT5���I%Ml� D�C� g!���E�L���i�VCPU_AVAILB�VO�EX7�!BQNL��(���A�� Q��Qq ��ƀ�  Qp�C���@$TO�OL6�$�_JM�P� �I�u�$SS�!&; SHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3��(���w�2u��Pr{t��%�DJU��~|#�WAIT�������%ONE���YBOư ?�� $@p%�vC�SBn)TPE��NEC��x"�$t$��.�*B_T��R��% �qR� ���sB�%�tM�+��t�.�F�R!�݀��OPm�MAS��_DOG�OaT	�D����C3S�	�O2DELAY���e2JO��n8E��Ss4'#�J�aP6%�����Y_��O2� �2���5���`? kPZ�ABCS��  �$�2��J�
����$$CLAS��O���A����{ @VIRT��O.@ABS�$�1� <E� < *A tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R��d�v�����M@[�AX�Lր�&A�dC  ����IN��ā��P#RE������LARMRECO�V <I䂥�N�G�� \K	 �=#�
J�\�M@PoPLIC�?<E��E�Ha�ndlingTo�ol �� 
V�7.50P/28� *A�(m���
�_SW�� U�P*A� ��F0�ڑ����A)@��O 20��*A���y:����x(B� 7DA5 '@)�m@����Non�e������ ���T��*A4olx��P_���V����g�UT�OB�ค����HGAPON8@��LA�ѽU��D 1<EfA����������� Q 1שI Ԁ��Ԑ�:��i�n����#B�)B ���\��HE�Z�r�HTTHKY��$BI�[�m� ����	�c�-�?�Q� o�uχϙϫϽ����� ���_�)�;�M�k�q� �ߕߧ߹�������� [�%�7�I�g�m��� �����������W�!� 3�E�c�i�{������� ��������S/A _ew����� ��O+=[a s������� K//'/9/W/]/o/�/ �/�/�/�/�/�/G?? #?5?S?Y?k?}?�?�? �?�?�?�?COOO1O OOUOgOyO�O�O�O�O �O�O?_	__-_K_Q_���(�TO4�s���DO_CLEAN��|&��SNM  9� �9oKo]ooo��o�DSPDRY�R�_%�HI��m@ &o�o�o#5GY k}����"����p�Ն �ǣ�qX�Մ��ߢ��g�PLU�GGҠ�Wߣ��PRUC�`B`9��o��=�OB��o&�SEGF��K������o %o����#�5�m���LAP�oݎ������ ����џ�����+��=�O�a���TOTA�L�.���USENUʀ׫ �X���R�(�RG_STRI�NG 1��
��M��Sc��
��_ITEM1 �  nc��.�@� R�d�v���������п �����*�<�N�`��r�I/O S�IGNAL���Tryout M�ode�Inp���Simulat{ed�Out��OVERR�`� = 100�In cycl����Prog A�bor�����S�tatus�	H�eartbeat���MH FauylB�K�AlerU� ��s߅ߗߩ߻�����8���� �S�� �Q��f�x���� ����������,�>��P�b�t�������,�WOR������V��
 .@Rdv�� �����*8<N`PO��6� ���o����� //'/9/K/]/o/�/ �/�/�/�/�/�/�/�DEV�*0�?Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO��O�O�OPALT B��A���O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:o�OGRI�p��ra�OLo �o�o�o�o�o�o *<N`r��� ���`o��RB�� �o�>�P�b�t����� ����Ώ�����(��:�L�^�p����PREG�N��.������ ��*�<�N�`�r��� ������̯ޯ����&����$ARG_���D ?	����i�� � 	$��	+[}�]}���Ǟ��\�SBN_CON?FIG i��������CII_SAVE  ���۱Ҳ\�TCEL�LSETUP �i�%HOME�_IO�͈�%M�OV_�2�8�RE�P���V�UTOB�ACK
�ƽFRA:\��� �Ϩ���'`�!��������� ����$�6�c�Z�8lߙ��Ĉ������ �������!凞��M� _�q����2����� ����%�7���[�m� �������@�������`!3E$���J�o�������I�NI�@��ε~��MESSAG�����q��ODE_!D$���O,0.ޜ�PAUS�!�~i� ((Ol� ������� / �//$/Z/H/~/l/�/�'akTSK � q�����UP3DT%�d0;�WSM_CF°�i�еU�'1GRgP 2h�93 |��B��A�/S�XSC�RD+11
1; 	����/�?�?�?  OO$O��߳?lO~O �O�O�O�O1O�OUO_  _2_D_V_h_�O	_X�>��GROUN0O��SUP_NAL��h�	�ĠV_ED�� 11;
 �%�-BCKEDT�-�_`�!oEo%����a��o����,�ߨ���e2no_��o�o�b���ee�o"�o�oED3�o��o ~[�5GED4�n#�� ~�j���ED5Z��Ǐ�6� ~���}���ED6����k�ڏ ~G���!�3�ED7��Z���~� ~�V�şןEDa8F�&o��Ů}p����i�{�ED9���W�Ư
}3�����CRo�����3��տ@ϯ����P�PNO�_DEL�_�RGE?_UNUSE�_�T�LAL_OUT �q�c�QWD_ABOR� �΢Q��ITR_RTN�=���NONSe����CAM_PARAM 1�U�3
 8
SO�NY XC-56� 2345678�90�H � �@���?���(O АV�|[r�u�~�X�HR5k�p|U�Q�߿�R57�����Aff��K�OWA SC31�0M|[r�̀�d @6�|V�� _�Xϸ���V��� ����$�6��Z�l��CE�_RIA_I8j57�F�1��tR|]��_LIO4YW=� ��P<~��F<�GP 1�,���_GYk�*C*  ��CU1� 9� @� G� Z�CLC]� d� l� s�R� ��U[�m� v� � }�� �� C�� ő"�|W��7�HEӰONFI� ��<�G_PRI 1�+P�m®/���������'CHK�PAUS�  1E� ,�>/P/:/ t/^/�/�/�/�/�/�/ �/?(??L?6?\?�?"O�����H�1�_MOR�� }��PBZ?����5 	 �9 O�?�$OOHOZK�2	��H�=9"�Q?55��CR�PK�D3P����>��a�-4�O__|Z
�OG_�7�P O�� ��6_��,xV�A�DB���='�)
�mc:cpmidcbg�_`��S:�)�	���Yp�_)o�S`�BBi�P�_mo8j�)�Koo�oV9i�)��og�o�o�m�of�oGq:�I�ZDEF �f8��)�R6pbuf.txtm�]nd�@����# 	`)н��A=L���zM-C�21�=��9����4�=�n׾�C�z  BHBCCP�UeB��C�F�;.<C�?��C5rSZE@�D�nyDQ���D��>���D�;D�����F��>F��$G}RB�oGzր��SYR��!�vqG���E�m�)�.��)�b)��<�q�G�x2ʄ�Ң �� a�D��j���E�e��EX��EQ�EJP� F�E�F�� G�ǎ^F� E�� FB�� H,- Ge�߀H3Y��� � >�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE d�O c
�(�;�"�G  <�6�z�R���?�j�C4��SZm� W��{�m��C��B-G�C�`@�$�q��T{�FP?ROG %i����c�I��� �Ɯ�f��KEY_TBL � �vM�u� �	
��� !"�#$%&'()*+,-./01c��:;<=>?@A�BC�pGHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������p����͓���������������������������������耇���������������������!j�LCK��.�j����STAT���_AUTO_DO����W/�INDT_'ENB߿2R��9��+�T2w�XSTO�P\߿2TRLl�L�ETE����_S�CREEN ~ikcsc���U��MMENU �1 i  <g\��L�SU+�U�� p3g���������� ��2�	��A�z�Q�c� ��������������. d;M�q� �����N %7]�m�� �/��/J/!/3/ �/W/i/�/�/�/�/�/ �/�/4???j?A?S? y?�?�?�?�?�?�?O �?O-OfO=OOO�OsO �O�O�O�O�O_�O_�P_Sy�_MANU�AL��n�DBCO�U�RIG���DB'NUM�p��<����
�QPXWORK 1!R�ү�_o�O.o@oRk�Q_AW�AY�S��GCP� ��=��df_AL�P�db�RY��������X_�p 1"�� , 
�^���o( xvf`MT�I^�rl�@�:sONTIM6������Zv�i�
õ�cMOTNE�ND���dRECO_RD 1(R�a��ua�O��q�� sb�.�@�R��xZ��� ����ɏۏ폄��� #���G���k�}����� <�ş4��X���1� C���g�֟�������� ӯ�T�	�x�-���Q� c�u����������>� ���)Ϙ�Mϼ�F� ࿕ϧϹ���:����� ��%�s`Pn&�]�o��� ��~ߌ���8�J���� ��5� ��k����ߡ� ��J�����X��|�� C�U�����������0�����	��dbTO�LERENCqdB�Ⱥb`L�͐PC�S_CFG )��k)wdMC:�\O L%04d.'CSV
�pc�)s[A �CH� z�p�)~���hMR�C_OUT *��[�`+P SGN� +�e�r��#��10-MAY-�20 09:27~*V27-JANj�21:48�k P;���)~��`pa�m�?�PJPѬ�VERSION �SV2.�0.�6tEFLO�GIC 1,�[ 	DX�P7)�P�F."PROG_E�NB�o�rj ULS�ew �T�"_WRSTJNEp�V�r`d�EMO_OPT_�SL ?	�es
� 	R575 )s7)�/??*?<?'>�$TO  �-�l�?&V_@pEX�W�d�u�3PATHw ASA\�?��?O/{ICT�aF�o`-�gds�egM%&AST?BF_TTS�x�Y�^C��SqqF�PM�AU� t/XrMSWR.�i6.|S/�Z!D_N�O0__�T_C_x_g_�_�tSB�L_FAUL"0��[3wTDIAU 1�6M6p�A�12345678#90gFP?Bo Tofoxo�o�o�o�o�o �o�o,>Pb��S�pP�_ �� �_s�� 0`��� ��)�;�M�_�q��� ������ˏݏ��|)gUMP�!� �^��TR�B�#+�=�P�MEfEI�Y_TE{MP9 È�3@8�3A v�UNI�.(�YN_BRK �2Y)EMGDI�_STA�%WЕN�C2_SCR 3��1o"�4�F�X� fv���������#��ޑ14����)��;�����ݤ5�����x�f	u�ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/߭P�b�t��  ��xߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N���r������� ��������&8 J\n����� ���"`�FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/4 ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O?�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�O�O�o�o�o 
.@Rdv� �������� *�<�N�`�r����o�� ��̏ޏ����&�8� J�\�n���������ȟ�ڟ����H�ETM�ODE 16��]� ��ƨ�
R�d�v�נRRO�R_PROG �%A�%�:߽�  ���TABLE  A������#�L��RRSEV_NU�M  ��Q���K�S���_AU�TO_ENB  q��I�Ϥ_NOh�� 7A�{�R��  *������������^�+��Ŀֿ迄�HISO���I��}�_ALM 18.A� �;�����+�e�wωϛϭ����_H���  �A���|��4�TC�P_VER !�A�!����$EXTLOG_REQ�s�{�V�SIZ_�~Q�TOL  ���Dz��=#�~��XT_BWD��p��r���n�_DI��7 9��}�z�x��m���STEP�����4��OP_DO����ѠFACTORY_TUN��dG�EATURE� :����l��HandlingTool ���  - CE�nglish D�ictionar�y��ORDE�AA Vis�� ?Master����96 H��nal?og I/O����H551��uto� Softwar�e Update�  ��J��mat�ic Backu�p��Part�&�ground �Edit��  8�\apCam�era��F��t\;j6R�ell����LOADR�omm���shq��TI"� ��co��
!� o���pane��� 
!��t�yle sele�ct��H59��n�D���onitorf��48����tr��?Reliab����adinDiagnos"�����2�2 ual Ch�eck Safe�ty UIF l�g\a��hanc�ed Rob S�erv q ct�\��lUser sFrU��DIF���Ext. DIOm ��fiA d���endr Err� L@��IF�rd��  �П�90���FCTN MeneuZ v'��74� �TP In��fa�c  SU (�G=�p��k Excn g�3���High-Spe�r Ski+�  s�O�H9 � mmun�ic!�onsg�tFeur� ����V�����conn���2��EN��In{crstru�����5.fdK�AREL Cmd7. L?uaA� �O�Run-TiN� Env����K� ���+%�s#�S/W���74��Lice�nseT�  (�Au* ogBoook(Sy��m)���"
MAC�ROs,V/Of�fse��ap��MqH� ����pfa5��MechStop� Prot��� �d�b i�Shiyf���j545�!�xr ��#��,+{�b ode Sw�itch��m\eҙ!o4.�& p#ro�4��g��Multi-T7�G��net.�Pos Regi���z�P��t Fsun���3 Rz1��Numx ������9m�1�  Adjyuj��1 J7�7�* ����6tat�uq1EIKR�DMtot��scove�� ��@Bxy- }uest1��$Go� � U5\?SNPX b"��x�YA�"Libr�����#�� �$~@h��pd]0�Jts in VCCM�����0�  �u!��23 R�0�/I�0�8��TMILIB^�M J92�@P�gAcc>�F�97��TPTX�+�BRS�QelZ0�M8 Rpm��q%��692���Unexcept�r motnT  �CVV�P���KC�����+-��~K  �II)�VSP C7SXC�&.c�� e��"�� t�@W9ew�AD Q�8bsvr nmen�@��iP� a0y�0��pfGridAplay !� nh�@�*�3R�1M-10iA(B201 �`�2V"  F���sc{ii�load��/83 M��l�����Guar�d J8	5�0�mP'�L`���;stuaPat�&]$�Cyc���|0oryi_ x%Data'P3qu���ch�1�h�g`� j� RLJ�am�5���IMI� De-B(\A�cP�" #^0C  �etkc^0assswo%q�)650�A1pU�Xnt��P�ven�CTqH�5��0YELLO�W BO?Y��� A;rc�0vis��Ch�WeldQc�ial4Izt�Oap� ��gs�` 2@�ma��poG yR�jT1 NE�#HT�� xyWb��! �p�`gd`���p\�� =P��JPN A7RCP*PR�A��� OL�pSup̂fil�p��J��� ��cro�670`�1C~E�d��SS�p]e�tex�$ �P�� So7 t� ssKagN5 <Q�BP:d� �9 "0�QrtQ�C��P�l0dpn��笔�rpf�q�e�pp�mascbi�n4psyn�' �ptx]08�HEL�NCL VIS? PKGS �Z@�MB &��B J�8@IPE GE�T_VAR FI�?S (Uni� L�U�OOL: AD}D�@29.FD�TiCm���E�@DVp���`A�ТNO WTWTEST ��� 6�!��c�FOR� ��ECT �a!�� ALSE AL�A`�CPMO-1�30��� b D: �HANG FRO�Mg��2��R70�9 DRAM A�VAILCHEC?KS 549��m�VPCS SU֐�LIMCHK��P��0x�FF POS� F�� q8�-12 CHAR�S�ER6�OGRA� ��Z@AVEH�A;ME��.SV��В�אn$��9�m "�y�TRCv� SH�ADP�UPDAT� k�0��STAT�I��� MUCH� ���TIMQ �MOTN-003���@OBOGU�IDE DAUG�H���b��@$to�u� �@C� �0��P�ATH�_�MOV{ET�� R64���VMXPACK �MAY ASSE�RTjS��CYCL�`�TA��BE C�OR 71�1-�A�N��RC OPT?IONS  �`���APSH-1�`fix��2�SO��B�0�XO򝡞�_T��	��i��0j��du�byz p wa��y�٠#HI������U�pb XSPD TB/��F� \hchΤBl0���END�CE�0�6\Q�p{ smOay n@�pk���L ��traff�#�	� ��~1fr�om sysva_r scr�0R� ���d�DJU���H��!A��/��SET� ERR�D�P7�����NDANT �SCREEN U�NREA VM 4�PD�D��PA����R�IO JNN��0�FI��B��G�ROUNנD Y��Т٠�h�SVI�P 53 QS��D�IGIT VERqS��ká�NEW�� P06�@C�1I�MAG�ͱ���8�� DI`���pSS�UE�5��EPLA�N JON� DE�L���157QאD��CALLI���Qx��m���IPND}��IMG N9 P�Z�19��MNT/Υ�ES ���`LocR Hol߀=��2:�Pn� PG:��=�M��can����~С: 3D mE2�view d XL��ea1 �0b�pwof Ǡ"HCɰ��ANNOT A�CCESS M �cpie$Et.Qs� a� loMdFl�ex)a:��w$qmWo G�sA9�-'p�~0��h0pa��eJ? AUTO-�0���!ipu@Т<ᡠI/ABLE+� 7�a ?FPLN: L�gpl m� MD<��VI�и�WIT �HOC�Jo~1Q�ui��"��N��U�SB�@�Pt & remov���D�v�Axis FT_t7�PGɰCP:�OS-144 � ?h s 268QՐ�OST�p  CR�ASH DU��$�P��WORD.$>�LOGIN�P���P:	�0�046 issueE�H�: Slow +st�c�`6����໰IF�IMPR���SPOT:Wh84���N1STY��0�VMGR�b�N�CkAT��4oRRE��9 � 58�1���:%�RTU!Pe -\M a�SE:�@pp�H��AGpL��m�@all��*0a�O�CB WA���"3 CNT0 T9D�WroO0alarqm�ˀm0d t�0M�"0�2|� o�Z@�OME<�� ��E% w #1-�SRE���M�st}0g   �  5KANJ�I5no MNS�@�INISIToALIZ'� E��f�we��6@� dr��@ fp "��S�CII L�afa�ils w��SYSTE[�i���  � Mq�1QG;ro8�m n�@vA����&��n�0q���RWRI OF �Lk��� \ref�"�
�up� de-�rela�Qd 0k3.�0SSchő�betwe4�IN�D ex ɰTPFa�DO� l� ��ɰGigE�sop�erabil`p l,��HcB��@]��le�Q0cflxpz�Ð���OS {�����v4pfigi GCLA�$�c2�7H�� lap�0ASBֻ If��g�2 lC\c�0�/�E��? EXCE 㰁�!P���i�� o0��Gd`]Ц�fq�l �lxt��EFal���#0�i�O�Y�n�CwLOS��SRNq1+NT^�F�U��Fq�KP�ANIO V7�/ॠ1�{����D�B �0��ᴥ�EDN��DET|�'� �}bF�NLINEb�GBUG�T���C"R�LIB��A��ABC JARKY@���� rkey�`I)L���PR��N��ITWGAR� D$�R  �Er *�T��a��U�0��h�[�ZE �V� TASK op.vr�P2" 8.�XfJ�srn�S谎�dIBP	c���B�/��BUS��UNN� j0-�{��c�R'���LOE�DIVS�CULs$cb����BW!��R~�0W`P�����IT(঱�tʠ�OF��UN#EXڠ+���p�Ft}E��SVEMG3`NML 505� �D*�CC_SAF�E�P*� �ꐺ� P�ET��'P�`�F  !���IR����c� i S>� K��K��H GUNCH�G��S�MECH���M��T*�%p6�u��tPORY L�EAK�J���S�PEgD��2V 74\GRI��Q�gޙ�CTLN��TR�e @�_�p ���EN'�IN������$��̸r��T3)�i�ST%O�A�s�L��͐!X	���q��Y� ���TO2�J m��0F0<�K����DU�S��%O��3 9�J �F�&���SSVG�N-1#I���RS	RwQDAU�Cޱ� �T�6�g��� 3�]���BRKCTR/"� �q\j5��_�Q�S�q�INVJ0D ZO �Pݲ���s��г�Ui �ɰ̒�a�DUAL�� J50e�x�RVO117 AW��TH!Hr%�N�24�7%�52��|�&aol ���R���at�S�d�cU���P,�LE�R��iԗQ0�ؖ  CST���Md�Rǰ�t� \fosB�A��0Np�c����{�U>��ROP 2�b�p}B��ITP4M��b !AUt c0< >� plete�N@�� z1^qR63�5 (AccuC�al2kA���I)C "�ǰ�1a\�Ps��ǐ� bЧ0P��������ig\cbacul "A3p�_ �1��ն���et�aca��AT���PaC�`�����_p��.pc!Ɗ��:�c�ircB���5�tl0��Bɵ�:�fm+��Ċ�V�b�ɦ�r�upfrm.����ⴊ��xed��Ί�~�pe�dA�D �}b�pt�libB�� �_�r!t��	Ċ�_\׊���6�fm�݊�oޢ� e��̆Ϙ���c�Ӳ�b5�j>�����tcȐD��	�r����mm 1��T�sl^0��T�1mѡ�#�rm3��qub Y�q�std}�f�pl;�&�ckv�=�r�vf�䊰��9�cvi����ul�`h�0fp�q �.f���� daq; i D�ata AcquWisi��n�
�h�T`��1�89����22 DMCM� RRS2Z�75���9 3 R71Y0�o59p5\�?��T "��1 #(D�T� nk@�� ������E Ƒȵ��Ӹ��etdmm ��ER����gE��1�q\mo?۳�= (G���[(

�2��` ! �@JMA�CRO��Skip?/Offse:�a���V�4o9� &qR�662���s�H�
 6Bq8�����9Z�43 J77z� 6�J783��o ��n�"v�R5�IKCBq2 PgTLC�Zg R�w3 (�s, �0������03�	з�JԷ\sfmnmc "MNMC�����ҹ�%mnf�F�MC"Ѻ0ª et�mcr� �8����� ,+{�D6{   �874\prdq�>,jF0���ax�isHProce�ss Axes �e�rol^PRA�
�Dp� 56 J8m1j�59� 56oa6� ���0w�690 s98� [!IDV�1Ĵ�2(x2��2ont�0�
����m2���?C��etis "ISD��9��^ FpraxRAM�Pp� D��defB��,�G�isbasicHB�@޲{6��� 708�6��(�Acw:������D
��/,��AMOX�� ��D@vE��?;T��>Pi� �RAFM';�]�!PAM �V�W�Ee�U�Q'
�bU�75�.�ce�Ne� nterfGace^�1' 5&!�54�K��b(Devam±�/�#���/<��Tane`"DNE�WE���btpdnu�i �AI�_s2�d_rsono���b�AsfjN��bdv_arFvf�xhpz�}w抰hkH9xstc8��gAponlGzv{�ff��r����z�3{q'Td>p�champr;e�p� ^5977��	܀�4}0��mɁ�/������lf�!�pcchmp]aMP&B�� �mpev������pcs��YeS�� _Macro�OD��16Q!)*�:$�2U"�_,��Y�(PC  ��$_;������o��J��gegemQ@GE�MSW�~ZG�ges�ndy��OD�ndd1a��S��syT�KɆ��su^Ҋ���n�mx���L��  ����9:p'ѳ޲��sp?otplusp����`-�W�l�J�s��t8[�׷p�key�ɰ��$��s�-Ѩ�m���\�featu 0FEqAWD�oolo�srn'!2 p����a�As3��tT.� (N. A.)�@�!e!�J# (j��,��oBIB�oD �-�.�n��k9�"AK��u[-�_���p� "PSEqW��~��wop "sE� ��&�:�J������y� |��O8��5��Rɺ�� ��ɰ[��X������ �%�(
ҭ�q HL�0k�
�z�a!�B�Q�"(g�Q��� ��]�'�.�����&���`<�!ҝ_�#��tpJ� H�~Z��j�����y�� ����2��e������Z ����V��!%���=��]�͂��^2�@iRV�� on�QYq͋J�F0� 8ހ�`�	(|^�dQueue����X\1�ʖ`�+F1tp/vtsn��N&��f�tpJ0v �RDV �	f��J1 Q����v�en��kvs�tk��mp��btkclrq���get����r<��`kack�XZ��strŬ�%�satl��~Z�np:! �`���q/�ڡ6!!l�/Yr�mc�N+v3�_� �����.v�/\jF��� �`Q�΋ܒ�N5?0 (FRA��+���͢frapar�m��Ҁ�} 6�J�643p:V�ELS�E
#�VAR �$SGSYSCF�G.$�`_UNITS 2�DG~°@��4Jgfr��4A�@FRL-��0ͅ�3ې�� �L�0NE�:�=�?@@�8�v�9~Qx304�8�;�BPRSM~Q�A�5TX.$VNUM_OL��5��D�J507��l� Functʂ"qwAP8��琉�3 H�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6N�k�AP����S��"T�PPR���QA�prnaSV�ZS��AS^8Dj510U�-�`�cr�`8 ��ʇ�DJ�R`jYȑH  k�Q �PJ6�a�21��48A�AVM 5�Q�b0y lB�`TUP xbJ545 `b��`616���0�VCAM 9��CLIO b1��5 ���`MSC�8�
rP R`\s�STYL MN{IN�`J628Q;  �`NREd�;@��`SCH ��9pD�CSU Mete>�`ORSR Ԃ�a�04 kREI�OC �a5�`542�b9vpP<�nP�a��`�R�`7�`�MASK Ho��.r7 �2�`OCO	 :��r3��p�b�p����r0X��a�`13�\mn�a39 H�RM"�q�q���LCHK�uOPLsG B��a03 �q=.�pHCR Ob�p=CpPosi�`fP�6 is[rJ5594�òpDSW�bM�qD�pqR�a37 }Rfjr0 �1�s4 �R�6�7��52�r5 \�2�r7 1� P6�~��Regi�@�T�uFRDM�uStaq%�4�`930�u�SNBA�uSHL]B̀\sf"pM��NPI�SPVC��J520��TC��`"MNрTMI�L�IFV�PACy W�pTPTXp�6.%�TELN oN Me�09m3?UECK�b�`�UFR�`��VCO�R��VIPLpq8�9qSXC�S�`VV9F�J�TP �q���R626l�u S��`Gސ�2IGsUI�C��PGSt�=\ŀH863�S�qX�����q34sŁ684���a�@b>�33 :B��1 T���96 .�+E�51� y�q53�3�b1� ���b1 n�jr9y ���`VAT ߲�q75 s�F��`�s�AWSM��`TO3P u�ŀR52p����a80 
�ށXY� q���0 ,b�`8k85�QXрOLp�}�"pE࠱tp�`L�CMD��ETSS����6 �V�CP�E oZ1�VRC�d3
�NLH�h��0c01m2Ep��3 f���p��4 /165�C��6l���7PR���008 tB��9� -200�`U02�pF�1޲1 ��޲A2L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�~J�7 rbcfA��L�8\PC����"�3!2m0u�n�K�Rٰn�5 5EW
n�s9 z��40 kB���3 ��6ݲ�`0/0iB/��6�u��	7�u��8 µ�������sU0�`�t �1 �05\rb��2 �E���K���j���5˰��60��a�HУ`:�63�jAF�_���F�#7 ڱ݀H�8�eH�L���cU0��7�p���1u��8u��9� 73������D7�� ��5t�97 ���8U�1��2��1R�1:���h��1np��"��8(�U1��\pyl��,࿱v ��.B�854��1V���ZD�4��im��1� <���>br�3pr�q4@pGPr�6 B��H�цp��1����1�`�͵155ض157 �2��62�S�����1b��2����1dΠ"�2���B6`2�1<c�4 7B��5 DR��8_�B/���187 uJ�8w 06�90 rB�n�1 (��202_ 0EW,ѱ2^�4�2��90�U2�p�2���2 b��4��2N�a"RB����9\��U2�`w�l���4 60Mp��7������Xb�s
5 ��3��x��pB"9 3 ��؆�`ڰR,:7  �2��V�2��5���2�^��a^9���qr����n�5����5�D��"�8a�Ɂ}�5B�"��5����`UA���d� ��86 �6 S��0��5�p�2�#�529 �2^�b1P�5~�2`���T&P5��8��5���u�!�5��ٵ544J��5��R�ąP nBX^z�c (�4�������U5J�V�5��1�1^��%����:��5 b21��lgA��58W82� �rb��5N�E�58�90r� 1�95 �"������c8"a�@�|�L ���!J"5|6��^!�6��B�"�8�`#��+�8%�6�B�AME�"1 i�C��622�Bu�6hV��d� 4��84�`�ANRSP�e/S� C�5� �6� ��� \� �6� �V� �3t��� T20CA�R��8� Hf� �1DH�� AOE� ��� ,+|��� �0\�� �!64�K��ԓrA� �1 (�M-7�!/50T@�[PM��P�Th:1 �C�#Pe� �3�0� }5`M75T"� �D8p� �0Gc� u��4��i1-710i��1� Skd�7j�?6�:-HS,� �RN��@�UB�f�X�=m�75sA*A6an����!/CB�B2.6A  �0;A�CIB�A�2�QF1ԣUB2�21� /7!0�S� �4����Aj1�3p���r#0 B'2\m*A@C��;bi"i1K�u"A~AAU� ?imm7c7��ZA�@I�@�Df�A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A�EA��5B�4>\77
B7@=Q�D�2�Q$B�E7�CJ�D/qAHEE�W7�_ |`jz@� 2�0�EBjc7�`�E"l7�@�7�A
1�E�V~`�W2�%Q�R9ї@0L_�#����"A���b��9H3s=rA/2�R5 nR4�74rNUQ1ZU�A�s\m9
1M92�L2�!F!^Y�ps� 2cci��-?�qhimQ �t  w043�C�p2�mQ0�r�H_ �H20�Evr0�QHsXBSt62�q`s������ ��Pxq3g50_*A3I)�2��d�u0�@� '4TX��0�pa3i1A3`sQ25�c��st�r"�VR1%e�q0
�� j1��O2 �A�UEi�y�.�‐ �0Ch20$CXB79#A�ᓄM 8Q1]�~�� 9�Q�� ?PQ��qA!Pvs� 5 	15aU���?PŅ�8��ဝQ9A6�zS*�7�qb5�1����QN��00P(��V7]u �aitE1���ïp?7�� !?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ���y00\ry�"�R2BL�tN  ���� �1D�6{�2�qeR�5����_b�3�X]1m1lcqP1�a�E�Q� �5F����!5���@M-16Q�� f���r� �Q�e� ��� PN�LT_�1��i1��94�53��@�e�|�b1l>F1u*AY2�
��R8�Q����RJ�cJ3�D}T� 85
Q g�/0��*A!P�*A��Ȑ𫿽�2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt ]1^u�ajrI�B�����~�|I�b��yI�\m�Qb�I�uz�A�c3A�pa9q� B6S��S0��m���}�85`N�>N�  �(M ���f1���6����16�1��5�s`�SC��U��A����5\s�et06c����10�y�h8��a6���6��9r�2HS @���Er���W@}�a�� I�lB���Y�ٖ�m�u�C����5�B��B��h`�F���X0��@�A:���C�M��AZ��@��4�6i����� e�O�-	���f1�� �F �ᱦ�1F�Y	���T6HL3��U66�~`���U�dU�9D20Lf0��Qv� ��f jq��N������0v
�� ��i	�	��72lqQ2������� �\chngmove.V��d���@2l_arf	�f ~��6������9C��Z���~���kr4�1 S���0��V��t������U�p7n�uqQ%�A]��V�1E\�Qn�BJ�2 W�EM!5���)�#�:�64��F�e50S�\��0�=�PV ���e������E��x���m7shqQSH"U��)��9�!A��(����� ,+{�ॲTcR1!��,�60e"=�4F�����2��	 R-��������Ӏ��Ж��4���LS`R�)"�!lOA��Q�) %!� 16�
 U/��2�"2�E�9p��|�2X� SA/i��'�
7F�H�@!B�0 ��D���5V��@2c@VE����T��pt���1L~E�#�F�Q��9E�#De/��RT��59���	�A�EiR��������9\m20�20��+�-u�19r4�`�E1�=`O9`@�1"ae��O�2���_$W}am41�4��3�/d1c_stAd��1)�!�`_T���r�_ 4\jdg �a�q�PJ%!~`-�r��+bgB��#c30�0�Y�5j�QpQb1��bq��vB��v25��U�����qm43 � �Q<W�"PsA�� e����t�i�P �W.��c�FX.�he�kE14�44��~6\j4�44�3sj��r�j4up@���\E19�h�PA�T �=:o�APf��coW�o!\�2a��2A;_2��QW2�bF�(�V11�23�`��X,5�Ra21�J*9$�a:88J9X�l5�m1a첚��*���(85�&������ �P6���R,52&AĀ���,fA9IfI50	\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP1���vB)e�m�����1pw� �1D6{�2�7�F�KAREL� Use S��F�CTN��� J9a7�FA+�� (�Q`޵�p%�)?�Vj9F?�(�j�Rtk208� "Km�6Q�y�j��iæPr�9�s#���v�krcfp�RC�Ft3���Q��kcc7tme�!ME�g�����6�main�dV�� ��ru��kD��c���o����J�d�t�F �»�.v!rT�f�����E%�!���5�FRj73B�K����UER�HJ�O  J�� (ڳF���F�q�Y�&T��p�F�z��19�tkvBr��ĄV�h�9p�E�y�<�k�������;�v���"CT��f����)�
� ���)�V	�6���! ��qFF��1q���=� ����O�?�$"���$���je���TCP �Aut�r�<520w H5�J53E1k93��9��96�!�8��9��	 �B57�4��52�Je�(�� Se%!Y������u��ma�Pqtoo�l�ԕ������c�onrel�Ftr�ol Relia'ble�RmvCU!��H51����� a�551e"�CNRE¹I�c��&��it�l\sfutst "UTա��"X�\u��g@��i�6Q]V0�B,Eѝ6A� �Q�)C���X@��Yf�I�1|6s@;6i��T6IU��vR�d�
$e%1��2�C#58�E6��8�Pv�iV4OFH58SOeJ� �mvBM6E~O58 �I�0�E�#+@�&�F �0���F�P6a���)/�++�</N)0\tr�1�����P ,+{�ɶ�rmaski�m#sk�aA���ky'd��h	A	�P�sDis�playIm�`v�����J887 (�"A��+HeůצprCds��I�:���h�0pl�2�R2��:�G9t�@��PRD�TɈ �r�C�@Fm��D�Q�A'scaҦ� V<Q0&��bVvbrl�eۀ�@��^S��&5Uf�j38710�yl	��Uq���7�&�p�p���P^@�P�firm Q����Pp�2�=bk�6��r�3��6��tppl��PL���O�p<b�ac�q	��g1J�U�`�d�J��gait_ 9e��Y�&��Q���	��Shap��era�tion�0��RG67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G���q.F�205p�5S��ɜՁ�retsap�BP��O�\s� "G�CR�ö? �qngda�G��V��s"t2axU��Aa]�Ɔbad�_�btp�utl/�&�e���t�plibB_��=�2�.����5���cir�d�v�slp��x�h3ex��v�re?�Ɵ�x�key�v�pm���x�us$�6�gcr��F������[�q�27j92�v�ol7lismqSk�9O|�ݝ� (pl.��$�t��p!o��29$Fo�8��cg7no@�tp�tcls` CLS0�o�b�\�km�ai_B
�s>�v�o	�t�b���ӿ�E�H���6�1enu501:�[m��utia|$�calmaUR��C�alMateT;R51%�i=1]@-��/ V� ��Z�� �fq1�9 "K9E�L����2m�CLMT�q�S#��et �L�M3!} �F�c�n�spQ�c���c_mioq��� ��c_e������su��ޏ �_� �@�5�G�join��i�j��oX���&c`Wv	 ���N�ve��C�clm�&Ao# �~|$finde�0�STD te�r FiLA�NG���R��
p��n3��z0Cen����r,������J�� ��� ���K��Ú�=���_Ӛ��r� "FNDR�� 3����f��tguid��䙃N�."��J�tq �� �������������J����_������c���	m�Z��\fndr.��n#>
B�2p��Z�CP M1a�����38A��� c��6� (���N� B������� 2�$�81��m_���"ex�z5�.Ӛ��c��bSа�e�fQ��	��RB�T;�OPTN  �+#Q�*$�r*$��*$ r*$%/s#C�d/.,P���/0*ʲDPN`��$���$*�Gr�$�k Exc�'IF��$MASK�%93� H5�%H558��$548 H�$4 -1�$��#1(�$�0 E�$��$-b�$��>�!UPDT �B�4 �b�4�2�49�0�4a��3�9j0"M�49�4�  ��4�4t�psh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4��3�adq\�5K97�9":E�ajO l "DQ^E^�3i�D!q ��4ҲO ?R�? ��q�5��T��32rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F���4��.�5y N� �2i�l(in�4��31� JH1�2Q4�251<ݠ�4rmal� �3)�REo�Z_�æOx�����4��^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg0���4�$HCd\�fͲ �eڱ�4�REM���4�yݱ"u@�RER59�32fO��47Z��5lity,�U��e"�Dil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe� =$�^�
E��u�IAymptm�U��BU��vste�y\�3��m e�b�DvI�[�Qu�:F��Ub�*_�
E,�sIu��_ Er���ox���4huse�E-�?�sn�������8FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��@�b���(��1� ��c��Y�R�� �>� P���W��������'�0ɵ�[��͂����  � ,�+@� �A^�bumpšf��B*�Box%��7A�ǰ60�BBw���MC�� (6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`����)��\bbk96�8 "�4�ω�b5b�9va69����'etbŠ��X����F�ed	�F��u�Lf� �sea"������'�\��,���b�Dѽ�o6�H�
�x�$�f���!y���Q[�! tperr��fd� TPl0o� _Recov,��3|D��R642 � 10��C@}s� N@��(U�rro���y�u2r��  �
�  ����$�$CLe� ��������������$z�_DIGIT\������� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_@�_�_ oo$j��+c�:PRODUCT�M�0\PGSTK�D��V&ohozf9�9��D���$�FEAT_IND�EX��xd���  
�`I�LECOMP ;���#��`�c�SETUP2 �<�e�b� � N �a�c_AP2BCK 1=�i?  �)wh0"?{%&c����Q �xe%�I�m� ��8��\�n���� !���ȏW��{��"� ��F�Տj���w���/� ğS���������B� T��x������=�ү a������,���P�߯ t������9�ο�o� ϓ�(�:�ɿ^��� Ϗϸ�G���k� �� ��6���Z�l��ϐ�� ����U���y���� D���h��ߌ��-��� Q���������@�R� ��v����)�����_� ����*��N��r ��7��m��&�3\�i
pP� 2#p*.cVRc�*���� /��PC�/1/FR6:D/].��/+T�` �/�/F%�/�,�`r/?�*.F�8?	H#&?e<�/�?;STM �2�?�.K ��?�=iPe�ndant Pa'nel�?;H�?@O��7.O�?y?�O:GIF�O�O�5�OoO�O_:JPG _J_�56_��O_�_�	PAN?EL1.DT�_��0�_�_�?O�_2 �_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEIN�S.XML���0\���qCus�tom Tool�bar	��PA?SSWORDy?FRS:\L��� %Passw�ord Config���֏e�Ϗ� B0���T�f������ ����O��s������ >�͟b��[���'��� K��򯁯���:�L� ۯp�����#�5�ʿY� �}��$ϳ�H�׿l� ~�Ϣ�1�����g��� �� ߯���V���z�	� s߰�?���c���
�� .��R�d��߈��� ;�M���q������<� ��`������%���I� �������8���� n���!��W� {"�F�j| �/�Se�� /�/T/�x//�/ �/=/�/a/�/?�/,? �/P?�/�/�??�?9? �?�?o?O�?(O:O�? ^O�?�O�O#O�OGO�O kO}O_�O6_�O/_l_ �O�__�_�_U_�_y_ o o�_Do�_ho�_	o �o-o�oQo�o�o�o �o@R�ov�� ;�_���*�� N��G������7�̏ ޏm����&�8�Ǐ\� 돀��!���E�ڟi� ӟ���4�ßX�j��� �����įS��w��𛯭�B�#��$FI�LE_DGBCK� 1=��/���� (� �)
SUMM?ARY.DGL���OMD:������Diag Su�mmary��Ϊ
CONSLOG��������D�ӱCo�nsole lo�gE�ͫ��MEMCHECK:�!ϯ����X�Memor?y Data��ѧ߁{)��HADOW�ϣϵ�J����Shadow ChangesM��'�-��)	F�TP7Ϥ�3ߨ����Z�mment T�BD��ѧ0=4)�ETHERNE�T�������T�ӱ�Ethernet� \�figura�tionU�ؠ��DCSVRF�߽߫������%�� v�erify alyl��'�1PY���DIFF�����[����%��dif!f]������1R�9�K��� ���{X��CHGD������c��r���2ZAS� 1��GD����k��z��F�Y3bI[� 1�/"GD����s/����/*&�UPDATES.�� �/��FRS:�\�/�-ԱUpd�ates Lis�t�/��PSRBW�LD.CM(?����"<?�/Y�PS_R?OBOWEL��̯ �?�?��?&�O-O�? QO�?uOOnO�O:O�O ^O�O_�O)_�OM___ �O�__�_�_H_�_l_ o�_�_7o�_[o�_lo �o o�oDo�o�ozo �o3E�oi�o� ��R�v��� A��e�w����*��� я`���������O� ޏs������8�͟\� ����'���K�]�� �����4���ۯj��� ���5�įY��}��� ���B�׿�x�Ϝ� 1���*�g�����Ϝ� ��P���t�	�ߪ�?� ��c�u�ߙ�(߽�L� ���߂���(�M��� q� ���6���Z��� ���%���I���B�� ���2�����h����$FILE_� {PR� ��������MDONLY 1�=.�� 
 ���q������� ���~%�I� m�2��h ��!/�./W/�{/ 
/�/�/@/�/d/�/? �//?�/S?e?�/�?? �?<?�?�?r?O�?+O =O�?aO�?�O�O&O�O JO�O�O�O_�O9_�O�F_o_
VISBC�KL6[*.V�Dv_�_.PFR:�\�_�^.PVi�sion VD file�_�O4oFo \_joT_�oo�o�oSo �owo�oB�of �o�+���� ���+�P��t�� ����9�Ώ]�򏁏�� (���L�^������� 5���ܟk� ���$�6� şZ��~�����
�MR_GRP 1�>.L��C4�  B���	 �W�����*u����RHB� ��2 ���� ��� ��� B�����Z�l���C����D�������Ŀ��J�8�L�8�J�� F�5U���R�p���ֿ �Gn�E���.E88�-���:u�{@ �����@A�A���)f�?h!A��تr��E�� F@ ������ھ���NJk�H�9�Hu��F!��IP�s��?����(�9�<�9�89�6C'6<,6\b��+�&�(��a�L߅�p�A��A� �߲�v���r������ 
�C�.�@�y�d��� �����������?��Z�lϖ�BH�� A�Ζ�������
0��PJ��P�K�0��ܿ� �B���/ ���@�33:���.�gN�UUU�U���q	>u.�?!rX��	��-=[z�=��̽=V6<��=�=�=$�q�����@8��i7G��8��D�8@9!�7�:�����D�@ D�� �Cϥ��C������'/0-��P/��� �/N��/r��/���/� ??;?&?_?J?\?�? �?�?�?�?�?O�?O 7O"O[OFOOjO�O�O �O�O�гߵ��O$_�O H_3_l_W_�_{_�_�_ �_�_�_o�_2ooVo hoSo�owo�o�i��o �o�o��);�o_ J�j����� ��%��5�[�F�� j�����Ǐ���֏� !��E�0�i�{�B/�� f/�/�/�/���/��/ A�\�e�P���t����� ���ί��+��O� :�s�^�p�����Ϳ�� �ܿ� ��OH��o� 
ϓ�~ϷϢ������� ���5� �Y�D�}�h� �߳ߞ��������o� 1�C�U�y��߉�� �����������-�� Q�<�u�`��������� ������;&_ J\�������� ��ڟ�F�j4� �������� !//1/W/B/{/f/�/ �/�/�/�/�/�/?? A?,?e?,φ?P�q?�? �?�?�?O�?+OOOO :OLO�OpO�O�O�O�O �O�O_'__K_�o_ �_�_�_l��_0_�_�_ �_#o
oGo.okoVoho �o�o�o�o�o�o�o C.gR�v� ����	���<� `�*<��`��� ��ޏ��)��M�8� q�\�������˟��� ڟ���7�"�[�F�X� ��|���|?֯�?���� �3��W�B�{�f��� ��ÿ��������� A�,�e�P�uϛ�b_�� ���Ϫ_��߀�=�(� a�s�Zߗ�~߻ߦ��� ����� �9�$�]�H� ��l���������� ��#��G�Y� �B��� ����z�������
ԏ :�C.gRd�� ����	�? *cN�r��� ��/̯&/�M/� q/\/�/�/�/�/�/�/ �/?�/7?"?4?m?X? �?|?�?�?�?�?��O !O3O��WOiO�?�OxO �O�O�O�O�O_�O/_ _S_>_P_�_t_�_�_ �_�_�_�_o+ooOo :oso^o�o�op��o��  ��$��o �o�~����� ��5� �Y�D�}�h� ������׏���� 
�C�.�/v�<���8� �����П����?� *�c�N���r������� �̯��)��?9�_� q���JO�����ݿȿ ��%�7��[�F�� jϣώ��ϲ������� !��E�0�i�T�yߟ� ���߮��߮o�o��o >�t�>��b�� ���������+��O� :�L���p��������� ����'K6o Z�Z�|�~���� �5 YDi� z������/ 
//U/@/y/@��/�/ �/�/���/^/??? Q?8?u?\?�?�?�?�? �?�?�?OO;O&O8O qO\O�O�O�O�O�O�O��O_�O7_��$F�NO ����VQ��
F0fQ kP F�LAG8�(LRR�M_CHKTYP�  WP��^Pk�WP�{QOM�P�_MIN�P���}�P�  XNP�SSB_CFG �?VU ��_���S oo�IUTP_DEF__OW  ��R>&hIRCOM�P8o��$GENOVRoD_DO�V�6�nflTHR�V d�e�dkd_ENBWo �k`RAVC_G�RP 1@�WCa X"_�o_1 U<y�r��� ��	��-��=�c� J���n��������ȏ ����;�"�_�F�X�\��ibROU�`FVX.�P�&�<b>&�8�?������������  �D?�јs���@@g�B�7�p�)�ԙ����`SMT�cG�m�M���� �LQHOS�TC�R1H���Ps��at�SM���f�\���	_127.0��1��  e��ٿ��� ��ǿ@�R�d�vϙ��0�*�	anonymous�������ό���0�[�� � �����r����ߨ� ������-���&�8� [�I�π������ ���1�C��W�y��� `�r������ߺ����� ��%�c�u�J\n ��������� M�"4FX��i� �����7// 0/B/T/���m/� �/�/�/??,?�/ P?b?t?�?�/�?��? �?�?OOe/w/�/�/ �?�O�/�O�O�O�O�O =?_$_6_H_kOY_�? �_�_�_�_�_'O9OKO ]O__Do�Ohozo�o�o �o�O�o�o�o
?o }_Rdv���_�_ oo!�Uo*�<�N� `�r��o������̏ޏ �?Q&�8�J�\���~>�ENT 1I��� P!􏪟  ����՟ğ���� ���A��M�(�v��� ^�����㯦��ʯ+� � �a�$���H���l� Ϳ�����ƿ'��K� �o�2�hϥϔ��ό� �ϰ�������F�k� .ߏ�R߳�v��ߚ��� ����1���U��y�<�QUICC0��b�t����1�����%���2&���u�!ROUTERv��R�d���!PCJ�OG����!1�92.168.0�.10��w�NAM�E !��!R�OBOTp�S_�CFG 1H��� �Au�to-start{ed�tFTP�������  2D��hz�� ��U��
//./A�#����~/� ���/�/�/�/� ? 2?D?V?h?�/?�?�? �?�?�?�?���@O ?dO�/�O�O�O�O�? �O�O__*_MON_�O r_�_�_�_�_	OO-O �_A_&ouOJo\ono�o �o=o�o�o�o�oo �o4FXj|�_�_ �_o�7o��0� B�T�#x�������� ��e�����,�>�� ���ŏ���Ο�� ����:�L�^�p� ����'���ʯܯ� � O�a�s�����l����� ����ƿؿ����� � 2�D�g��zόϞϰ� ���#�5�G�I��}� R�d�v߈ߚ�iϾ��� �����)߫�<�N�`��r��XST_ER�R J5
���P�DUSIZ  j��^J����>��?WRD ?t���  guest}��%�7��I�[�m�$SCDMNGRP 2Ktw�������V$�K�� 	�P01.14 8~��   y�����B   � ;����� ����������
 �������?�����~����C.gR|����  i  ��  
��������� +�������
���l �.r���"�l��� m
d����|��_GROU��]L�� �	�����07EQUPD'  	պ�J��TYa ����T�TP_AUTH �1M�� <!iPendany���6�Y!K?AREL:*��
-KC///A/ �VISION �SETT�/v/� "�/�/�/#�/�/
? ?Q?(?:?�?^?p>�CTRL N�����5�
�F�FF9E3�?��FRS:DEFA�ULT�<FA�NUC Web �Server�:
 �����<kO}O�O�O��O�O��WR_CONFIG O��� �?��IDL_CPU_PC@��B��7P�BHUMIN(\��<T?GNR_IO�������PNPT_S_IM_DOmVw[�TPMODNTO�LmV �]_PRT�Y�X7RTOLNK 1P����_o�!o3oEoWoio�RMA�STElP��R�O�_CFG�o�iUO���o�bCYCLE��o�d@_ASG s1Q����
 ko ,>Pbt��� ������sk�bNUM����K@�`�IPCH�o��`R?TRY_CN@oR<��bSCRN����Q��� �b�`�b�R���Տ��$J�23_DSP_E�N	����OB�PROC�U�iJ[OGP1SY@��?8�?�!�T��!�?*�POSRE��zVKANJI_@�`��o_�� ��T�L��6͕����CL_�LGP<�_���EYL_OGGIN�`�����LANGU�AGE YF7ReD w���LG��YU�?⧈�x� ������=P��'�0��$ NM�C:\RSCH\�00\��LN_D?ISP V��
�0�������OC�R.R;DzVT=#�K@9�BOOK W
{���i��ii��X �����ǿٿ����1�"��6	h������e�?�G_BU_FF 1X�]��2	աϸ����� ������!�N�E�W� ��{ߍߺ߱�����������J���DC�S Zr� =����^�+�ZE���������a�IO 1[�
{ ُ!� � !�1�C�U�i�y����� ����������	- AQcu��������EfPTM  �d�2/ASe w������� //+/=/O/a/s/�/8�/��SEV���]�TYP`�/??y͒�RS@�"��×�FL 1\
������?�?�?`�?�?�?�?/?TP6���">�NGN�AM�ե�U`�UP�S��GI}�𑪅�mA_LOAD�G� %�%DF_MOTN���O�@�MAXUALRM <��J��@sA�Q����QWS ��@C �]m�@-_���MP2�7�^
{� ر�	�!�P�+ʠ�;_/��R1r�W�_�WU�W�_ ��R	o�_o?o"oco Noso�o�o�o�o�o�o �o�o;&Kq\ �x������ �#�I�4�m�P���|� ��Ǐ���֏��!�� E�(�i�T�f�����ß ��ӟ���� �A�,� >�w�Z�������ѯ�� ��د���O�2�s� ^�������Ϳ���ܿ��'��BD_LDX�DISAX@	��M�EMO_APR@E� ?�+
  � *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT ��Q�c�Ϝ߇��ߧ� ����w����>�)�b� t�[����{����� �����:���I�[�/� �����������o��� ��6!ZlS� �s����2 �AS'�w�� ��g��.//R/�d/�_MSTR �`�-w%SCD 1am͠L/�/H/�/ �/?�/2??/?h?S? �?w?�?�?�?�?�?
O �?.OORO=OvOaO�O �O�O�O�O�O�O__ <_'_L_r_]_�_�_�_ �_�_�_o�_�_8o#o \oGo�oko�o�o�o�o �o�o�o"F1j Ug������ ���B�-�f�Q����u�����ҏh/MKC_FG b�-�~�"LTARM_���cL�� �σQ�N�<�METsPUI�ǂ���)�NDSP_CMN�Th���|�  	d�.��ς�ҟܔ�|�POSCF�����PSTOL 1�e'�4@�<#�
5�́5�E�S�1�S� U�g�������߯��ӯ ���	�K�-�?���c��u�����|�SING_CHK  ��^;�ODAQ,�f���Ç��DEV }	L�	MC:!̟HSIZEh��-���TASK %�6�%$123456789 �Ϡ��TRIG 1g�+ l6�%���ǃ`�����8�p�YP[�� ��EM_INF� 1h3� �`)AT&�FV0E0"ߙ�)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ������H�����A���AI�q�,��|���� ���ߵ�����J� ��n������W����� ������"����X� �/����e��� ���0�T;x� =�as��/� ,/c=/b/�/A/�/ �/�/�/��?�� �^?p?#/�?�/�?s? }/�?�?O�?6OHO�/ lO?1?C?U?�Oy?�O �O3O _�?D_�OU_z_�a_�_�ONITO�R��G ?5�  � 	EXEC�1Ƀ�R2�X3�X4��X5�X���V7�X8
�X9Ƀ�RhBLd�R Ld�RLd�RLd
bLdb Ld"bLd.bLd:bLdFb�Lc2Sh2_h2kh2�wh2�h2�h2�h2��h2�h2�h3Sh3�_h3�R�R_GRP_SV 1in�z��(ͅ�
�Åo��ۯ_MOx��_D=R^��PL_NAME !6���p�!Def�ault Per�sonality� (from FwD) �RR2eq� 1j)TUX)�TX��q��X d Ϗ8�J�\�n������� ��ȏڏ����"�4��F�X�j�|������2 '�П�����*�<�N�`�r��<������ ��ү�����,�>��P�b� �Rdr 1o��y �\�, ��3���� @D7�  ��?������?䰺��A'�6x����;�	lʲ�	 �x7J������ �< ��"�� �(pK��K ��K�=*�J���J?���JV���Z�����rτ́p�@j�@T;f���f��ұ]�lï�I��p������������b��3���´  �
`��>����bϸ�z���꜐r�Jm��
� B�H�˱]Ӱ�t�q�	� p_�  P�pQ�p}��p|  Ъ��g���c�	'� �� ��I� ��  ����:��È
�È=̣��"�s��	�В�I  �n �@B�cΤ�\��ۤ���tq�y߁rN��� � '�����@2?��@������/�C��C�C�G@ C������O
�A�W�@<�UP�R�
h�B�"b�A��j�����:���Dz۩��߹������j��( �� -���C���'�7������q�Y����� �?�ff ��gy> ����Ёq:a��
>+�  	PƱj�(�����7	���|�?�嚧�xZ�p<
6�b<߈;܍��<�ê<� <�&Jσ��AI�ɳ+���?f7ff?I�?&�k��@�.��J<?�`�q�.� ˴fɺ�/��5/��� �j/U/�/y/�/�/�/��/�/?�/0?q��F�?l??�?/�?�+)�?�?�E�� �E�I�G+� F��?)O�?9O_OJO��OnO�Of�BL޳B �?_h�.��O�O��%_ �OL_�?m_�?�__�_��_�_�_�
�h��<�g>��_Co��_goRodo�o�GA��ds�q�C�o�o�o|����$]H�q���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?�$��?�K�0±�
=ç>�����3�W
=�#��W��e��9������{�����<��(��B�u��=�B0�������	L��H�F��G���G���H�U`E����C�+���I#��I��HD��F��E���RC�j=��
�I��@H��!H�( E<YD0q�$�� H�3�l�W���{����� ���՟���2��V� A�z���w�����ԯ�� ������R�=�v� a������������߿ ��<�'�`�Kτ�o� �Ϻϥ��������&� �J�\�G߀�kߤߏ� �߳�������"��F� 1�j�U��y����� �������0��T�?��Q����(�1���3/E�����5�������q3�8������q4Mgs8&IB+2D��a���{� ^^	������JuP2P7Q4_�A��M0bt��R������/   �/�b/P/ �/t/�/ *a)_3/�/�/�%1a?�/?p;?M?_?q?  �?��/�?�?�?�?O 2� F�$�vGb	�/�A��@�a�`�qC��C@�o�O2��~�OF� DzH@��� F�P DC���O�O�ys<O�!_3_E_W_i_s?̯��@@pZ.tR22!2~
 p_�_�_�_	o o-o?oQocouo�o�op�o�o��Q ��+���1��$MS�KCFMAP  ��5� ��6�Q�Q"~�cON�REL  
�q3�bEXCFENB?w
s1uXq�FNC_QtJOG_OVLIM?wdIp�Mrd�bKEY?w��u�bRUN�|��u�bSFSPD�TY�avJu3sSI�GN?QtT1MO�T�Nq�b_CE_GRP 1p�5s\r���j��� ��T��⏙������ <��`��U���M��� ̟��🧟�&�ݟJ� �C���7�������گ��������4�V�`T�COM_CFG 1q}�Vp�����}
P�_ARC_\r�
jyUAP_C�PL��ntNOCH�ECK ?{ 	r��1� C�U�g�yϋϝϯ����������	��({NO_WAIT_L�l	uM�NTX�r{z�[m�_ERRY�s2sy3� &�������r�c� �^�T_MO��t��,  �
$�k�3�_PARAM��u{��V[��!�u?��� =9@345678901��&� ��E�W�3�c�����{�0������ �����=�UM_RSPACE �Vv���$ODRDSP����jxOFFSE?T_CARTܿ��DIS��PEN_FILE� �q���c֮�OPTION�_IO��PWO_RK v_�msC �P(�R$0puj.j	 ��H�j(6$� RG_DSBL  �5�Js�\��RIE�NTTO>p9!C���Pq=#�UT_SIM_D�
r�b� V� LCT ww�bc��|U)+$_PEXE�d&RATp �vju�p���2X�j)TUX�)TX�##X d-�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O�H2�/oO�O�O�O�O@�O�O�O�O_]�<^O ;_M___q_�_�_�_�_��_�_�_o���X�O�U[�o(��(����$o�,� ��IpB` @oD�  Ua?�[cbAa?��]a]�DWcxUa쪋l;�	lmb��`�x�J�`�����a�< ��`�� ��b, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�b���� �N U�B[�'!o�:q�pC\�C�@@sBq�|���= m�
�A\��h@ߐ�n����Z��B\��A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�'!��(p �?�ffo��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��W ��Ӱ�|�ɆDT Qy-����D � ��,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�T�(�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_j��_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ�_ ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������//�"#�$PGTRA�CELEN  �#!  ���" �8&_UP z���g!�o S!h 8!_�CFG {g%Q#"!x!�$J �#�|"DEFSPD �|�,!!J ��8 IN TRL +}�-" 8�%�!�PE_CONFI�� ~g%��g!�$�%�$LID�#�-74GRP� 1�7Q!��#!A ���&f�f"!A+33D��� D]� C�O� A@+6�!�" �d�$�9�9*1*0� 	 +9�(�&�"��? ´	C�?�;B @3AO�?OIO3OmO�"!>�T?�
�5�O�O�N�O =?��=#�
�O_ �O_J_5_n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_ Roxoco�o�o�o�o�o �o�o>)bM���;
V7.1�0beta1�$�  A�E>�rӻ�A " �p�?!G��q>�嚻r��0�q��޻qBQ��qA\��p�q�4�q�p�"�BȔ2�D�V�h�w�!�p�?�?)2{ȏ w�׏���4��1� j�U���y�����֟�� ����0��T�?�x� c�������ү����!o �,�ۯP�;�M���q� ����ο���ݿ�(π�L�7�p�+9��sF@ �ɣͷϥ�g% ������+�!6I�[� �������ߵߠ����� ����!��E�0�B�{� f����������� ��A�,�e�P���t� ����������� =(aL^��� ����'9$ ]�Ϛ��ϖ����� ��/<�5/`�r߄� �ߏ/>�/�/�/�/�/ ?�/1??U?@?R?�? v?�?�?�?�?�?�?O -OOQO<OuO`O�O�O �O�O���O_�O)__ M_8_q_\_n_�_�_�_ �_�_�_o�_7oIot ���o�o���o�o �o(/!L/^/p/�/{ *o������� ��A�,�e�P�b��� �������Ώ��+� =�(�a�L���p����� �Oߟ񟠟� �9�$� ]�H���l�~�����ۯ Ư���#�No`oro�o n��o�o�o�oԿ�� �8J\ng���� vϯϚ�������	��� -��Q�<�u�`�r߫� ���ߺ�������;� M�8�q�\�������� z������%��I�4� m�X���|��������� ��:�L�^���Z�� ���������$� 6�H�Swb� ������// =/(/a/L/�/p/�/�/ �/�/�/?�/'??K? ]?H?�?��?�?f?�? �?�?O�?5O OYODO }OhO�O�O�O�O�O�O &8J4_F_��� �_�_��_�_"4 -o�O*ocoNo�oro�o �o�o�o�o�o) M8q\���� �����7�"�[� m��?����R�Ǐ��� ֏�!��E�0�i�T� ��x��������_$_ V_ �2�l_~_�_������R�$PLID_�KNOW_M  ��T�|����SV ��U�͠�U ��
��.�ǟR�=�O������mӣM_GROP 1��!`0u���T@ٰo�ҵ�
���Pзj��` ���!�J�_�W�i�{� �ϟϱ����������V��MR�����T��s�w� s��ߠ޴� �߅��ߩ߻�����A� ��'������ ��������=��� #���������}�������S��ST��1 1Ն�U# ���0�_ A .��,> Pb������ ��3(iL^�p�����2r*���<-/�3/)/;/M/4 f/x/�/�/5�/�/�/�/6??(?:?�7S?e?w?�?8�?�?�?�?MAD  d#`�PARNUM  �w�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a��OT_CMP_0��B@�P@'˥T�ER_CHK'U���˪?R$_6[RS8l�¯��_MOA@�_�U_�_RE_RES_G ��>�o o8o+o\oOo�oso�o �o�o�o�o�o�o�W �\�_%�Ue B af�S� ����S 0����SR0�� #��S�0>�]�b��S�0�}������RV 1�x����rB@c]��}t�(@c\��}��D@c[�$����RTHR_IN�Rl�DA��˥d,�M�ASS9� ZM�M�N8�k�MON_QUEUE ���X˦��x� RDNP�UbQN{�P[��ENqD���_ڙEXE韌ڕ�@BE�ʟ��O�PTIOǗ�[��P�ROGRAM %��%��ۏ�O��?TASK_IAD0�OCFG ���xtO��ŠDATA��]�Ϋ@��27� >�P�b�t���,����� ɿۿ�����#�5�G�^��INFOUӌ�������ϭϿ����� ����+�=�O�a�s� �ߗߩ߻��������4^�jč� yġ~?PDIT �ί|c���WERFL
���
RGADJ ��n�A����?�����@���IORI�TY{�QV���MPGDSPH�����Uz�y���OTOEy��1�R� (!�AF4�E�P]����!tcph����!ud��!�icm��ݏ6�XYm_ȡ�R��ۡ)� *+/ ۠�W:F�j ������%@7[B�*��OPORT#�BC۠�����_CAR�TREP
�R� S�KSTAz��ZSS�AV���n�	2500H863��P�r�$!�R����q�n�}/�/�'^� URGE�B��6rYWF� DO{�r�UVWV��$�A�WR�UP_DELAY� �R��$R_HOTk��%O]?�$�R_NORMAL�k�L?�?p6SEMI�?�?�?3AQSKI�P!�n�l#x 	1/+O+ OROdO vO9Hn��O�G�O�O�O �O�O_�O_D_V_h_ ._�_z_�_�_�_�_�_ 
o�_.o@oRoovodo �o�o�o�o�o�o�o *<Lr`����n��$RCVT�M�����pDC�R!�LЈqC�`N�C���C��Q?��>r��<|�{4M��g�&��/���Z��t�����l4�{��4Oi��O <
6�b<߈;܍��>u.�?!<�&{�b�ˏ ݏ��8�����,�>� P�b�t���������Ο ���ݟ��:�%�7� p�S������ʯܯ�  ��$�6�H�Z�l�~� ������ƿ���տ� ��2�D�'�h�zϽ��� ����������
��.� @�R�d�Oψߚ߅߾� ����������<�N� ��r��������� ����&�8�#�\�G� ����}����������� S�4FXj|� �������� 0T?x�u� ���'//,/>/ P/b/t/�/�/�/�/�/ �/�?�/(??L?7? p?�?e?�?�?��?�?  OO$O6OHOZOlO~O �O�O�?�?�O�O�O�O  __D_V_9_z_�_�? �_�_�_�_�_
oo.o�@oRodovo�X�qGN_ATC 1��� AT&�FV0E0�k�ATDP/6/9�/2/9�hAT�A�n,AT�%G1%B960��i+++�o,��aH,�qIO_TYPE  �u��sn_�oREFP�OS1 1�P{O x�o�Xh_ �d_�����K� 6�o�
���.���R�����{{2 1�P{ ���؏V�ԏz����q3 1��$�6�p���ٟ���S4 1�����˟���n���>%�S5 1�<�N��`�����<���S6 1�ѯ���/������ѿO�S7 1� f�x���ĿB�-�f��S8 1������Y�������y�SMA�SK 1�P  q
9�G��XNOM����a~߈ӁqMO�TE  hܗ�_CFG ���������rPL_RANG�ћQ����OWER� ��e���S�M_DRYPRG %i�%��J��TART �
��X�UME_PRO�'�9��~t_EXE�C_ENB  <�e��GSPD����8��c��TDB���sRM��MT_!��T�ߓaOBOT�_NAME �i���iOB_O�RD_NUM ?�
�\qH?863  �T���������bPC_TIMEOUT��{ x�`S232���1��k L�TEACH PE�NDAN �ǅ��}���`Mai�ntenance Cons�R}�m
�"{�dKCL/!Cg��Z ��n�� No Us�e}�	��*NPqO��х��ӽ(CH_L����]���	�mMAVAIL��{����SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�M7��%aR  ��ϰ�P{_��P_INTVAL��@����JR_OPoTION�V �E�BpVAT_GR�P 2�����(y_Ho � e_vo�o�oYo�o�o�o �o�o*<�bOo NDpw����� �	���?�Q�c�u� ����/���ϏᏣ��� �)�;���_�q����� ����O�ɟ���՟ 7�I�[�m�/������� ǯٯ믁��!�3��� C�i�{���O���ÿտ ���ϡ�/�A�S�e� 'ωϛϭ�oρ����� ��+�=���a�s߅� Gߕ߻����ߡ��� '�9�K�]��߁��� ��y����������5��G�Y��E�$SCAN_TIM�AYue�w�R �(ӿ#((�<0.a�aPaP
Tq>��Q��oa�����OOE2/���d;D2BaR��WY���^���^R^	r � P��� �  8�P�	<�D��G Yk}���������Qp�/@/R//)P;��o\T��Qpg-�t�_DiKT|��[  � l v%������/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OWW�#�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_olO~Od+No`o ro�o�o�o�o�o�o�o &8J\n�������u�  0�"0g�/�-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ����$o��˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�����Do������ ��ҿ�����,�>� P�b�tφϘϪϼ���`������w
�  5 8�J�\�n߀ߒߜկ� ��������	��-�?�Q�c�u����� ��-����� � 2�D�V�h�z��������������������& ��%	�12345678^�" 	��/� `r��������(: L^p����� �� //$/6/H/Z/ l/~/��/�/�/�/�/ �/? ?2?D?V?h?�/ �?�?�?�?�?�?�?
O O.O@Oo?dOvO�O�O �O�O�O�O�O__*_ YON_`_r_�_�_�_�_ �_�_�_ooC_8oJo \ono�o�o�o�o�o�o �oo"4FXj�|������� ��	��s3�E�W��{�Cz  Bp���   ��2����z�$SCR_�GRP 1�(��U8(�\x�^ @ > 	!��	  ׃���"�$� ���-��+��R�w����D~�����#�����O���M-�10iA 890�9905 Ŗ5 M61C >4��J*ׁ
� ����0�����#�1�	�"�z�������¯Ҭ ���c��� O�8�J��������!�����ֿ��B�By���������A��$�  @��<� �R�?��d���Hy�u�O����F@ F�` �§�ʿ�϶������� %��I�4�m��<�l�`�߃ߕߧ߹�B��� \����1��U�@�R� ��v������������;���*<=�
�F���?�d�<�>HE�����@�:��� B���ЗЙ����EL_DEFA�ULT  ���_�B��MIPOWERFL  �$1 oWFDO $���ERVENT �1�����"��pL!DUM_�EIP��8��j!AF_INE <�=�!FT����!��4 ���[!RPC�_MAIN\>�8J�nVISw=y���!TP��PU��	d�?/!�
PMON_PR'OXY@/�e./�/�"Y/�fz/�/!RDM_SRV�/r�	g�/#?!R dC?�h?o?!
p�M�/�i^?�?!?RLSYNC�?8��8�?O!ROS�.L�4�?SO" wO�#DOVO�O�O�O�O �O_�O1_�OU__._ @_�_d_v_�_�_�_�_�o�_?oocoiICE_KL ?%y� (%SVCPRG1ho8��e��D�o�m3�o�o�`4 D�`5(-�`6PU�`7x}�`���l9��{�d:?� �a�o��a�oE��a�o m��a���aB���a j叟a���a�5� �a�]��a����a3� ���a[�՟�a�����a ��%��aӏM��a��u� �a#����aK�ů�as� ��a��mob�`�o�` 8�}�w�������ɿ�� �ؿ���5�G�2�k� VϏ�zϳϞ������� ���1��U�@�y�d� �߯ߚ��߾������ �?�*�Q�u�`��� ����������;� &�_�J���n������������sj_DEV� y	�M{C:(!`OUT",?REC 1�Z� �d   	 	������

 �Z�{ 0H6lZ�~� ����� //D/ 2/h/z/\/�/�/�/�/ �/�/�/?�/,?R?@? v?d?�?�?�?�?�?�? �?OO(ONO<OrOTO fO�O�O�O�O�O�O_ &__J_8_Z_\_n_�_ �_�_�_�_�_�_"oo Fo4oVo|o^o�o�o�o �o�o�o�o0T Bxf����( ���,��P�>�`� ��h���������Ώ� �(�:��^�L���p� ������ܟ���� � 6�$�Z�H�~���r��� ��دƯ����2�� &�h�V���z�����Կ �ȿ
�����.�d� RψϚ�|ϾϬ����� ����<��`�N�p� �߄ߺߨ�������� �8�&�\�J�l��joV 1�w P�l�	� � ��F��
TYP�EVFZN_C�FG �x��d7�GR�P 1�A�c �,B� A� D;� B���  �B4RB2�1HELL:�4(
 X���>�%RSR���� E0iT�x� �����/�Sew�  ��%w������#����)�A�2#�d�����HK 1��� ���m/h/z/�/�/ �/�/�/�/�/
??E? @?R?d?�?�?�?�?��?OMM ����?���FTOV_EN�B ���+�HOW_?REG_UIO��IMWAITB\�JKOUT;F���LITIM;E��ΆOVAL[OMC_U�NITC�F+�MO�N_ALIAS �?e�9 ( he�s_(_:_L_^_�� _�_�_�_�_j_�_�_ oo+o�_Ooaoso�o �oBo�o�o�o�o�o '9K]n�� ��t���#�5� �Y�k�}�����L�ŏ ׏������1�C�U� g����������ӟ~� ��	��-�?��c�u� ������V�ϯ��� ���;�M�_�q���� ����˿ݿ����%� 7�I���m�ϑϣϵ� `�������ߺ�3�E� W�i�{�&ߟ߱����� �ߒ���/�A�S��� w����X������ ����=�O�a�s��� 0������������� '9K]��� �b���#� GYk}�:�� ����/1/C/U/  /f/�/�/�/�/l/�/ �/	??-?�/Q?c?u? �?�?D?�?�?�?�?O �?)O;OMO_O
O�O�O �O�O�OvO�O__%_�7_�C�$SMON�_DEFPRO ����`Q� *S�YSTEM*  �d=OURECA�LL ?}`Y �( �}4cop�y md:prg�state.dg� virt:\t�emp\=>192.168.4�P�46:3892 a2>_�_�_o}3�Uconslog�_��_ �_eowo�oiio�_<oNo�o�o�f�2�Uerrall.ls�o�n�oew�`9�Rfrs:�orderfil�.dat1umpback<Nt�����j0�Tb:*.*�� �b�t���c�6��x9�P873C6 W������.��*.d��ƎϏ`�r�|��e
xyzr�` 61 +�=�O�����e����ӑ�� ҟc�u�����5�͇ ٯ����"���̈ѯ�b�t���c4x��:\)���;�S�U����.
� }5��a���� Άֿg�yϋϞ���9� T�����	����@��� c�u߇ߚ�-�?�п�� ���ϩ߻�N�_�q� ��Ϩ�1�������� �&���J�[�m���� ��7����������"� ��F���i{����+�=O���)�8504 *�cu ����5�6��� �"��5�b/t/�/𙏫���P2164 W/�/�/�/��/�) �/`?r?�?���;?M? �?�?O'�4�?�? cOuO�O��5/�'�O �O�O/"/�O�(�Ob_ t_�_����QCU_�_ �_
o�_�_NQ�_ho zoo�O�O:_�_�o�o 
_�oA_�odv� �_.o;�_���o ��Oo`�r����o�o 2�oޏ���'�K\�n������$S�NPX_ASG �1�������� P 0� '%R[?1]@1.1����?���%֟��&� 	��\�?�f���u��� �����ϯ��"��F� )�;�|�_�������ֿ ��˿���B�%�f� I�[Ϝ�Ϧ��ϵ��� ����,��6�b�E߆� i�{߼ߟ�������� ���L�/�V��e�� �����������6� �+�l�O�v������� ��������2V 9K�o���� ���&R5v Yk�����/ ��<//F/r/U/�/ y/�/�/�/�/?�/&? 	??\???f?�?u?�? �?�?�?�?�?"OOFO )O;O|O_O�O�O�O�O �O�O_�O_B_%_f_ I_[_�__�_�_�_�_ �_�_,oo6oboEo�o io{o�o�o�o�o�o �oL/V�e� �������6� �+�l�O�v��������PARAM ������ �	U��P�����OFT_KB_CFG  ヱ����PIN_SIM  ���C�U�g������RVQSTP/_DSB,�򂣟|����SR �/��� &  UL�TIROBOTT�ASK�����T�OP_ON_ER/R  ����PTN /��@�A	�RI�NG_PRM� ���VDT_GR�P 1�ˉ�  	������������ Я�����*�Q�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߣ� �߲����������� 0�B�i�f�x���� ���������/�,�>� P�b�t����������� ����(:L^ p�������  $6HZ�~ �������/  /G/D/V/h/z/�/�/ �/�/�/�/?
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8___\_���VPRG_COUNT��@���R'ENBU��UM�S���__UPD 1�>/�8  
s_� oo*oSoNo`oro�o �o�o�o�o�o�o+ &8Jsn��� ������"�K� F�X�j���������ۏ ֏���#��0�B�k� f�x���������ҟ�� ����C�>�P�b��� ������ӯί������UYSDEBU)G�P�P�)�d�YH�SP_PASS�U�B?Z�LOG [��U�S)�9#�0�  ��Q)�?
MC:\��6���_MPC���U�$��Qñ8� �Q趿SAV ���ج�ǲ&�ηSV�;�TEM_TIM�E 1��[ (�m��&����}YT1SVGUNS�P֕U'�U���AS�K_OPTIONДP�U�Q�Q��BC?CFG ��[u�� n�A�a�` a�gZo��߃ߕ��߹� ������:�%�^�p� [��������� � ����6�!�Z�E�~�i� ��������&����� ��&8��nY� }�?��ԫ � �(L:p^� ������/ / 6/$/F/l/Z/�/~/�/ �/�/�/�/�/�/2?8  F?X?v?�?�??�? �?�?�?�?O*O<O
O `ONO�OrO�O�O�O�O �O_�O&__J_8_n_ \_~_�_�_�_�_�_�_ o�_ o"o4ojoXo�o D?�o�o�o�o�oxo .TBx��j �������� ,�b�P���t�����Ώ ��ޏ��(��L�:� p�^�������ʟ��� �o��6�H�Z�؟~� l�������د���ʯ  ��D�2�h�V�x�z� ��¿���Կ
���.� �>�d�Rψ�vϬϚ� �Ͼ�������*��N� �f�xߖߨߺ�8��� ������8�J�\�*� ��n���������� ��"��F�4�j�X��� |������������� 0@BT�x� d�����> ,Ntb���� ��/�(//8/:/ L/�/p/�/�/�/�/�/ �/�/$??H?6?l?Z? �?~?�?�?�?�?�?O �&O8OVOhOzO�?�O �O�O�O�O�O
__�O @_._d_R_�_v_�_�_ �_�_�_o�_*ooNo <o^o�oro�o�o�o�o �o�o J8n $O�����X����4�"�X�B�v���$TBCSG_G�RP 2�B��  �v�� 
 ?�   ������׏�������@1��U�g�z���ƈ��d, ���?~v�	 HC��d��>����e�CL  B���Пܘ��w���\)���Y  A�ܟ$�B�g�B�Bl�i�X��ɼ���X��  DA	J���r�����C�����үܬ���D�@ v�=�W�j�}�H�Z����ſ���������v�	V3.0�0��	m61c�	*X�P�u�g�&p�>���v�(:��� ��p͟�  O����p�����z�JCFG �B���� �����������=��=�c�q�K�qߗ߂� �ߦ��������'�� $�]�H��l����� ��������#��G�2� k�V���z��������� �����p*<N ���l����� ��#5GY} h����v�b�� >�// /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?d?R?t?v?�? �?�?�?�?O�?*OO :O`ONO�OrO�O�O� �O�O�O_&__J_8_ n_\_�_�_�_�_�_�_ �_�_�_oFo4ojo|o �o�oZo�o�o�o�o�o �oB0fT�x �������,� �P�>�`�b�t����� Ώ�������&�L� �Od�v���2�����ȟ ʟܟ� �6�$�Z�l� ~���N�����دƯ� � �2��B�h�V��� z�����Կ¿���� .��R�@�v�dϚψ� ���Ͼ�������<� *�L�N�`ߖ߄ߺߨ� ���ߚ�������\� J��n������� ���"���2�X�F�|� j��������������� .TBxf� ������ >,bP�t�� ���/�(//8/ :/L/�/�ߚ/�/�/h/ �/�/�/$??H?6?l? Z?�?�?�?�?�?�?�? O�?ODOVOhO"O4O �O�O�O�O�O�O
_�O _@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<oro`o�o�o�o�o �o�o�o&�/>P �/������ ���4�F�X��(� ��|�����֏���� Ə0��@�B�T���x� ����ҟ������,� �P�>�t�b������� ��������:�(� ^�L�n�������2d �����̿�$�Z�H� ~�lϢϐ��������� �� ��0�2�D�zߌ� �߰�j���������� 
�,�.�@�v�d��� �����������<� *�`�N���r������� ������&J\ �t��B��� ���F4j| ��^����/��  2 6# �6&J/6"�$TB�JOP_GRP �2���?  ?�X,i#��p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�x�'�!�!>���
5�59>�0+1�33=�CL� �fff?+0?�ffB� J1�%Y?d7�.���/>��2�\)?0�5����;��hCY� ��  @� �!B� � A�P?�?�3EC�  D�!�,�0�*BOߦ?�3JB���
:���Bl�0��0�$�1�?O6!?Aə�AДC�1sD�G6�=q�E�6O0�p��B�Q�;�A�� �ٙ�@L3D	��@�@__�O�O>BÏ\JU�OHH�1ts}�A@33@?1� C�� �@�_�_&_8_>��D�UV_0��LP�Q30<{�zR� @�0�V�P!o3o �_<oRifoPo^o�o�o �oRo�o�o�o�oM (�ol�p~���p4�6&�q5	�V3.00�#m761c�$*(��$�1!6�A� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,IR�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^S@;Q��|8�E`rz@/&�8�6&�<��1�w�^$ES�TPARS  �*({ _#HR��AB_LE 1�p+Z�6#|�Q� � 1�|��|�|�5'=!|�	�|�
|�|�˕6!�|�|�|���RDI��z!ʟܟ� ��$���O������ ¯ԯ�����S��x# V���˿ݿ��� %�7�I�[�m�ϑϣ� �����������U-�� ��ĜP�9�K�]�o���-�?�Q�c�u���6�N�UM  �*z!� >  Ȑ�����_CFG ������!@b IMEBF_TT����x#��a�VER��b�w�a�R 1�p+
' (3�6"1 ��  6!����������  �9�$�:�H�Z�l�~� ���������������^$��_��@x�
�b MI_CHAN�m� x� kDBGLV;0o�x�a!n �ETHERAD �?�� �y��$"�\&n ROUmT��!p*!�*�SNMASK��x#�255.�h�fx^$OOL�OFS_DI���[ՠ	ORQCTRL �p+;/�� �/+/=/O/a/s/�/ �/�/�/�/��/�/�/�!?��PE_DET�AI��PON_�SVOFF�33P_MON �H��v�2-9STRTC_HK ����42VTCOMPA�Ta8�24:0FPR�OG %�%�MULTIROB�OTTO!O06�P�LAY��L:_IN�ST_MP GL�7YDUS���?�2L�CK�LPKQUIC�KMEt �O�2SC�RE�@�
tps��2�A�@�I���@_Y���9�	S�R_GRP 1Ҿ� ��� \�l_zZg_�_�_�_�_�_�^�^�oj�Q'O Do/ohoSe��oo�o �o�o�o�o�o! WE{i�������	1234�567��!���X��E1�V[
 �}�ipnl/a�g?en.htmno���������ȏ~�P�anel setup̌}�?��0�B�T�f� ��񏞟 ��ԟ���o���� @�R�d�v������#� Я�����*���ϯ ůr���������̿C� �g��&�8�J�\�n� ����϶��������� uϣϙ�F�X�j�|ߎ� �����;��������0�B��*NUALR�Mb@G ?�� [���������� �� ��%�C�I�z�m�������v�SEV � ����t�E?CFG Ձ=]�/BaA$   B�/D
 ��/C� Wi{�����@�� PRց;C �To\o�I�6?K0(%����0 �����//;/ &/L/q/\/�/�/�/lƇD �Q�/I_��@HIST 1׾�9  ( � ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1 Ec0p?p�?�?�?/C�� >?P=962n?�?
OO0.O�?�?�136c?|O �O�O�OAOSO�?�O_ _0_�O�O_Lu_�_�_ �_:_�/�_�_oo)o ;o�__oqo�o�o�o�o Ho�o�o%7I~��a81�ou��� ���o���)�;� M��q���������ˏ Z�l���%�7�I�[� ��������ǟٟh� ���!�3�E�W���� ������ïկ�v�� �/�A�S�e�Pb�� ����ѿ������+� =�O�a�s�ϗϩϻ� ������ߒ�'�9�K� ]�o߁�ߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y��� v�����������	 �?Qcu��( ����)� M_q���6� ��//%/�I/[/ m//�/�/�/D/�/�/ �/?!?3?�/W?i?{? �?�?�?�����?�?O O/OAOD?eOwO�O�O �O�ONO`O�O__+_ =_O_�Os_�_�_�_�_ �_\_�_oo'o9oKo �_�_�o�o�o�o�o�o jo�o#5GY�o�}������?���$UI_PAN�EDATA 1������  	�}��0�B�T�f�x��� ) ����mt�ۏ���� #�5���Y�@�}���v� ����ן�������1���U�g�N������ �1��Ïȯگ� ���"�u�F���X�|� ������Ŀֿ=���� ��0�T�;�x�_Ϝ� �ϕ��Ϲ������,���M��j�o߁ߓ� �߷������`��#� 5�G�Y�k��ߏ��� �����������C� *�g�y�`��������� F�X�	-?Qc ����߫���� ~;"_F� �|�����/ �7/I/0/m/�����/ �/�/�/�/�/P/!?3? �W?i?{?�?�?�?? �?�?�?O�?/OOSO eOLO�OpO�O�O�O�O �O_z/�/J?O_a_s_ �_�_�_�O�_@?�_o o'o9oKo�_oo�oho �o�o�o�o�o�o�o# 
GY@}d�� &_8_����1�C� �g��_��������ӏ ���^���?�&�c� u�\�������ϟ��� ڟ�)��M����� ������˯ݯ0��� ��7�I�[�m������ ����ٿ�ҿ���3� E�,�i�Pύϟφ���0����Z�l�}���1� C�U�g�yߋ�)߰� #������� ��$�6� ��Z�A�~�e�w��� ��������2��V��h�O�����v�p��$�UI_PANEL�INK 1�v��  ��  ��}12�34567890 ����	-?G � ��o�����a ��#5G�	�����p&���   R�����Z� �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?.O@O ROdOvO�O O�O�O�O �O�O_�O�O<_N_`_0r_�_�_�0,���_ �X�_�_�_ o2ooVo hoKo�ooo�o�o�o�o �o�o��,>r} ��������� ���/�A�S�e�w� �������я���t v�z����=�O�a� s�������0S��ӟ� ��	��-���Q�c�u� ������:�ϯ��� �)���M�_�q����� ����H�ݿ���%� 7�ƿ[�m�ϑϣϵ� D��������!�3�E� �_i�{�
�߂����� �������/��S�e� H���~��R~'�'� a��:�L�^�p��� ������������  ��6HZl~�� �#�5��� 2 D��hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?�/ �?�?�?�?�?�?m?O O&O8OJO\O�?�O�O �O�O�O�O�O[�_�� 4_F_)_j_|___�_�_ �_�_�_�_o�_0oo Tofo��o��o��o �o�o,>1b t����K�� ��(�:����{O ������ʏ܏�uO� $�6�H�Z�l������� ��Ɵ؟����� �2� D�V�h�z�	�����¯ ԯ������.�@�R� d�v��������п� ��ϕ�*�<�N�`�r� ���O�Ϻ�Io������ ���8�J�-�n߀�c� �߇����߽����o 1�oX��o|���� ���������0�B� T�f������������ ��S�e�w�,>Pb t��'���� �:L^p� �#���� // $/�H/Z/l/~/�/�/ 1/�/�/�/�/? ?�/ D?V?h?z?�?�?�??? �?�?�?
OO.O��RO dO�߈OkO�O�O�O�O �O�O_�O<_N_1_r_ �_g_�_7OM�m��$UI_QUI�CKMEN  >��_Ao�bRESTORE� 1�?  �|��Rto�o�im�o�o�o�o �o:L^p� %������o� ���Z�l�~����� E�Ə؏���� �Ï D�V�h�z���7����� ��/���
��.�@�� d�v�������O�Я� ����ßͯ7�I��� m�������̿޿��� �&�8�J��nπϒ� �϶�a�������Y�"� 4�F�X�j�ߎߠ߲� �����ߋ���0�B�T�gSCRE`?�#mu1s]co`u2��3��U4��5��6��7��y8��bUSERq�dv��Tp���ks����4��5��6��7���8��`NDO_�CFG �#k � n` `PDA�TE ����NonebSE�UFRAME  ��TA�n�RTO?L_ABRTy�l�Α�ENB����GR�P 1�ci/aCz  A�����Q@�� $6HR�d��`U�����MSK  �����MNv�%�U�%����bVISCAN�D_MAX�I���FAIL_�IMG� �PݗP#���IMREGN�UM�
,[SI�Z�n`�A�,~VONTMOU��@���2���a��a��~��FR:\� � MC{:\�\LOG�7B@F� !�'/�!+/O/�Uz �MCV�8#U�D1r&EX{+�S|�PPO64_���0'fn6PO��LIb�*�#9V���,f@�'�/�� =	�(SZV��.����'WAI��/STAT 	����P@/�?�?�:�$�?�?��2DW�P  ��P yG@+b=��� H��O_JMPE�RR 1�#k
 � �2345678901dF�ψO{O �O�O�O�O�O_�O*_�_N_A_S_�_
� M�LOWc>
 �_�TI�=�'M�PHASE  ���F��PSHI[FT�1 9�]@<�\�Do�U#oIo �oYoko�o�o�o�o�o �o�o6lCU �y����� �@�	�V�-�e2����	VSFT1�2�	VM�� ��5�1G� ���%A_�  B8̀̀E�@ pكӁ˂�у���z�ME@�?��{��!c>&%�aM�1��k�0�{ �$�`0TDINEND��\�O� �z���S��w��P��=�ϜRELE�Q���Y���\�_ACT�IV��:�R�A ���e���e�:�R�D� ���YBOX� �9�د�6���02���1�90.0.�83v��254�:�QF�	 �X��j��1�ro�bot���  � p�૿�5pc��̿������7�����-�f�ZABC�����,]@U��2 ʿ�eϢωϛϭϿ� ���� ���V�=�zߐa�s߰�E�Z��1� Ѧ