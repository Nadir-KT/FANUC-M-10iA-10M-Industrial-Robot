��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ��&�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�� W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2�� XD�#
 �d $CARD�_EXIST4�$FSSB_TY�PuAHKBD_YS�B�1AGN Gn� $SLOT�_NUMJQPREV,DBU� g1� �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��AETE_OK�RUS�P_CR�Q$;4�V� 0LACIw1�RAP�k �1x@ME@$D�V�Q�Pv�Ah{oQL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa4 hq;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I9�TY!1�@,P*2 �`w@� �!R*�HD�cJ* C��2���3��4��5��6���7��8��94:�qO�$ <� �$6xK3 1w`O_M|�@�C t � �E#6NGP�ABA� �c��ZQ���`����@nr��� ��P��0����x�p��PzPb26����"J��_R��BC�J��3�JVP��tB�S��}Aw��"�tP_�*0OFSzR @�� RO_K8���aIyT�3��NOM_�0Ҝ1ĥ3�ACPT �� $���AxP��K}EX�� �0�g0I01��p�
$TyFa��C$MD3���TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF0�vF�40CPp@�a�2 
P$A`PU8�3N)#�dR�*�AX�!sDETAI�3BUFV��p@�1 |�p۶�pP�IdT� PP[�M�Z�Mg�Ͱj�F[�SIMQSI�"0��A�.�����lw T�p|zM��P�B�F�ACTrbHPEW�7�P1Ӡ��v��MC�d� �$*1JqB�p<�*1DECH����H��(�c� �� +PNS_EMP��$GP���,P!_��3�p�@Pܤ��TC��|r��0�s�� b�0�� �B���!
����JR� ��SEGF�R��Iv �aR�TrkpN&S,�PVF4|��� &k� Bv�u�cu��aE�� !2���+�MQ��E�SIZ�3����T��P���|��aRSINF� ����kq���������LX�����F�CRCMu�3CClpG�� p���O}���b�1����P���2�V�DxIC��C���r����P��{�� EV �zF_J��F�pNB0�?�������A�! � r�Rx����V�lp�2���aR�t�,�g�R>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!�@$SK��2G �� �"�"�@�PR8� 
 ��D���# l>�q1$��$��
+�L9$?(�V�)%@?R4C&_?R4gENE��'~?�(�� RE�pY2(�H �OS��#$L�3$$3R�h�;3�MVOk_D@!V�ROScrr�w�S����CRIGGER�2FPA�S��7�ET�URN0B�cMR_���TUː[��0EkWM%���GN>`���RLA���Eݡ<�P�&$P�t�'�@4a��C�DϣV��DXQ��4�1��MVG�O_AWAYRM�O#�aw!�D�CS_)  `IS#� �� �s 3S�AQ汯 4Rx�@ZSW�AQ�p�@1UW��NcTNTV)�5RV
a����|c�éWƃ��J�B��x0��SAFE�ۥ�V_SV�bEX�CLUU�;��ONL��cYg�~az��OT�a{�HI_V�? �!0Q, M�_ #*�0� ��_z�2�o CdSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc��@Sp�i�a+ �j�f \Ca�pOGIx2,���$F�b�$ѐOT��@A $DUMMY��Ft��Ft±�06U- ` !�HE�|s��~b�c�B@ SUFFI���4PCA��Gs5Cw6CrZ0M�SWU. 8!�KgEYI��5�TM�10�s�qoA�vINޱE�Ca, / D��H7OST�P!4����<���<�°<��p<�E�M'���Z�0SBL�� UL��0  ��	��w��DT��01 � $|��9USAMPL�@��/���決�$ I@|갯 $SUBӄ���w0QS�����#��SAV�����c�S< X9�`�fP$�0E!�� YN_B�#2 M0�`DI�d�pO|��m��#$F�R_I�C� �ENC2s_Sd3  ��< 3�9���� cgp����4�"��2�A9��ޖ5���`ǻ�@Q@K&D-!�a�AVER�q��λ�DSP
���PC�_�q��"�|�ܣ�V7ALU3�HE�(��M�IP)���OP5Pm �TH�*�D�S" T�/�Fb��;�d����d ���&���ET6 }H(rLL_DUǀ��a�@��k���֠O�T�"U�/��o�@@N_OAUTO70�C$}�x�~�@s��*|�Cp��C� 2�iaz�L�� 8/H *��L� � ��Բ@sv��`� �� � ����Xq��cq���q��T�q��7��8��9���0���1�1 �1�-�1:�1G�1T�1*a�1n�2|�2��U2 �2-�2:�2G�U2T�2a�2n�3|ʥ3�3� �3-�3�:�3G�3T�3a�3�n�4|�v�����9� <���z�ΓKI`����H硵��FEq@�{@: ,��&a?g P_P?��>�����E�@��ia�QQ��;fp$T�P�$VARI�����,�UP2Q`< W�߃TD��g�����`������q��BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P�"�l@``>t� ;��6����ST����T��M ����0	��i���F����������kRt ����F?ORCEUP�b܂�FLUS
pH(N𒰚 ��6bD_CM�@E�7N� (�v\�P��REM� Fa���@j���
Kr�	N���EFF/�̎�@IN�QOVܣ�OVA�	TR3OV DT)��DTMX:e �P :/��Pq�vXpCLN _�p��@ �2�	_|��_T: �*|�&PA�QDI���1��0�Y0RQm�_+qH���M���CL�d#�R�IV{�ϓN"EAR6/�IO�PCP��2BR��CM�@N �1b 3GCLF��!DY�(��a�#5T�DG���� :�%��FSS� )��? P(q1�1��`_1"811�E�C13D;5D6�GSRA���@�����PW�ON2EBUG�S�2�C`g�ϐ_E A x��@a��TERM�59B�5�qORIw�0C�9SM_-`���0�D�:A�9E�5����UP��F�3 -QϒA�P�3>�@B$SEGGJ� �EL�UUSEPNFI��pBx��1@�<�4>DC$UF�P���$���Q�@C����G�0T�����SN;STj�PATۡg���APTHJ�A�E *�Z%qB\`F�{E��F��q�pARxPY�aSH�FT͢qA�AX_SGHOR$�>��6 @�$GqPE���OV�R���aZPI@P@$Uz?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi�[Y )��G�@R��i�e���i�R�!P�uASY1M���uqAWJ�G)��E��Q7i�RD�U�[d�@i�U��C�%UP����P���WOR�@Mv��k0SMT���G��GR��3�aP�A�@��p5�'�H ׸ j�A�TO�CjA7pP]Pp$OPd�O��C�%�pe�O!��RE.p�R�C�AO�?��Be5pR�EruIx'QG��e$PWR) IM�du�RR_$s  ��b�B Iz2H|8�=�_ADDRH�?H_LENG�B�q��q:�x�R��So�J6.�SS��SK���`��� ��-�SE*ܕ�$��HSN�MN1K	�j�5�@r�֣OL��\�WpW�<Q�>pACRO�p�� �@H ����Q� ��OUPW3�b_>�I��!q�a1������ ��|��������-����:���iIOX2S�=�D�e��]����L $��p�!_O�FF[r_�PRM_���aTTP_��H��M (�pOcBJ�"�pG�$H��LE�C��ٰN � 9�*�AB_�T��
�S�`�S��LV��KRW"duH�ITCOU?BGi�LO�q����`d� Fpk�GpSS� ����HWh�wA��O�.��`INCPU>X2VISIO��!���¢.�á<�á-� ��IOLN)�P �87�R'�[p$S�L�bd PUT_&��$dp�Pz ��� F_AS2Q/�$LD���D�aQ"T U�0]P�A������PHYG灱Z���5�UO� 3R ` F���H�Yq�Yx�ɱvpP�Sdp���x��,ٶ%�UJ��S����;NE�WJOG�G �'DIS��&�KĠ��&3T |��AV��`�_�CTR!S^�FL�AGf2&�LG�dU� �n�:��3LG_SIZ��ň�X��=���FD��I�� ��Z �ǳ��0�Ʋ�@s ��-ֈ�-�=�-���-�x�0-�ISCH_��Dq��N?���V���EE!2�C��n�Uȡ����`L�Ӕ�DAU��EA��Ġt�����GHr��I�BO}O)�WL ?`��� ITV���0\�R;EC�SCRf 0��a�D^�����MARG��`!P�)�T�/ty�$?I�S�H�WW�I�ܩ�T�JGM��MN�CH��I�FNKEuY��K��PRG���UF��P��FWDv��HL�STP���V��@�����RS"S�H�` �Q�C�T1� ZbT�R ���U����@��|R��t�i���G��8PPO��6�F�1�Mޘ�FOCU��RG�EXP�TUI��IЈ�c��n��n ����ePf���!p6�ePr7�N���CANAI��jB��VAIL��C�Lt!;eDCS_H!I�4�.��O�|!"�S Sn�y�0I�BUFF1�XY��PT�$��� �v��fĘ�1�A
�rYY��P ������pOS1�2�3���0Z � � ��aiE�*��IKDX�dP�RhrO�X+��A&ST��R���Yz�<! Y$EK&CK+���Z&m&�OS�5�0[ L��o�0��]PL�6p wq�t^����t�0��7�?_ \ �`�Р瀰�7��#�0C��]{ ��CLDP��>;eTRQLI�jd8.�094FLGz�0�r1R3�DM�R7��LqDR5<4R5ORG.� ��e2(`���V�8.��T8<�4�d^ �q�<4(��-4R5S�`T00m���0DFRCLM�C!D�?�?3I@��M9IC��d_ d����RQm�q�DSTB	�  �Fg�H�AX;b �H�LE/XCESZr�� rB)Mup�a`��B;dP��rB`��`a��F_A�J��$[�O�H0K�db \��ӂS�7$MB��LIБ}S?REQUIR�R>qx�\Á�XDEBU��*oAL� MP�c�ba���P؃ӂ!BoAND���`�`d�҆�c�c3DC1��IN�����`@�(h?Nz�@q��o��UPST8� �e�rLOC�RYI�p�EX�fA�px��A�AODAQP�7f X��ON��[rMF�����f)�"I�`�%�e��T���FX�@�IGG� g �q��"E�0��#���$R�a%;#7y��Gx�VvCPi�DATAw�pE:�y��RFЭ��NVh t $+MD�qIё)�v+�tń�tH�`�P�u�<|��sANSW}��t(�?�uD�)�r��	@Ði �@CU���V�T0'QoARR2�j Dɐ�Qނ~�Bd$CALI�@�F�G�s�2�RI�N��v�<��NTE���kE���,�V�����_Nl��ڂ���kDׄRm�DIVFiFDH�@ـn��$V��'c!$��$Z������~�[��oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS�@#2L�q�Ɣ83ಀ����� ��PAT!H��������3̒Vp�A_�Q�.�4�B��Cᐈ�_MGh��$DDQ���G�$FWh��p��m������b�DE��PPAB�NԗROTSPE!ED����00J�Я�8��@���$US�E_��P��s�S�Y��c�A kqYNru@Ag��OFF�qn�MOUN�NGg��K�OL�H�INC *��a��q��Bj�L@�BENCS��q'RđX���D��IN#"I(�0��4�\BݠVEO�w�>Ͳ23_UPE�߳/LOWL���00����D��'RwP���� �1RCʀƶMO3SIV�JRMO���@�GPERCH  �OV��^��i� <!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸUPp������TRKr�>"AYLOA'a��  Q-�(�<�1Ӣ`0 ���RTI$Qx�0 MO ���МB R�0J��D���s�H����b�DU�M2(�S_BCKLSH_C(���>� =�q�#�U��ԑ���2�<t�]ACLALvŲp�1n�P�CHK00:'%SD�RTY4�k���y�1�q_6#2�_�UM$Pj�Cw�_�S�CL��ƠLMT_OJ1_LO�'P���q��E�����๕�幘SPC��7���L���PCo���H� ȰPU�m�C/@�"XT\_�c�CN_��N��Le���SFu���V��&#����9�(���=�C�u�SH6#��c��� �1�Ѩ�o�0�͑
��f_�PAt�h�_Ps�W�_10��4�R�01D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�sR0Hљ��_W��-ԁ_=��C��I��I*�I�II�F�`�aJLA.�1[�VC��0�D�BO1U�@i�B\JRKU��~	@DBL_SMd�:BM%`_DLC�BGRV��C��I���H_� �*CcOS+\�(LN� 7+X>$C�9)I�9)u*c,)�Z2 HƺcMY@!�( "TH&-��)THET0�N�K23I��"=�A C-B6CB=�C�A�B�(261C�616SB8C�T25GTS QơC��aS$" �4c#<�7r#$DUD�EX��1s�t��B�6���AQ�|r�f$NE�DpI B U�\B5��$!��!�A�%E(G%(!LCPH$U�2׵�2SX pCc%pCr%�2�&�C�J�&!�VAHV6H3�YLUVhJVuKV�KV�KUV�KV�KV�IHAH@ZF`RXM��wXuKH�KUH�KH�KH�KH�I�O2LOAHO�YWNO�hJOuKO�KO�KO*�KO�KO�&F�2#1�ic%�d4GSPBA?LANCE_�!�c�LEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%�Ċ1ky�UTO_<?�jT1T2Cy��2N&�v�ϰctw�gѠp�0Ӓ~���T��O����� INSEGv�!�REV�v!���gDIF��1l�w6�1m�0OB�q
����MIϰ1��L�CHWAR����A�B&u�$MEC�H,1� :�@�U�AX�:�P��Y�G$�8pn� 
Z��|���RO�BR�CR��N�|&�MSK_�`�f�p P Np_���R����΄ݡ�1 ��ҰТ΀ϳ��΀"��IN�q�MTC�OM_C@j�q � L��p��$ONORE³5����$�r 8� GRl�E�SD�0ABF��$XYZ_DAx5A���DEBU�qXI��Q�s �`$�wCOD�� ���k�F�f�$BU�FINDXР � ��MOR��t $-�U��)��rРB��������Gؒu� � $SIMULT ��~�� ����OBJE�` �AD�JUS>�1�AY_	Ik��D_����C��_FIF�=�T � ��Ұ��{��p� ��З��p�@��D�FRiI��ӥT��RO� Ұ�E�{�͐OPsWO�ŀv0���SYSBU�@ʐ$�SOP����#�U<"��pPRUN�I�PA�DH�D����_OU�=��qn�{$}�IMAG��iˀ�0P�qIM��Ơ�IN�q���RGOVRDȡ:���|�aP~���Р�0L_6p0���i��RB���0e��M���EDѐ*F� ��N`M*���3x�̰SL�`ŀ�w x $OV�SL�vSDI��DEXm�g�e�9w�����V� ~�N���w�����Ûǖȳ�M��͐�q<��� x� HˁE�F�ATUS���C�0àǒN��BTM����If����4����(�ŀy DˀEz�g���P�E�r�����
���EXE��V��E�Y�$Ԝ� ŀz @ˁ��U�P{�h�$�p��X�N���9�H� ��PG"�{ h $SUB��c�@�_��01\�MPWAeI��P����LO���<�F�p�$RCVFAIL_C恎f�BWD"�F���D�EFSPup | Lˀ`�D�� U�UNI��S��ѱR`���_L�pP$����P�ā}��� @B�~���|��`ҲN�`�KET��y���Pԙ $�~���0SI�ZE�ଠ{���S�<�OR��FORMAT/p � F���r�EMR��y�UX8���@�PLI7�ā�  $�P�_SWI��Ş_�PL7�AL_ )�ސR�A��B�(0uC��Df�$Eh�[���C_=�U� � � ����~�J3�0����TWIA4��5��6��MOM������4 �B�AD��*���* PU70NR W��W ��V������ A$PI �6���	��) �4l�}69��Q���c�_SPEED�PGq� 7�D�>D�����>tMt[��SAM�`痰>��MOV���$��p�5���5�D�1�$2��������{�Hip�IN?,{�F( b+=$�H*�(_$�+�+�GAMM�f�1{��$GET��ĐH�D�����
^pLIBRt�ѝI��$HI��!_��Ȑ�B6E��*81A$>G086LW=e6 \<G9�686��R��ٰ�V��$PD#CK�Q�H�_����;"��z�.%�7��4*�9� ��$IM_SRO�D`�s"���H�"�LE��O�0\H��6@�bp��U� �ŀ�P�q?UR_SCR�ӚA�Z��S_SAVEc_D�E��NO��CgA�Ҷ��@�$��� �I��	�I� %Z[�  ��RX" ��m���" �q�'"�8�H ӱt�W�UpS��хDM��O㵐.'}q�� Cg���@ʣ�ߑ�R��M�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PL�M���	� 0h�H�{�X��O��z�Z�eT�M����� pS��C ��O__0_B_�a��_%�� |S����@ 	�v��v �@���w�v��EM��% v(R�fr�B�ː��ft�P��PM��QU.� �U�Q��A�f�QTH=�HOLޛ�QHYS�ES��,�UE��B��O.#��  -�P0�|��gAQ���ʠu���O��ŀ�ɂv�-�A;ӎ�ROG��a2�D�E�Âv�_�ĀZ�INFO&��+�����b�R�OI킍 =((@SLEQ/��#������o���DS`c0O�0�01�EZ0NUe�_�AUyT�Ab�COPY�P�Ѓ�{��@M��N������1�P�
� ��RiGI�����X_�P�l�$�����`�W��P��j@�G���EXT_CYCtb!���p����h�7_NA�!$�\��<�RO�`]�� � m��PORp�ㅣ���SRVt��)����DI �T_ l���Ѥ{�ۧ��ۧ Ъۧ5٩6٩7٩8����AS�B쐒���$�F6���PL8�A�A^�TAR��@ E `�Z�����<��d7� ,(@FLq`hѦ�@YNL���M�C���PWRЍ��=�e�DELAѰ��Y�pAD#qX� ��QSKIP�� iĕ�x�O�`NT!���P_x���� �@�b�p1�1�1� ��?� �?��>��>��&�>�3�>�9�Js2R;쐖 4��EX� TQ����ށ �Q���[�KFд�R�wRDCIf� �U`
�X}�R�#%M!*��0�)��$RGEAR�_0IO�TJBFL1G�igpERa��T�C݃������2TH�2N��� 1��b��Gq T�0 I����M���`Ib�\���REF�1�� l�h��ENA9B��lcTPE?@�� ��!(ᭀ����Q�#��~�+2 H�W���2�Қ���"�4�F�X�
j�3�қ{����(����j�4�Ҝ��
���.�@�R�j�5�ҝ�u�����������j�6�Ҟ��(:L
j�7�ҟo���(��j�8�Ҡ���"4Fj�SMS�K�����a��E��A��MOTE������@ "1�L�Q�IO�5"%I���P��POWi@쐣  �����X�gpi��쐤��Y"$DSB_SIGN4A�Qi��̰C���tRS23�2%�Sb�iDEVICEUS#�R�R�PARIT�!O�PBIT�Q��O?WCONTR��QXⱓ�RCU� M�S�UXTASK�3NxB��0�$TATU�PK�S@@쐦F��6�_�PC}�$F�REEFROMS8]p�ai�GETN@S��UPDl�ARB��S�P%0���� !>m$USA���a8z9�L�ERI�0f�&�pRY�5~"_�@f�qP�1�!�6WRK�D9�F9ХFR�IEND�Q4bUFx��&�A@TOOLHF�MY5�$LEN�GTH_VT��FCIR�pqC�@�E� �IUFIN�R����RGI�1�AITI:�xGX��I�FG2�7G1a����3��B�GPRR�DA��Oa_� o0e�I1RER�0đ�3&���TC���AQJV�G|�.2���F��1�!d�9Z�8 +5K�+5��E�y�L0�4��X �0m�L
N�T�3Hz��89��%��4�3G��W�0�W�RdD�Z��Tܳ���K�a3d��$cV �2���1��I1TH�02K2sk3K3Jci�aI�i�a�0L��SL��R$Vؠ�B�V�EVk�]V*R��� �,6Lc���9V2�F{/P:B��PS_�E���$rr�C�ѳ3$A0��wPR���v�U�cSk�� {���2���� 0���VX`�!�tX`��0P��ꁂ
�5SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V��� �S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD��<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C���:c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQkfC�ѷ =	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�qG �X��ȑ����$.A$�1$�c1Ó���� x~�EG�0ݓ��q!AR����09p>B�%��AXE���ROB��W�A4�_�-֣SY���!6��&MS�'WR���-1���STR��5�9�E�� 	5B��=QB90�@6������kOT�0o 	$�ARY8�w20����	%�FI��;�$�LINK�H��1��a_63�5�q�2XYZ"��;�q�3�@��1�2�8{0B�{D��� CFI��6G��
�{�_J��6��3a'OP_O4Y;5�Q#TBmA"�BC
�z��DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ ��@�5<:7�� +1�?0K�Mc�6�8Cb�vrb�4�ORQ��X�>8�#op�� ����wq�Uf�����T'OVE�Q��M;�@E#�UK#�UQ"�VW�Z Q�W���Tυ� ;� ���QH�!`�ҽ��U�Q��WkeK#kecXER��	GE	0��S�dAWaǢ:D���7!�!AX�rB! {q��1uy-!y �pz�@z�@z6Pz \Pz� z1v�y �y�+y�;y�Ky �[y�ky�{y��y��q�yDEBU��$����L�!º2WG`  AB!�,��S9V���� 
w��� m���w����1���1�� �A���A��6Q��\Q����!�m@��2CLAB3B�U�����So  ÐER��>�� � $�@� mAؑ!p�PO���Z�q0w�^�_MR}Aȑ� d  9T�-�ERR��TYz�B�I�V83@�cΑTOQ�d:`L� �d2�p ��˰�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	�SFZN�_CFG_!� 4 ��?º�|�ų����@�<ȲW iV ��\$� �n���Ѵ��09c�Q��(�FA�He�,�XEDM�(���H��!s�Q�g�P{R�V HELLĥ�� 56�B_BAS!�RSR��ԣo E�#S��[��1r�U%��2ݺ3ݺ4ݺU5ݺ6ݺ7ݺ8ݷ��ROOI䰝0�03NLK!�CAB� n��ACK��IN��T:�1�@�@ z�m�7_PU!�CO� ��OU��P� Ҧ) ���޶��TPFWD�_KARӑ��R�E~��P��(��Q�UE�����P
��C�STOPI_AL �����0&���㰑�0GSEMl�b�|�M��6d�TY|�SOK�}�DI�����(����_TM\�MANR�Q�ֿ0E+�|�$�KEYSWITCaH&	���HE
�OBEAT����E� �LEҒ���U��F�O�����O_HOuM�O�REF�P�PRz��!&0��Cr+�OA�ECO��xB�rIOCM�D8׵�]���8�` G� D�1����U���&�MH�»P�CFOsRC��� ���OM�  � @�V��|�U,3P� 1(-�`� 3-�4���NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F��V ��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��C@�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7sE&��VP��UPD�� � ��|�԰��YS�LOǢ� �  z��и���o�E��`>�8^t��АALUץ�����CU���wFOqIgD_L�ӿuHI�z�I�$FILE_����t��$`�JvS�A��� h���E_BLCK�#�C>,�D_CPU<�{� <�o����tJr���R ��
PWl O� ��LA���S��������RUN F�Ɂ��Ɂ����F�����ꁬ�M�TBC�u�C� �X ;-$�LENi���v������I��G�L�OW_AXI�F)1��t2X�M����hD�
 ��I�� ���}�TOR����Dh��� L=��⇒�8s���#�_MA`�8ޕ��ޑTCV����T���&��ݡ�����J�����J����MDo���J�Ǜ ����
���2��� v���l��F�JK��VKi�hΡv�Ρ3��J0㤶ңJJڣJJ�A�ALң�ڣ��42�5z�&�N1-�9�(��␅�L~�_Vj�x������ ` ��GROU�pD��B>�NFLIC��REQUIREa�EBUA��p����2¯�����c��� \��APP�R��C���
�E�N�CLOe��SC_M v�,ɣ�
�ޣ�� ���MCp�&���g�_MG�q�C� �{�9���|�wBRKz�NOL��t|ĉ R��_LI|�H�Ǫ�k�J����P
� ��ڣ�����&���/�"��6��6��8���|���� ���8�%�W�2�e�PATHa�z�p�z�=�vӴ��ϰ�x�CN=�CaA�����p�IN��UC��bq��CO�U�M��YZ������qE�%���2������PA�YLOA��J2L�3pR_AN��<�L���F�B�6�R�{�R_?F2LSHR��|�LOG��р��ӎ���ACRL_u��������.���H�p�$yH{���FLEX
���J�� :�/����6�2�`����;�M�_�F16� ����n���������ȟ��Eҟ�����,� >�P�b���d�{�������������5�T��X��v���E ťmFѯ����� ��&�/�A�S�e�D�}Jx�� � ��0����j�4pAT����6n�EL  �%ø�J���ʰJE��C�TR�Ѭ�TN��F�&��HAND_V�B[
�pK�� $F2{�6� �r�SW$#s�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�+p�K�� &0�_��ER!V9�SQASYM$��] �����x�������_SHl����� ��sT�(����(�:�JA���S�cir��_VI�#Oh9�``V_UNI��td�~�J���b�E�b��d ��d�f��n�������H��uN���D�2�H������"Cq3EN� a�DI��>�Obtas�Dpx�S� ��2IxQA�� ��q��-��s �� s�ܒ��� ��OMME��rr/�TVpPT�P ���qe�i����P�x ��y�T�Pj� $D�UMMY9�$7PS_��RFq�0;$:� s����!~q� X����K��STs�ʰSBR���M21_Vt�8�$SV_ERt�O���z���CLRx�A�  O�r?p? Oր �� D $GgLOB���#LO�ЀՅ$�o��P�!S;YSADR�!?p��pTCHM0 �� ,����W_NA��/�e���Q�SR��l (:]8:m�K6�^2 m�i7m�w9m��9���� ���ǳ���ŕߝ�9ŕ ���i�L���m���_�_�_�TtqXSCSRE�ƀ�� ��3STF���}�pТR6�sq] _v AŁ�� T����TYP �r�K��u�!u����O�@IS�!���tC�UE{t� �����H�S���!R�SM_�XuUNE�XCEPWv��CpS_��{ᦵ�ӕ���÷���COU ���o 1�O�UET��փr���PROG�M� FLn!$C�U��PO*q��c�I�_�pH;� � �8��N�_HE
p���Q��pRY ?A���,�J�*��;��OUS�� � �@d���$BUT�T��R@���COL�UM�íu�SERyVc#=�PANEv �Ł� � �PG�EU�!�F��9�)�$HELP��WRETER��)״�� �Q������@�0 P�P �IN��sE�PNߠw v�1�y���� ���;LN�� ����9_��k�$H��M �TEX�#����FLyAn +RELV��D4p�������M��?,��ӛ$�����P=�USRVI;EWŁ� <d��puU�p0NFIn �i�FOCU��i�PRI# m+�q���TRIP)�m�sUNjp{t� QP<��XuWARNWud�_SRTOLS�ݕ������O|SORNN��RAUư��T���%��VI|�zu�� $�PATyHg��CACH�LOG6�O�LIM�ybM���'��"�HO;ST6�!�r1�=R�OBOT5���KIMl� D�C� g!���E�L���i�VC�PU_AVAIL�B�O�EX7�!BQN L�(���A�� Q��Q� ��ƀ�  �QpC���@$T�OOL6�$�_J;MP� �I�u�$SS�!$sqV�SHIF��|s�AP�p�6�s���R�^��OSURW�p�RADIz��2�_ �q�h�g! �q)��LUza$OUT?PUT_BM��IML�oR6(`)�@wTIL<SCO�@Ce�;��9��F ��T��a��o�>��3�����w�2u�.�PV�zu��%�D�JU��|#�WA�IT������%�ONE��YBO�ư �� �$@p%�C�SBn)T;PE��NEC��x"p�$t$���*B_T��R��%�qR� ���s	B�%�tM�+��t�.`�F�R!݀��OPm�wMAS�_DOG�OaT	�D����C3�S�	�O2DELAY���e2JO��n8E� �Ss4'#J�aP6%�����Y_��O2$��2����5��`? ��ZABCS�� � $�2��J�
�b��$$CLAS>�����AB�xb�'@@VIRT��O.@ABS�$�1� <E� < *A tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R��d�v�����M@[�AXmLր ���dC7  ���IN��ā���PRE������LARMRE?COV <I䂶��NG�� \K	? A   J�\��M@PPLIC�?�<E�E��Handling�Tool �� �
V7.50P/�28[�  �H����
�_SW UP*A� F��F0ڑ����A@~�� 20���*A���:�����FB 7wDA5�� #'@?I�@���None������� ��T��~*A49�xl�E_��V����g�UTOB�ค����?HGAPON8@���LA��U��D 1<EfA����������� Q 1"שI Ԁ��Ԑ��:�i�n����#B{)B ����\�HE�Z�r�HTTHKY��$BI� [�m�����	�c�-� ?�Q�o�uχϙϫϽ� �������_�)�;�M� k�q߃ߕߧ߹����� ���[�%�7�I�g�m� ������������ W�!�3�E�c�i�{��� ������������S /A_ew��� ����O+= [as����� ��K//'/9/W/]/ o/�/�/�/�/�/�/�/ G??#?5?S?Y?k?}? �?�?�?�?�?�?COO O1OOOUOgOyO�O�O �O�O�O�O?_	__-_0K_Q_��(�TO4�s����DO_CLEA�N��e��SNM  9� �9oKo�]ooo�o�DSPDgRYR�_%�HI��m@&o�o�o#5 GYk}����0"���p�Ն �ǣ��qXՄ��ߢ��g�PLUGGҠ�Wߣ��WPRC�`B`9��o�=�OB��oe�/SEGF��K���� ��o%o����#�5�m���LAP�oݎ�� ��������џ������+�=�O�a���TO�TAL�.���USWENUʀ׫ �X����R(�RG_STRING 1���
�M��S�c�
��_ITE;M1 �  nc�� .�@�R�d�v������� ��п�����*�<��N�`�r�I/O SIGNAL���Tryout� Mode�I�np��Simul�ated�Ou�t��OVER�R�` = 100��In cyc�l���Prog� Abor���~��Status��	Heartbe�at��MH F�aulB�K�AlerUم�s߅ߗߩ߻����������  �S���Q��f�x�� ������������� ,�>�P�b�t�������,�WOR������V� ��
.@Rdv ��������*<N`PO ��6ц��o��� ��//'/9/K/]/ o/�/�/�/�/�/�/�/�/�DEV�*0� ?Q?c?u?�?�?�?�? �?�?�?OO)O;OMO�_OqO�O�O�OPALTB��A���O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o:o�OGRI�p��ra �OLo�o�o�o�o�o�o *<N`r�������`o��R B���o�>�P�b�t� ��������Ώ���� �(�:�L�^�p����PREG�N��.��� �����*�<�N�`� r���������̯ޯ����&����$AR�G_��D ?	����i���  	$���	[}�]}����Ǟ�\�SBN_C�ONFIG �i�������CI�I_SAVE  ���۱Ҳ\�TC�ELLSETUP� i�%HO�ME_IO�͈�%MOV_�2�8��REP���V�UT�OBACK
��ƽFRA:\�� �Ϩ���'` ��������� ����$�6��c�Z�lߙ��Ĉ�� �����������!凞 ��M�_�q����2� ��������%�7��� [�m��������@��������!3E$���Jo��������INI�@���ε��MESSA�G����q��OD�E_D$���Ox,0.��PAUS��!�i� ((Ol������� � /�//$/Z/H/�~/l/�/�'akTSK  q������UPDT%�d�0;WSM_CF°i�еU�'1�GRP 2h�93� |�B��A�/S�XoSCRD+11
1;' ����/�? �?�? OO$O��߳? lO~O�O�O�O�O1O�O UO_ _2_D_V_h_�O�	_X���GROUN�0O�SUP_NA�L�h�	�ĠV_�ED� 11;
 ��%-BCKEDT-�_`�!oEo$����a��o������ߨ���e2 no_˔o�o�b���eep�o"�o�oED3 �o�o ~[�5GED4�n#�� ~p�j���ED5Z� �Ǐ6� ~���}���ED6����k�ڏ ~pG���!�3�ED7�� Z��~� ~�V�şן�ED8F�&o��Ů�}����i�{�ED!9ꯢ�W�Ư
}3�����CRo���� �3�տ@ϯ����P�P?NO_DEL�_�R�GE_UNUSE��_�TLAL_OU�T q�c�QW?D_ABOR� ����Q��ITR_RT�N����NONS�e���CAM�_PARAM 1��U3
 8
�SONY XC-�56 23456�7890�H �� @���?�>��( АV�|[�r؀~�X�HR�5k�|U�Q�߿�R5y7����Aff���KOWA SC�310M|[r��>��d @6�|V ��_�Xϸ���V���  ���$�6��Z�l���CE_RIA_I�857�F�1���R|]��_LeIO4W=� ��P�<~�F<�GP 1.�,���_GxYk*C*  �V�C1� 9� @� iG� �CLC]� Ud� l� s�R� T��[�m� v� �� �� �� C�� �"�|W��7�{HEӰONFI� ���<G_PRI 1�+P�m®/���������'C�HKPAUS�  ;1E� ,�>/ P/:/t/^/�/�/�/�/ �/�/�/?(??L?6?h\?�?"O������H�1_MOR��� �XaBiq-<���5 	 �9 O �?$OOHOZK�2	���=9"�Q?55���C�PK�D3P��|����a�-4�O__|Z
�OG_�7@�PO�� ��6_��,xV��ADB���='�)�
mc:cpmi�dbg�_`��S:�"(�����Up�_)o��S  �3Pq����R�P�_mo8j�����Oko�oV9i�(�=(�>Ok�g�o�o�l�Kof��oGq:I�ZDEFg f8��)�R�6pbuf.txt m�]n�@����# �	`(Ж�A=L�m��zMC�21�=�a� :���4�=��n׾�Cz  BH�BCCPUeB��_B�y;���>C���Cn�aSWE@E?{hD�]^Dْ?�r����D��^���G	��F���F��Cm	�fF�O�F��I�SY���vqG����Em�(�.����1(��<�q�G�x�2��Ң �� a�D��j���ES\��X��EQ�EJ�P F�E�F�� G���F�^F E�� F�B� H,- Ge��H3Y�����`�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE ��O@b 
�(�;��"�  <�6�z�Rb���?�j�C4�(�aSWm� W��{�Jm�C��B-G�Cu��@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"��_ , 
�^����o xvf`MT�I�^�rl@�:sONT�IM�������Zv�i
õ�cMOT�NEND���dRECORD 1(R�qa��ua�O��q ��sb�.�@�R��x Z�������ɏۏ� ����#���G���k�}� ����<�ş4��X�� �1�C���g�֟���� ����ӯ�T�	�x�-� ��Q�c�u�������� ��>����)Ϙ�M� ��F�࿕ϧϹ���:� ������%�s`Pn&�]� o��ϓ�~ߌ���8�J� ����5� ��k��� �ߡ��J�����X�� |��C�U�������� ���0�����	��db�TOLERENC�qdBȺb`L����PCS_CFG �)�k)wdM�C:\O L%04�d.CSV
�`cl�)sA �CH� z�`)~���h�MRC_OUT �*�[�nSG�N +�e�r���#�10-MAY�-20 10:4�6*V15-JAN�j51�k P/Vt��)~�`�pa�m��P�JPѬVE�RSION �SV2.0.�8.|EFLOGI�C 1,�[ 	DX�P7)�PF."�PROG_ENB��o�rj ULSew ��T�"_WRST�JNEp�V�r`dEM�O_OPT_SL� ?	�es
 ?	R575)s7)��/??*?<?'�$TO  �-��?&[V_@pEX�Wd�u��3PATH ASA\�?�?O�/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C��SqqF�PMAU�� t/XrMSWR.D�i�a.|S/�Z!D_N�O0__T_C_�x_g_�_�tSBL_/FAUL"0�[3w/TDIAU 16M�a�p�A12�34567890gFP?BoTofo xo�o�o�o�o�o�o�o ,>Pb�S�p-P�_ ���_s �� 0`����� )�;�M�_�q����������ˏݏ��|)UM�P�!� �^�T�R�B�#+�=�PME�fEI�Y_TEMP9 È�3@�3A �v�UNI�.(YN_BRK 2Y�)EMGDI_S�TA�%WЕNC2_SCR 3��1o"�4�F�X�fv����������#��ޑ14����)�;���t��ݤ5��� ��x�f	u�ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /߭P�b�t�� ��x� �߰���������
�� .�@�R�d�v���� ����������*�<� N���r����������� ����&8J\ n������� �"`�FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/4?,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O? �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �o�O�O�o�o�o
 .@Rdv��� ������*�<� N�`�r����o����̏ ޏ����&�8�J�\� n���������ȟڟ�����H�ETMODoE 16���W ��ƨ
R��d�v�נRROR_PROG %A��%�:߽�  ��TABLE  A�������#�L�RR�SEV_NUM � ��Q���K�S���_AUTO_ENB  ���I�Ϥ_NOh� �7A�{�R�  �*������������^�+��Ŀֿ迄��HISO�͡I�}�_�ALM 18A�� �;�����+ �e�wωϛϭϿ��_H���  A��|��4�TCP_�VER !A�!�����$EXTLO�G_REQ��{�V�SIZ_�Q�T�OL  ͡Dz���A Q�_B�WD����r���n�_�DI�� 9���}�z�͡m���ST�EP����4��OP�_DO���ѠF�ACTORY_T�UN�dG�EAT?URE :�����l�Han�dlingToo�l ��  - C�Englis�h Dictio�nary��ORD�EAA Vi�s�� Masteyr���96 H���nalog I/yO���H551���uto Soft�ware Upd_ate  ��J���matic Ba�ckup��Par�t&�ground Edit���  8\ap�Camera��F���t\j6R�elyl���LOADR�7omm��shq��oTI" ��co��
! o���p�ane�� 
!���tyle s�elect��H5�9��nD���oni7tor��48�����tr��Relia�b���adin�Diagnos�"����2�2 ual� Check S�afety UI�F lg\a��h�anced Ro�b Serv q� ct\��lUs�er FrU��D�IF��Ext. oDIO ��fiAs d��endr �Err L@��I%F�r��  �П��90��FCTN /MenuZ v'���74� TP In���fac  S�U (G=�p���k Excn g��3��High-wSper Ski+�  sO�H9 � m�munic!�on5sg�teur� �����V����c�onn��2��ENމ�Incrst�ru���5.fd�KAREL �Cmd. L?u�aA� O�Runw-Ti� Env��R��K� ��+%�s#�S/W��74��L?icenseT��  (Au* ogBook(Sy���m)��"
MACROs,V�/Offse��a�p��MH� ����p�fa5�MechS�top ProtL��� d�b i��Shif���j545�!xr ��#���,K�b ode Switch��m\e�!o4.�& pro�4���g��Multi�-T7G��net�.Pos RGegi��z�P���t Fun���3s Rz1��Numx ������9m�1�  �Adjuj��1 J7�7�* ����6�tatuq1EIK�RDMtot���scove�� ���@By- }uest1�$Go� � U5�\SNPX �b"���YA�"Li�br����#�� �$~@h�pd]0�J�ts in VCCCM�����0�  �u!��2 R�0�/�I�08��TMI�LIB�M J92:�@P�Acc>�F�{97�TPTX�+6�BRSQelZ0�M�8 Rm��q%��6�92��Unexc�eptr motn>T  CVV�P���KC����+-��~K  II)�VS�P CSXC�&.ac�� e�"�� t�@�Wew�AD� Q�8bvr nm�en�@�iP� a�0y�0�pfGri�dAplay !�� nh�@*�3R�1M-�10iA(B20k1 �`2V"  F����scii�lo{ad��83 M��yl����Guar�dO J85�0�mP'��L`���stuaPa9t�&]$Cyc����|0ori_ x%Da�ta'Pqu���cAh�1��g`� j� RLJam�5���IMI De-B(�\A�cP" #^0C~  etkc^0�asswo%q�)6�50�ApU�Xn�t��Pven�CT�qH�5�0YELLOW BO?Y���� Arc�0vi�s��Ch�Wel=dQcial4Izt�Op� ��gs�`k 2@�a��poG3 yRjT1 NEf�#HT� xyWbF��! �p�`gd`����p\� =P��JP�N ARCP*P�R�A�� OL��pSup̂fil��p��J�� ��cro�670�1C~E�d���SS�pe�tex��$ �P� So7 t^� ssagN5 <Q"�BP:� �9 "0�Q#rtQC��P�l0dpn�笔�rpf�q��e�ppmas�cbin4psy=n�' ptx]08��HELNCL �VIS PKGS9 �Z@MB &���B J8@IPE� GET_VAR� FI?S (Un�i� LU�OOL:� ADD�@29.KFD�TCm���E�@�DVp���`A�ТN�O WTWTEST �� V�!��c��FOR ��ECT� �a!� ALSE� ALA`�CPMO-130��� b �D: HANG FROMg��2���R709 DRA�M AVAILC�HECKS 54�9��m�VPCS �SU֐LIMCH�K��P�0x�FF WPOS� F�� q�8-12 C�HARS�ER6�O�GRA ��Z@AV�EH�AME��.SV��Вאn$��9�wm "y�TRCv�� SHADP�UP�DAT k�0��S�TATI��� M�UCH ���TI�MQ MOTN-�003��@OB�OGUIDE DAUGH���b��@�$tou� �@C� <�0��PATH�_��MOVET�� R�64��VMXPA�CK MAY A�SSERTjS��C�YCL`�TA��B�E COR 71��1-�AN��RC �OPTIONS � �`��APSH-�1�`fix��2�S�O��B��XO򝡞�_�T��	�i��0j��d�u�byz p wa��y�٠HI�������U�pb XSPD �TB/�F� \hcehΤB0���END�[CE�06\Q�p{ }smay n@��pk��L ��tr'aff#�	� ���~1from sy�svar scr��0R� ��d�DJUD���H�!A��/��SET ERR��D�P7����NDA�NT SCREE�N UNREA �VM �PD�D��P�A���R�IO gJNN�0�FI��}B��GROUNנD Y�Т٠�h�SVIP 53 Q�S��DIGIT �VERS��ká�N{EW�� P06�@=C�1IMAG�ͱ4���8� DI`����pSSUE�5��EPLAN JON�� DEL���157�QאD��CALL�I���Q��m���IP�ND}�IMG N�9 PZ�19��MwNT/��ES ���`LocR Hol�߀=��2�Pn� PG�:��=�M��can�����С: 3D� mE2view gd X��ea1 ��0b�pof Ǡ"�HCɰ�ANNO�T ACCESS? M cpie$E�t.Qs a� lo^MdFlex)a:���w$qmo G�sA�9�-'p~0��h0pa���eJ AUTO1-�0��!ipu@Т|<ᡠIABLE+�� 7�a FPLN:9 L�pl m� �MD<�VI�и�W�IT HOC�Jo~1Qui��"���N��USB�@�Pt� & remov����D�vAxis �FT_7�PGɰC�P:�OS-14�4 � h s 2968QՐOST�p � CRASH D�U��$P��WOR�D.$�LOGI�N�P��P:	�0�0�46 issue�E�H�: Slo[w st�c�`�6����໰IF�I�MPR��SPOT�:Wh4���N1STyY��0VMGR�\b�N�CAT��4oR�RE�� � 5�8�1��:%�RTU�!Pe -M a�SE:B�@pp���AGpL��r�m@all���*0a�OCB WA����"3 CNT0� T9DWroO0a�larm�ˀm0d� t�M�"0�2|� 9o�Z@OME<�� ���E%  #1-�S�RE��M�st}0g�     5K�ANJI5no �MNS@�INISITALIZ'�3 E�f�we��6@�� dr�@ fp �"��SCII L��afails w|��SYSTE[��i��  � Mq��1QGro8�m �n�@vA����&��nx�0q��RWRI �OF Lk��� \gref"�
�up� de-rela�Q_d 03.�0SS�chőbetwe�4�IND ex 6ɰTPa�DO� �l� �ɰGigE��soperabi]l`p l,��Hc�B��@]�le�Q0c�flxz�Ð���O�S {����v4pfigi GLA�$�c2z�7H� lap�0�ASB� If��g�2 l\c�0��/�E�� EXCE	 㰁�P���i��� o0��Gd`]Ц�f<q�l lxt��EFal��#0�i�O�Y�n�CLOS��S[RNq1NT^�F��U��FqKP�ANIO' V7/ॠ1�{����DB �0���v��ED��DET|��'� �bF�NLI;NEb�BUG�T�:��C"RLIB��A���ABC JAR�KY@��� rkeMy�`IL���PR���N��ITGAR� D$�R �Er *�T��a�U�0��h�[��ZE V� TASK p.vr��P2" .�XfJ�srqn�S谥dIBP	c����B/��BUS.��UNN� j0-��{��cR'���LO�E�DIVS�CUL`s$cb����BW!���R~�W`P�����I�T(঱tʠ�OF��UNEXڠ+����p�FtE��SVE�MG3`NML 5�05� D*�CC_SAFE�P*� ���� PET��'P�`��F  !���IR(����c i S>� �K��K�H GU�NCHG��S�M�ECH��M��T�*�%p6u��tPOR�Y LEAK�J���SPEgD��2�V 74\GRI���Q�g��CTLN��TRe @�_�p ��6�EN'�IN���`���$���r��T3)�.i�STO�A�s�	L��͐X	���q��1Y� ��TO2�J �m��0F<�K����D)U�S��O��3	 9�J F�&���S?SVGN-1#I�N��RSRwQDAU�C@ޱ� �T6�g��� 3��]���BRKCTR8/"� �q\j5��_��Q�S�qINVJ0D ZO�Pݲ���s���г�Ui ɰ̒�a�D�UAL� J50�e�x�RVO117 AW�TH!Hr%�nN�247%�52��|�&aol ���R��(�at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���M�d�Rǰt� \fosB�A�0Np�c�����{�U��ROP �2�b�pB��ITP�4M��b !AU�t c0< � plet9e�N@� z1^q�R635 (Ac�cuCal2kA���I) "�ǰ�1
a\�Ps��ǐ� b���0P򶲊���ig�\cbacul "A3p_ �1��ն����etaca��AT���PC�`�����;_p�.pc!Ɗ�<�:�circB����5�tl��Bɵ�:�f!m+�Ί�V�b�ɦ�~r�upfrm.����ⴊ�xed��Ί�N~�pedA�D �}b>�ptlibB�� �_�rt��	Ċ�a_\׊ۊ�6�fm�� ��oޢ�e��̆Ϙ���c�Ӳ�5�j>�����#tcȐ��	�r���ʸ�mm 1��T�sl�^0��T�mѡ�#�r�m3��ub Y�q�s3td}��pl;�&�cckv�=�r�vf������9�vi����Cul�`�0fp�q ��.f��� daq�; i Data A�cquisi��nB�
��T`��1��89��22 D�MCM RRS2�Z�75��9 3 �R710�o59�p5\?��T "��1 (D�T� nk@��������E Ƒ�ȵ��Ӹ�etdm�m ��ER����gxE��1�q\mo? ۳�=(G���[0(

�2�` ! �@�JMACRO��S�kip/Offs�e:�a��V�4o9<� &qR662����s�H�
 6Bq8�����9Z�43 �J77� 6�J783�o ��n�"vv�R5IKCBq?2 PTLC�Z�g R�3 (�s�, �������0�3�	зJԷ\sf�mnmc "MN�MC����ҹ�%mnf�FMC"Ѻ0�>� etmcr� ��8���� ,�K�DV� �  874\p'rdq>,jF0�ޢ�axisHPr�ocess Axwes e�rol^�PRA
�Dp� 56o J81j�59� 56o6� ���0w��690 98� [!I#DV�1��2(x2��2ont�0�
�����m2���?C��e�tis "ISD���9�� Fprax�RAM�P� D��d�efB�,�G�is_basicHB�@p޲{6�� 708�6��(�Acw:�������D
�/,��AMOX �� ��DvE��?;T��2>Pi� RAFM';�]�!PAM�V�W�Ee`�U�Q'
bU�75��.�ceNe� nt?erface^�1' 5&!54�K��b(Devam±�/�#����/<�Tane`"�DNEWE���btp_dnui �AI�_�s2�d_rsono���bAsfjN��bdv_arFvf�x0hpz�}w��hkH9x�stc��gApon1lGzv{�ff� �r���z�3{q'�Td>pchamp�r;e�p� ^597@7��	܀�4}0��mɁ��/�����lf�!�pcochmp]aMP&xB�� �mpev��8����pcs��Ye�S�� Macro�OD��16Q!)*��:$�2U"_,��Y�(PC ��$_;�������o��J�gegemQ@GEMSW�~ZG�gesndy��OD��ndda��S��s1yT�Kɓ�su^Ҋ�ĩ�n�m���L��  ���9:p'ѳ޲���spotplusp���`-�W�l�J��s��t[�׷p�key�ɰ�$��s�-Ѩ��m���\featu� 0FEAWD�o;olo�srn'!�2 p���a�As3��t�T.� (N. A.)��!e!�J#
 (j�,��oBIB��oD -�.�n��k9�"K��u[-�_����p� "PSE�qW����wop "sEЅ�&�:�J��� ���y�|��O8��5� �Rɺ���ɰ[��X� ������%�(
ҭ�q HL�0k�
�z�@a!�B�Q�"(g� Q�����]�'�.��� ��&���<�!ҝ_�#��tpJ�H�~Z��j��� ��y������2��e� �����Z����V��! %���=�]�͂��^2�@�iRV� on�Q$Yq͋JF0� 8ހ�`�	(^�dQueue���X\1�ʖ`�+~F1tpvtsn��YN&��ftpJ0v �RDV�	f��J1 iQ���v�en�^�kvstk��mp���btkclrq8���get�����r��`kacqk�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�m	c�N+v3�_� �����.v�/\jF��� �`Q�΋�ܒ�N50 (FR�A��+��͢fraparm��Ҁ�} =6�J643p:V��ELSE
#�V�AR $SGSY�SCFG.$�`_UNITS 2�D`G~°@�4Jgfr��4A�@FRL-��0ͅ �3ې���L�0NE�: �=�?@�8�v�9~Q�x304��;�BPR�SM~QA�5TX.�$VNUM_OLp��5��DJ507��~l� Functʂ�"qwAP��琉�3 �H�ƞ�kP9jQ�Q5 ձ� ��@jLJzBJ[ �6N�kAP����S>��"TPPR��\�QA�prnaSV��ZS��AS8Dj510U�-�`cr�`8 ���ʇ�DJR`jYȑH_  �Q �P�J6�a21��48�AAVM 5̕Q�b0 lB�`TU�P xbJ54s5 `b�`616����0VCAM ~9�CLIO b71�5 ���`gMSC8�
rP R`�\sSTYL� MNIN�`J6�28Q  �`NR�Ed�;@�`SCH ���9pDCSU M�ete�`ORSR� Ԃ�a04 kR�EIOC �a5.�`542�b9vpP@<�nP�a�`�R�`7�`��MASK 3Ho�.r7 �2�`OOCO :��r3� �p�b�p���r0X��a��`13\mn�a3?9 HRM"�q�q~��LCHK�u�OPLG B��a0�3 �q.�pHCR� Ob�pCpPosyi�`fP6 is[r�J554�òpDS�W�bM�D�pqR�a337 }Rjr0 �1�s�4 �R6�7��52�r5 �2�r7 1� P6���Regi��@T�uFRD�M�uSaq%�4�`9{30�uSNBA�u�SHLB̀\sf�"pM�NPI�S�PVC�J520v��TC�`"MNрoTMIL�IFV��PAC W�pTP�TXp6.%�TELN N Me��09m3UEC9K�b�`UFR�`���VCOR��VIPuLpq89qSXC�S��`VVF�J�TPy �q��R626l��u S�`Gސ�2�IGUI�C��P�GSt�\ŀH86�3�S�q�����q34:sŁ684���a��@b>�3 :B��1� T��96 .�+�E�51 y�q53̀3�b1 ���b1 �n�jr9 ���`VAsT ߲�q75 s�xF��`�sAWSMӞ�`TOP u�ŀRq52p���a80 
��ށXY q���0 \,b�`885�QXр�OLp}�"pE࠱t�p�`LCMD��EgTSS���6 �>V�CPE oZ1�gVRCd3
�NLH�h��001m2Ep���3 f��p��4 //165C��6l����7PR��008 �tB��9 -200��`U0�pF�1޲1	 ��޲2L"���p���޲4��5 \h�mp޲6 RBCF`�`ళ�fs�8 ������~�J�7 rbcfA�L�8\PC����"�32m0u�n�K��Rٰn�5 5EW�
n�9 z��4�0 kB��3 ��6|ݲ�`00iB/��I6�u��7�u��8 �0�������sU0�`�t� �1 05\rb��2 E���K���dj���5˰��60��a�HУ`:�63�jAF�_���F�7 ڱ݀H�a8�eHЋ��cU0���7�p��1u��8<u��9 73����&��D7� ��5t�W97 ��8U�1���2��1�1:���h���1np�"��8(�U=1��\pyl��,�p��v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6C B���цp��1��r��1�`͵155ض�157 �2��62 �S����1b��2$����1Π"�2����B6`�1<c�4� 7B�5 DR��8�_�B/��187 �uJ�8 06�9s0 rBn�1 (���202 0EW,�ѱ2^��2��90�U12�p�2��2 b��u4��2�a"RB����9\�U2�`w�l����4 60Mp��7�������b�s
5 ¿�3����pB"9 �3 ����`ڰR,:7 �2��V�2���5���2^��a^9����qr����n�5 ����5᥁"�8a�Ɂ}�5B���5����`!UA���� ��86 �+6 S�0��5�p�2<�#�529 �2^��b1P�5~�2�`���&P5��8"��5��u�!�5��ٵW544��5��R��P nB^z�c (4�����U5J�V�5��1�1^���%�����5 b2a1��gA��58W[82� rb��5N��E�5890r� 1�95 �"������ c8"a��|�L ���!�J"5|6��^!�6��B�"8�`#��+�58%�6B�AME�"�1 iC��622D�Bu�6V��d� 4��{84�`ANRSP�e/S� C�5 � �6� ��� \� �6�� �V� 3t��� �T20CA�R��8�� Hf� 1DH�� A�OE� �� ,K|�� �0\�� �!64K��ԓrA� ��1 (M-7�!/50T�[PM��P�Th:1�C�#Pe� ��3�0� 5`M75cT"� �D8p� �0�Gc� u�4��i1-7'10i�1� Skd�7�j�?6�:-HS, � �RN�@�UB�f<�X�=m75sA*A�6an���!/CB�B2.6A �0;A�CIB�A��2�QF1�UB2�21� /70�S� �4��A��Aj1�3p���8r#0 B2\m*A@�C��;bi"i1K�u"A�~AAU� imm7c�7��ZA@I�@�Df��A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5�*A�EA�5B�4>\77
B7=Q�D�2�Q$BR�E7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E
"l7�@7�A
1�E�V$~`�W2%Q�R9ї@0L_�#����"Aȉ��b��H3s=rA/2�R5nR4�74rNUpQ1ZU�A�s\m9
1M92L2�!F!^Y�ps� 2ci��-?�qhimQ�t  w043�C��p2�mQ�r�H_ �H2�0�Evr�QHsXBSt62�q`s����� �<�Pxq350_*A3#I)�2�d�u0�@� �'4TX�0�pa3i1A3sQ25�c��st�r�VR1%e�q0
��j1��O2  �A�UEiy�.�‐ �0dCh20$CXB79#A��ᓄM Q1]�~�� 9�Q��?PQ��qA!P vs� 5	15aU����?PŅ���ဝQ9A6�zS*�7�qb5�1p����Q��00P(��V7]u�aitE1���À�p?7� !?�z��r=bUQRB1PM=�Q�a9��H��QQ�25L��������Q��@L���8ܰ��y00\}ry�"R2BL�t�N  ��� �1DV��2�qeR�5���_b�3�X^]1m1lcqP1�a��E�Q� 5F����!5<���@M-16Q��  f���r��Q�e� ��8� PN�LT_�1��i1��9453��@�e�|�b1l>F1u *AY2�
��R8�Q����RJ�J3�D}T� 85
Qg�/0��*A!P@�*A�Ð𫿽�2ǿپ6t�6=Q���P�ȓ��� AQ�  g�*ASt]1^u�ajrI� B����~�|I�b��y&I�\m�Qb�I�uz��A�c3Apa9q� B6�S��S��m���}�8�5`N�N�  �(M���f1���6�����161��5�s`�SC��U��A�����5\set06c�����10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��� �5�B��B��h`�F� ��X0���A:���C�M�B��AZ��@��4�6i� ���� e�O�-	�� �f1��F �ᱦ�1pF�Y	���T6HL3���U66~`���U�dU�9D20Lf0��Qv � ��fjq��N���� ��0v
� ��i	�	.��72lqQ2�������� \chng�move.V��d����@2l_ar f	�f~��6��� ���9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�A]�,�V�1\�Qn�BJ�2W�EM!5�0��)�#:�64��F��e50S�\��0� =�PV���e�������E�����m7;shqQSH"U��)@��9�!A��(����� ,K��ॲTR1!��,�60e=�4F�����2��	 R-����� ������Ж��4���LSR�)"�!l�OA��Q�) %!� 16�
U/��2�"2��E�9p���2X� SA�/i��'�
7F�H �@!B�0��D���5V ��@2cVE��p��T�2�pt갖�1L~E�#ȚF�Q��9E�#De/��RT��59���	�A��EiR������9\7m20�20��+�-u�19r4�`�E1�= `O9`�1"ae��O2��_$W}am4�1�4�3�/d1c_std��1)�!�`_T��r�_ 4\jdg�a�q�PJ%! ~`-�r�+bgB��#Nc300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W�"Ps A��e���� t�i�P�W.��c�@FX.�e�kE14��44�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2a���2A;_2��QW2��bF�(�V11�23`�`��X5�Ra21�!J*9�a:88J99X�l5�m1a첚��*���(85�&��� ����P6���R,!52&A����,fA9INfI50\u�z�OV
 �v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&� �P1��vB)e�m������1p� �1D�V��27�F�KA�REL Use =S��FCTN��� J97�FA+�� (�Q޵�p%�)?�V�j9F?(�j�Rtk?208 "Km�6Q��y�j��iæPr�9��s#��v�krcfp�RCFt3���Q�¿kcctme�!M�E�g����6�mai�n�dV�� ��ru��kDº�c���o��L��J�dt�F ����.vrT�f������E%�!��5�FRj7%3B�K���UER�H�J�O  J�� (ڳF���F�q�Y�&T���p�F�z��19�tk vBr���V�h�9p�E�y�<�k������;�v���"CT��f�� ��)�
І��)�V	� 6���!��qFF��1 q���=�����O�?�$"����$��je���T?CP Aut�r�<�520 H5�J[53E193��9��+96�!8��9��	 n�B574��52�uJe�(�� Se%!�Y�����u��ma�Pqtool�ԕ��������conrel��Ftrol Re?liable�Rmv9CU!��H51���p�� a551e"<�CNRE¹�I�c�&��it�l\�sfutst "�UTա��"X�\u@��g@�i�6Q]V0�B$,Eѝ6A� �Q� )C���X��Yf�I�1�|6s@6i��T6AIU��vR�d�
$e%1��2�C58�E6���8�Pv�iV4OFH58�SOeJ� mvBM6E~O58�I�0�E�#+@ �&�F�0���F�P6a����)/++�</N)0�\tr1�����P �,K�ɶ�rmaski�msk�aA���Iky'd�h	A	�P�s�DisplayI�m�`v����J88G7 ("A��+Heůצprds��IϩǪ��h�0pl�2�R2Ƚ�:�Gt�@��PRD�TɈ�r�C�@Fm�8�D�Q�AscaҦ�� V<Q&��bVvbrl�eې@��^S��&5�Uf�j8710�yAl	��Uq���7�&��p�p��P^@�P�firmQ����Pp�2�=bk�6�r�3��6��otppl��PL���O�p<b�ac�q	��g 1J�U�d�J��gait_9e��Y�&��Qx���	�Shap��eration�0<��R67451j9:(`sGen�ms�42-f��r�p�5����2�rsgl�E��pp�G���qF�205p��5S���Ձ�retsdap�BP�O�\s�� "GCR�ö? ^�qngda�G��V��st2axU��A1a]��bad�_�>btputl/�&�|e���tplibB_��=�2.����5���gcird�v�slp���x�hex��v�rqe?�Ɵx�key��v�pm��x�us$�6�gcr��F���p���[�q27j92��v�ollismqS�k�9O�ݝ� (p#l.���t��p!o��A29$Fo8��cg7no~@�tptcls` �CLS�o�b�\�km�ai_
�s>�v�o�	�t�b���ӿ�E��H��6�1enu�501�[m��ut�ia|$calma�UR��CalMat�eT;R51%�i=1 ]@-��/V� ��Z��� �fq1�9 "K9�E�L����2m�C�LMTq�S#��et �LM3!} �F�c�nspQ�c���Oc_moq��� ��cc_e�����su���ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ���N�sve��C�clm��&Ao# �|$find�e�0STD� ter Fi�LANG���R���
��n3��z0C3en���r,���� ��J����� ���K ��Ú�=���_Ӛ���r� "FNDRК� 3��f��tguid�䙃N�."��J�tq�� �������@������J����_�� ����c��	m�Z�~�\fndr.��n#>
B2p��Z�C�P Ma�����3�8A��� c��6� ( ���N�B�������� 2�$�81��m_���"ex�z5 �.Ӛ��c��bS���efQ��	���RBT;�OPTN �+#Q�*$�r *$��*$r*$%/s#C��d/.,P�/0*ʲDPN��$���$*��Gr�$k Exc��'IF�$MASK��%93 H5�%H�558�$548 H�$4-1�$��#1(�$�0 E�$��$�-b�$���!UPDT �B�4�b�4�2�49��0�4a�3�9j0"Mx�49�4  ��4<�4tpsh���4<�P�4- DQ� �3 �Q�4�R�4�pR%0�2�r�4.b
E\���5�Ax�4��3adq\�5K979":E�ajO? l "DQ^E^�3i�Dq ��4ҲO) ?R�? ��q�5��T��3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F蠠�4��.�5y N|� �2il(in�4��31 JH1�2Q4�251ݠ�4rma	l� �3)�REo�Z_ �æOx����4��^F�?onorTf��7_ja��UZҒ4l�5rms�AU�Kkg���4�$HCd\�fͲ�eڱ�4�RE	M���4yݱ"u@�RE�R5932fO��47|Z��5lity,�Up��e"Dil\�5���o ��7987p�?�25 �3hk910 �3��FE�0=0P_>�Hl\mhm�5 ��qe�=$�^�
E�x�u�IAymptm�U0��BU��vste�y\ �3��me�b�DvI�[� Qu�:F�Ub�*_�
EL,�su��_ �Er��ox���4hGuse�E-�?�sn��������FE��,�box�����c݌,"� ������z��M��<g��pdspw)�	� �9���b���(��1���c��Y�R� � �>�P���W��������'�0ɵ�[���͂���  �� ,K@� ��A�bump�šf��B*�Box%��7Aǰ60�BBw�\��MC� (6�,f��t I�s� ST ��*��}B�����=w��"BBF
�>��`���)��\bb?k968 "�4��ω�bb�9va699����etbŠ��1X�����ed	�F�b�u�f� �sea""������'�\��,� ���b�ѽ�o6�H�
�x�$�f���!y�����Q[�! tpe�rr�fd� TP�l0o� Recov�,��3D��R64�2 � 0��C@}s�� N@��(U�rroč��yu2r��  �
  �����$$CLe� ��������������$z�_DI�GIT��������.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$j���+c:PROD�UCTM�0\PG/STKD��V&oho�zf99��D����$FEAT_�INDEX��xd���  �
�`ILECOM�P ;���#���`�cSETUPo2 <�e�b?�  N �a�c�_AP2BCK �1=�i  �)wh0?{%&c����Q�xe%�I �m���8��\� n����!���ȏW�� {��"���F�Տj��� w���/�ğS������ ���B�T��x���� ��=�үa������,� ��P�߯t������9� ο�o�ϓ�(�:�ɿ ^���Ϗϸ�G��� k� �ߡ�6���Z�l� �ϐ�ߴ���U���y� ���D���h��ߌ� ��-���Q������� ��@�R���v����)� ����_�����*�� N��r��7� �m�&�3\t�i
pP 2#p*.VRc�*��� /�ƗPC/1/F'R6:/].��/+T�`�/�/F%�/�,�`r/?�*.F��8?	H#&?e<x�/�?;STM �2��?�.K �?�=�iPendant? Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OpoO�O_:JPG _�J_�56_�O_�_�	�PANEL1.D	T�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�W�I��
TP�EINS.XML��0\���q�Custom T?oolbar	���PASSWOR�DyFRS:�\L�� %Pa�ssword Config���֏ e�Ϗ�B0���T�f� ���������O��s� �����>�͟b��[� ��'���K��򯁯� ��:�L�ۯp�����#� 5�ʿY��}��$ϳ� H�׿l�~�Ϣ�1��� ��g��ϋ� ߯���V� ��z�	�s߰�?���c� ��
��.��R�d��� ����;�M���q�� ����<���`������ %���I�������� 8����n���!� �W�{"�F �j|�/�S e��/�/T/� x//�/�/=/�/a/�/ ?�/,?�/P?�/�/�? ?�?9?�?�?o?O�? (O:O�?^O�?�O�O#O �OGO�OkO}O_�O6_ �O/_l_�O�__�_�_ U_�_y_o o�_Do�_ ho�_	o�o-o�oQo�o �o�o�o@R�ov ��;�_�� �*��N��G���� ��7�̏ޏm����&� 8�Ǐ\�돀��!��� E�ڟi�ӟ���4�ß X�j��������įS���w������B�#���$FILE_DG�BCK 1=���/���� ( �)
S�UMMARY.DyGL���MD:������Diag� Summary���Ϊ
CONSLOG�������D�ӱ�ConsoleO logE�ͫ���MEMCHECK�:�!ϯ���X�Me�mory Dat�a��ѧ�{)>��HADOW�ϣ����J���Shad�ow Chang�esM�'�-��)	FTP7Ϥ�3������Z�mmen�t TBD��ѧ0�=4)ETHERNET��������T�ӱEther�net \�figurationU��ؠ��DCSVRF��߽߫�����%��� verify� all��'�1P{Y���DIFF��p����[���%��diff]�������1R�9�K��� ����X��CH�GD������c��r����2ZAS�� ��GAD���k��z��FY3bI[�� �/"GAD���s/�����/*&UPDAT�ES.� �/��FORS:\�/�-Ա�Updates �List�/��PS�RBWLD.CM�(?���"<?�/Y�P�S_ROBOWEL��̯�?�?��?&� O-O�?QO�?uOOnO �O:O�O^O�O_�O)_ �OM___�O�__�_�_ H_�_l_o�_�_7o�_ [o�_lo�o o�oDo�o �ozo�o3E�oi �o���R�v ���A��e�w�� ��*���я`������ ���O�ޏs������ 8�͟\�����'��� K�]�쟁����4��� ۯj������5�įY� �}������B�׿� x�Ϝ�1���*�g��� ��Ϝ���P���t�	� ߪ�?���c�u�ߙ� (߽�L߶��߂��� (�M���q� ���6� ��Z������%���I� ��B�����2������h����$FIL�E_� PR� ���������MDONL�Y 1=.�� 
 ���q��� �������~% �I�m�2 ��h��!/�./ W/�{/
/�/�/@/�/ d/�/?�//?�/S?e? �/�??�?<?�?�?r? O�?+O=O�?aO�?�O �O&O�OJO�O�O�O_��O9_�OF_o_
VI�SBCKL6[�*.VDv_�_.POFR:\�_�^.P�Vision VD file�_ �O4oFo\_joT_�oo �o�oSo�owo�o B�of�o�+� ������+�P� �t������9�Ώ]� 򏁏��(���L�^�� �����5���ܟk� � ��$�6�şZ��~������
MR_GR�P 1>.L~��C4  B����	 W������*u����RHB ��2 ���� ��� ���B�����Z�l� ��C���D�������Ŀ���J�!LL#���J��;F��5US��"Qw�
����ֿ G��%�Fb��E���y.��9:�~�@]����A&�}A��O�f�?�2A���r��E�� F�@ ������ھ���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6�\b��B�Y<%���A�o=�@�0eߋ�^�A��߲� v���r������
�C� .�@�y�d������ ��������?�Z�l�v��BH�� ��R�@(��E��������
0�P=��P��V!��ܿ� �B���/ ��@�33�:��.�g&�@U�UU�U��q	>u?.�?!rX���	�-=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7��:����D�@ ?D�� Cϥ��+C������'/0- ��P/����/N��/r� �/���/�??;?&? _?J?\?�?�?�?�?�? �?O�?O7O"O[OFO OjO�O�O�O�OX�� ���O$_�OH_3_l_W_ �_{_�_�_�_�_�_o �_2ooVohoSo�owo �o�i��o�o�o�� );�o_J�j� ������%�� 5�[�F��j�����Ǐ ���֏�!��E�0� i�{�B/��f/�/�/�/ ���/��/A�\�e�P� ��t��������ί� �+��O�:�s�^�p� ����Ϳ���ܿ� � �OH��o�
ϓ�~Ϸ� �����������5� � Y�D�}�hߍ߳ߞ��� �����o�1�C�U� y��߉�������� ����-��Q�<�u�`� �������������� ;&_J\�� ��������ڟ� F�j4����� ����!//1/W/ B/{/f/�/�/�/�/�/ �/�/??A?,?e?,� �?P�q?�?�?�?�?O �?+OOOO:OLO�OpO �O�O�O�O�O�O_'_ _K_�o_�_�_�_l� �_0_�_�_�_#o
oGo .okoVoho�o�o�o�o �o�o�oC.g R�v����� 	���<�`�*< ��`�����ޏ�� )��M�8�q�\����� ��˟���ڟ���7� "�[�F�X���|���|? ֯�?�����3��W� B�{�f�����ÿ���� �����A�,�e�P� uϛ�b_�����Ϫ_�� ߀�=�(�a�s�Zߗ� ~߻ߦ�������� � 9�$�]�H��l��� ����������#��G� Y� �B�������z��� ����
ԏ:�C.g Rd������ 	�?*cN� r�����/̯ &/�M/�q/\/�/�/ �/�/�/�/�/?�/7? "?4?m?X?�?|?�?�? �?�?��O!O3O��WO iO�?�OxO�O�O�O�O �O_�O/__S_>_P_ �_t_�_�_�_�_�_�_ o+ooOo:oso^o�o �op��o�� ��$ ��o�o�~� ������5� � Y�D�}�h�������׏ ����
�C�.�/ v�<���8������П ����?�*�c�N��� r��������̯�� )��?9�_�q���JO�� ���ݿȿ��%�7� �[�F��jϣώ��� ��������!��E�0� i�T�yߟߊ��߮��� �o�o��o>�t� >��b��������� ��+��O�:�L���p� ������������' K6oZ�Z�|� ~�����5  YDi�z��� ���/
//U/@/ y/@��/�/�/�/���/ ^/???Q?8?u?\? �?�?�?�?�?�?�?O O;O&O8OqO\O�O�O �O�O�O�O�O_�O7_���$FNO ����VQ�
F0fQ} kP FLAG8��(LRRM_CHKTYP  WP���^P�WP��{QOM�P_MIN܇P����P� � XNPSSB_�CFG ?VU? ��_����S ooIUTP_�DEF_OW  ���R&hIRC�OM�P8o�$GE�NOVRD_DO�V�6�flTHR֨V d�edkd_E�NBWo k`RA�VC_GRP 19@�WCa X"_�o _1U<y� r�����	�� -��=�c�J���n��� �����ȏ����;��"�_�F�X���ibRO�U�`FVX�P��&�<b&�8�?��埘����>���  D?�јls���@@g�B�7��p�)�ԙ���`SMT
�cG�mM���� ��LQHOSTC�R19H���P��at��SM��f��\���	127.�0��1��  e ��ٿ�����ǿ@��R�d�vϙ�0�*�	a�nonymous������������(([�� � ����� r����ߨߺ�����-� ��&�8�[�I�π� ������1�C� �W�y���`�r����� �ߺ�������%�c� u�J\n������ ���M�"4F X��i����� �7//0/B/T/� ��m/��/�/�/ ??,?�/P?b?t?�? �/�?��?�?�?OO e/w/�/�/�?�O�/�O �O�O�O�O=?_$_6_ H_kOY_�?�_�_�_�_ �_'O9OKO]O__Do�O hozo�o�o�o�O�o�o �o
?o}_Rdv ���_�_oo!� Uo*�<�N�`�r��o�� ����̏ޏ�?Q&��8�J�\���>�ENT� 1I�� P!\􏪟  ���� ՟ğ�������A�� M�(�v���^������ ���ʯ+�� �a�$� ��H���l�Ϳ����� ƿ'��K��o�2�h� �ϔ��ό��ϰ���� ���F�k�.ߏ�R߳� v��ߚ��߾���1����U��y�<�QUICC0��b�t����A1�����%���2&����u�!ROU�TERv�R�d���!?PCJOG�����!192.168.0.10���w�NAME !���!ROBOT�p�S_CFG �1H�� ��Auto-s�tarted�tFTP���� ��� 2D�� hz����U� �
//./�v��� /���/�/�/�/�/ �!?3?E?W?i?�/? �?�?�?�?�?�?�� �AO�?eO�/�O�O�O �O�?�O�O__+_NO �OJ_s_�_�_�_�_
O O.OoB_'ovOKo]o oo�oP_>o�o�o�o�o o�o5GYk} �_�_�_��8o� �1�C�U�$y����� ���ӏf���	��-� ?�����Ə��� ϟ�����;�M� _�q���.�(���˯ݯ ��P�b�t�����m� ��������ǿٿ���� �!�3�E�h��{ύ� �ϱ����$�6�H�J� /�~�S�e�w߉ߛ�j� ���������*߬�=��O�a�s��YT_ERR J5
����PDUSIZ  ���^J����>~��WRD ?t���  guest}��%��7�I�[�m�$SCD�MNGRP 2K�t�������V$�K�� 	�P01.14 �8��   y�����B  �  ;����� ����������
 ������������~��`��C.gR|����  i  _�  
��������� +��������
���lZ .r���"�!l��� m
d�������_GROU���L�� �	����07EQUPOD  	պ�JV�TYa �����TTP_AUTH� 1M�� <!�iPendan�y��6�Y!KAREL:*��
-KC///A/� VISION SETT�/v/�"�/�/�/#�/�/ 
??Q?(?:?�?^?p>��CTRL Nв���5�
�.FFF9E3�?��FRS:DE�FAULT�<�FANUC We�b Server�:
�����<kO}O��O�O�O�O��WR_�CONFIG �O�� �?��I�DL_CPU_P5C@�B��7Pw�BHUMIN(\���<TGNR_IO������PNPT_SIM_DOmV�w[TPMODN�TOLmV �]_P�RTY�X7RTOL_NK 1P��� �_o!o3oEoWoio�RMASTElP��R>�O_CFG�o�i�UO��o�bCYC�LE�o�d@_AS�G 1Q����
 ko,>Pbt� ��������\sk�bNUM����<K@�`IPCH�o���`RTRY_CN�@oR��bSCRN(����Q��� �b�`��bR���Տ���$J23_DSP_EN	����?OBPROC�Un�iJOGP1SY�@��8�?��!�T�!�?*�POS�RE�zVKANJI_�`��o_�� ���T�L�6͕����C�L_LGP<�_���EYLOGGIN�`���LANGUAGE YF�7RD w���LeG��U�?⧈�x� �����=P�V�'0��$ N�MC:\RSC�H\00\��LN�_DISP V���
��������OC��R.RDzVTA{�O�GBOOK W�
{��i��ii��X�����ǿٿ���b��"��6	h������e�?�G_B�UFF 1X�]��2	աϸ���� �������!�N�E� W߄�{ߍߺ߱����߀�����J���D�CS Zr� =����^�+�ZE���������a�IO 1[
{ ُ!� �!�1�C�U�i�y��� ������������	 -AQcu�������EfPTM  �d�2/AS ew������ �//+/=/O/a/s/p�/�/��SEV�����TYP��/??y͒�RS�@"��×�FL 1\
������?�?��?�?�?�?�?/?TP�6��">�NG�NAM�ե�U`�UPS��GI}�𑪅}mA_LOAD��G %�%D?F_MOTN���O��@MAXUALRM<��J��@sA�Q�����WS ��@C �]�m�-_���MP2�7�^�
{ ر�	�!P�+ʠ�;_/��Rcr�W�_�WU�W �_��R	o�_o?o"o coNoso�o�o�o�o�o �o�o�o;&Kq \�x����� ��#�I�4�m�P��� |���Ǐ���֏��!� �E�(�i�T�f����� ß��ӟ���� �A� ,�>�w�Z�������ѯ ����د���O�2� s�^�������Ϳ����ܿ�'��BD_LDXDISAX@	��MEMO_APR@�E ?�+
 � *�~ϐϢϴ�����������@ISC ;1_�+ ��I� �T��Q�c�Ϝ߇��� ������w����>�)� b�t�[����{��� �������:���I�[� /������������o� ����6!ZlS� �s���� 2�AS'�w� ���g��.//�R/d/�_MSTR� `�-w%SCD 1am͠L/�/H/ �/�/?�/2??/?h? S?�?w?�?�?�?�?�? 
O�?.OORO=OvOaO �O�O�O�O�O�O�O_ _<_'_L_r_]_�_�_ �_�_�_�_o�_�_8o #o\oGo�oko�o�o�o �o�o�o�o"F1 jUg����� ����B�-�f�Q����u�����ҏh/MK�CFG b�-�㏕"LTARM_���cL��� σQ�N�<�ME�TPUI�ǂ����)NDSP_CM�NTh���|�  d�.��ς�ҟ|ܔ|�POSCF�����PSTOL �1e'�4@�<#�
5�́5�E�S�1� S�U�g�������߯�� ӯ���	�K�-�?����c�u�����|�SIN�G_CHK  ���;�ODAQ,�f���Ç��DEV �	L�	MC:>!�HSIZEh��-���TASK �%6�%$1234?56789 �Ϡ���TRIG 1g.�+ l6�%����ǃ�����8�p�YP�[� ��EM_IN�F 1h3�� `)AT?&FV0E0"ߙ��)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ������H�����A���AI�q�,��|���� ���ߵ����� J���n������W��� ��������"����X ��/����e�� ����0�T;x �=�as��/ �,/c=/b/�/A/ �/�/�/�/��?� ��^?p?#/�?�/�? s?}/�?�?O�?6OHO �/lO?1?C?U?�Oy? �O�O3O _�?D_�OU_�z_a_�_�ONIT�OR��G ?5� �  	EXESC1Ƀ�R2�X3�XE4�X5�X���V7�X8�X9Ƀ�RhBLd �RLd�RLd�RLd
bLd bLd"bLd.bLd:bLdTFbLc2Sh2_h2khU2wh2�h2�h2�hU2�h2�h2�h3Sh�3_h3�R�R_G�RP_SV 1i�n���(ͅ�
��3�8��r��6�_MOx�_D=R^���PL_NAME� !6��p�!�Default� Persona�lity (from FD) ��RR2eq 1j)TUX)TX��q��X dϏ8�J�\� n���������ȏڏ� ���"�4�F�X�j�|������2'�П��� ��*�<�N�`�r��<��������ү������,�>�P�b� �R�dr 1o�y �\��, �3��~�� @D�  ��?�����?䰺�㱏A'�6����;��	lʲ	 �xJ����� ��< �"�� ��(pK�K� ��K=*�J����J���J�V���Z�����rτ́p@j��@T;f���f���ұ]�l��I��p������������b��3��´  �
`�>����b����z���ΐr�Jm��
�  B�H�˱]Ӂt�q�	�� p�  �P�pQ�p��p| � Ъ�g���c�	�'� � ���I� �  {����:�È
�?È=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁ryN���  '�������@2��@�c����/�C��}C�C�@ C�������
�A���   U@<�P�R�
hǉB�b�A��j���0��������Dz۩���߹�����j���( �� -��C���'�7������q�Y����� �?�ff ���gy ��@���q+q��
>+�'  PƱj�(�����7	���|�?�����xZ�p<�
6b<߈;�܍�<�ê<� <�&J���AI�ɳ+����?fff?I�?&��k�@�.��?J<?�`�q� .�˴fɺ�/��5/ ����j/U/�/y/�/ �/�/�/�/?�/0?q��F�?l??�?�/�?+)�?�?�E��� E�I�G+� F��?)O�?9O�_OJO�OnO�Of�BL޳B�?_h�.��O�O ��%_�OL_�?m_�?�_�_�_�_�_�_�
�h��Îg>� �_Co�_goRodo�o�G#A�ds�q�C�o�o8�o|����$h]Hq���D��p3C���pCHmZZD7t���6q�q��ܶN�'�3A�A�A�R1AO�^??�$�?�K�0�±
=ç>�����3�W
=�#�W��e�����@����{����<���(�B�u�����=B0�������	L��H��F�G���G���H�U`E���C�+����I#�I���HD�F���E��RC�j=���
I��@�H�!H�( E<YD0q �$��H�3�l�W��� {��������՟��� 2��V�A�z���w��� ��ԯ�������� R�=�v�a��������� ���߿��<�'�`� Kτ�oρϺϥ����� ���&��J�\�G߀� kߤߏ��߳������� "��F�1�j�U��y� ������������0�@�T�?�Q����(�1g��3/E�����5������q�3�8�����q4�Mgs&IB�+2D�a���{�^^	���P���uP2P7Q4_A��M0bt��R����X��/   �/ �b/P/�/t/�/ *a@)_3/�/�/�%1a�?�/?;?M?_?q?  �?�/�?�?�?�?�O 2 F�$N�vGb�/�A��@X�a�`�qC��C@�o��O2���OF� �DzH@�� F�P D���O�O�ys<O!_3_E_W_i_~s?���@@pZ�.t22!:2~
 p_�_ �_�_	oo-o?oQoco�uo�o�o�o�o��Q ���+��1���$MSKCFMA�P  �5� �6�Q�Q"~��cONREL  �
q3�bE�XCFENB?w
8s1uXqFNC_Qt�JOGOVLIM�?wdIpMrd�bKE�Y?w�u�bRU�N�|�u�bSFSPDTY�avJu�3sSIGN?QtTO1MOT�Nq�b�_CE_GRP [1p�5s\r� ��j�����T��⏙� �����<��`��U� ��M���̟��🧟� &�ݟJ��C���7��� ����گ�������4��V�`TCOM_C_FG 1q}�V�p�����
P�_AR�C_\r
jyUA�P_CPL��ntN�OCHECK ?={ 	r ��1�C�U�g�yϋ� �ϯ���������	���({NO_WAITc_L�	uM�NTX��r{�[m�_E�RRY�2sy3�� &�������r��c� ��T_MO���t��, �s�$�k�3�PARAM:��u{��V[ﰽ�!�u?�� =9@3�45678901 ��&���E�W�3�c������{������� �����=�UM_RSPACE ��Vv��$ODR�DSP���jxOF�FSET_CAR9Tܿ�DIS���PEN_FILE�� �q��c֮�OPT?ION_IO���PWORK v_�ms �P(��R�Q
�j.j	 ���Hj&6$� R�G_DSBL  ��5Js�\��R�IENTTO>p�9!C��PqfA� UT_SIM_D�
r�b� V� LCT ww�bc��|U)+$_PEXE�d&RATp �vju�p���2X�j)TUX�)TX�##X d-�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O�H2�/oO�O�O�O�O@�O�O�O�O_]�<^O ;_M___q_�_�_�_�_��_�_�_o���X�O�U[�o(��(����$o�,� ��IpB` @oD�  Ua?�[cbAa?��]a]�DWcxUa쪋l;�	lmb��`�x�J�`�����a�< ��`�� ��b, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�"���� �N	 W��  '!o�:q�pC	 C�@@sBq�|�:�� m�
�!�h@ߐ�n����Z��B	 �A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�'!��(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��� ��3 ���Ӱ��ɆDT� Qy-����D � ��ӱ4�P :� L :�GP:�D :�@ :�U8�8�	8�
8�U8�8�8�8�Q8�X@:�8�8�8�8�8��:�E8�8�x�:�8�PP�:�d :�8�8�P��:�
�:�!8�"8�Q#8���:�%8�&8�U'8�(8�)8�*8�T��:�,8�-8�.8�/8�08�18�,��� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�X�(�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_d��_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п�_��� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p�������� //$)�$�PGTRACEL�EN  #!  ��" ��8&_UP z/���g!o S!�h 8!_CFG7 {g%Q#"!�x!�$J �" |"D�EFSPD |��,!!J �8 I�N TRL }�-" 8�(IPE�_CONFI� ~>g%�g!�$q�$�"8 LID�#��-74GRP s1�7Q!�#!�A ���&ff�"!A+33D��� D]� CÀ� A@+6�!�" d�$�9�9*1*0� �	 +9�-+6�? #´	C�?�;B@3A�O�?OIO3OmO"!>�T?�
5�O��O�N�O =��=#�
�O_�O_ J_5_n_Y_�O}_�_y_x�_�_�_  Dzco" 
oBo�_Roxo co�o�o�o�o�o�o �o>)bM��;�
V7.10b�eta1�$ � A�E�r�ϻ�A " �p?!{G��q>���r���0�q�ͻqB7Q��qA\�p�q��4�q�p�"�B�@�2�D�V�h�w��p�?�?)2{ȏw� ׏���4��1�j�U� ��y�����֟���� ��0��T�?�x�c��� ����ү����!o�,� ۯP�;�M���q����� ο���ݿ�(��L��7�p�+9��sF@ �ɣͷϥ�g%��� ���+�!6I�[߆��� ���ߵߠ��������� !��E�0�B�{�f�� ������������ A�,�e�P���t����� �������=( aL^����� ��'9$]�� ���ϖ������� /<�5/`�r߄ߖߏ/ >�/�/�/�/�/?�/ 1??U?@?R?�?v?�? �?�?�?�?�?O-OO QO<OuO`O�O�O�O�O ���O_�O)__M_8_ q_\_n_�_�_�_�_�_ �_o�_7oIot�� �o�o���o�o�o(/ !L/^/p/�/{*o� �������� A�,�e�P�b������� ���Ώ��+�=�(� a�L���p������Oߟ 񟠟� �9�$�]�H� ��l�~�����ۯƯ�� �#�No`oro�on��o �o�o�oԿ���8 J\ng����vϯ� ��������	���-�� Q�<�u�`�r߫ߖ��� ��������;�M�8� q�\��������z��� ���%��I�4�m�X� ��|����������� :�L�^���Z������ �����$�6�H� Swb��� ����//=/(/ a/L/�/p/�/�/�/�/ �/?�/'??K?]?H? �?��?�?f?�?�?�? O�?5O OYODO}OhO �O�O�O�O�O�O&8 J4_F_����_�_ ��_�_"4-o�O *ocoNo�oro�o�o�o �o�o�o)M8 q\������ ���7�"�[�m��? ����R�Ǐ���֏� !��E�0�i�T���x� �������_$_V_ ��2�l_~_�_�����R��$PLID_KNOW_M  �T?������SV ��U.͠�U��
� �.�ǟR�=�O������mӣM_GRP S1��!`0u��T�@ٰo�ҵ�
 ���Pзj��`��� !�J�_�W�i�{ύϟπ����������߱�MR�����T��s�w� s��ߠ޴߯߅� �ߩ߻�����A��� '��������� ������=���#��� ������}������S��{ST��1 1��U�# ���0�_ A .��,>Pb �������� 3(iL^p������2�*���<-/3 /)/;/M/4f/x/�/�/5�/�/�/�/�6??(?:?7 S?e?w?�?8�?�?��?�?MAD  �d#`PARNUM  qw�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a�OT>_CMP_��B@��P@'˥TER�_CHK'U��0˪?R$_6[RSl�¯���_MOA@�_�U_��_RE_RES_G ��>�oo8o +o\oOo�oso�o�o�o �o�o�o�o�W �\�_%�Ue Baf �S� ����S0� ���SR0��#��S �0>�]�b��S�0}���<���RV 1�����^rB@c]��t�_(@c\����_D@c[�$���RTHR_INRl��DA��˥d,�MASmS9� ZM�MN8��k�MON_QUEUE ���˦��Vx� RDNPUbQqN{�P[��END���_ڙEXE�ڕ�@�BE�ʟ��OPT�IOǗ�[��PROGRAM %���%��ۏ�O��TA�SK_IAD0�OCFG ���tO��^ŠDATA���Ϋ@��27�>�P� b�t���,�����ɿۿ������#�5�G���IWNFOUӌ���� ���ϭϿ�������� �+�=�O�a�s߅ߗ� �߻��������^�jč�� yġ?PDIT �ίc���WERFL
��
�RGADJ �&n�A����?�����@���IORITY�{�QV���MPDSQPH�����Uz��ޝ�OTOEy�1��R� (!AF�4�E�P]���!�tcph���!�ud��!icqm��ݏ6�XY_ȡ��R��ۡ)�� *+/ ۠� W:F�j�� ����%7�[B�*��POSRT#�BC۠�����_CARTR�EP
�R� SKS�TAz��ZSSAV����n�	2500H863���r�T$!�R���Áq�n�}/�/�'� U�RGE�B��rYW�F� DO{�rUVW�V��$�A�WRUP�_DELAY ��R��$R_HOT�k��%O]?�$R_?NORMALk�L?<�?p6SEMI?�?|�?3AQSKIP!��n�l#x 	 1/+O+ OROdOvO9H n��O�G�O�O�O�O�O _�O_D_V_h_._�_ z_�_�_�_�_�_
o�_ .o@oRoovodo�o�o �o�o�o�o�o*< Lr`���n��$RCVTM�v����pDCR!��LЈqCq��C�2ACĳ�u?�A�>�Rߐ<|�{4M�l��� ��´��ʿ��Ҿ�?�[�|��4Oi���O <
6b<�߈;܍�>�u.�?!<�&{�b�ˏݏ�� 8�����,�>�P�b� t���������Ο��� ݟ��:�%�7�p�S� �����ʯܯ� �� $�6�H�Z�l�~����� ��ƿ���տ���2� D�'�h�zϽ��ϰ��� ������
��.�@�R� d�Oψߚ߅߾ߩ��� ������<�N��r� ������������ �&�8�#�\�G����� }�����������S� 4FXj|��� ������0 T?x�u��� �'//,/>/P/b/ t/�/�/�/�/�/�/� ?�/(??L?7?p?�? e?�?�?��?�? OO $O6OHOZOlO~O�O�O �?�?�O�O�O�O __ D_V_9_z_�_�?�_�_ �_�_�_
oo.o@oRo�dovo�X�qGN_A�TC 1�� �AT&FV�0E0�kAT�DP/6/9/2{/9�hATA�n�,AT%G�1%B960�i�+++�o,�aH�,�qIO_TY�PE  �u�s�n_�oREFPOS�1 1�P{ x�o�Xh_�d_ �����K�6�o� 
���.���R����{{/2 1�P{����؏V�ԏz����q3 1��$�6�p��ٟ|���S4 1������˟���n���%�S5 1�<�N�`������<���S6 1�ѯ���/�����ѿ>O�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASKw 1�P  
9ߜG��XNOM����a~߈ӁqMOTE�  h�~t��_CFG ������рrPL_RANG����Q��POWER ���e��SM�_DRYPRG �%i�%��J��T?ART �
�X�UME_PRO'��9��~t_EXEC_ENB  �e��GSPD�����蜩c��TDB���R�M��MT_!�T����`OBOT�_NAME �i���iOB_O�RD_NUM ?�
�\qH?863  �T���������bPC_TIMEOUT��{ x�`S232���1��k L�TEACH PE�NDAN �ǅ��}���`Mai�ntenance Cons�R}�m
�"{�dKCL/!Cg��Z ��n�� No Us�e}�	��*NPqO��х��ӽ(CH_L��������	�mMAVAIL��{���ՙ�SPACE�1 2��| �d��(>��&����p��M,8�?�ep/eT/�/�/�/ �/�W//,/>/�/b/ �/v?�?Z?�/�?�9�e �a�=??,?>?�?b? �?vO�OZO�?�O�O�Os�2�/O*O <O�O`O�O�_�_u_�_�_�_�_[3_#_5_ G_Y_o}_�_�o�o�o �o�o[4.o@o Rodovo$�o�o��@��"�	�7�[5K ]o��A���菀	�̏�?�&�T�[6 h�z�������^�ԏ�� �&��;�\�C�q�[7��������͟{�� �"�C��X�y�`���[8����Ưدꯘ� �0�?�`�#�uϖ�}ϼ��[G �i�� �ϋ
G� ����$�6�H�Z�l� ~ߐ��8 ǳ���������d(���M� _�q�������� ���?���2�%�7�e� w��������������� �����!�RE�W�� ��������p?Q `�� @0��ߖrz	�V_��� ��
/L/^/|/2/d/ �/�/�/�/�/�/?�/ �/�/*?l?~?�?R?�? �?�?�?�?�?�?2O�?�
��O[_MO�DE  �˝IS ���vO,*Aϲ�O-_��	M_�v_#dCWORK_{AD�Ml[P%a/R  ��ϰ�P�{_�P_INTVA�L�@����JR_O�PTION�V ��EBpVAT_G�RP 2����(y_Ho �e_vo�o�oYo�o�o �o�o�o*<�bO oNDpw���� ��	���?�Q�c� u�����/���ϏᏣ� ���)�;���_�q��� ������O�ɟ��� ՟7�I�[�m�/����� ��ǯٯ믁��!�3� ��C�i�{���O���ÿ տ���ϡ�/�A�S� e�'ωϛϭ�oρ��� ����+�=���a�s� ��Gߕ߻����ߡ�� �'�9�K�]��߁�� ���y�����������5�G�Y��E�$SC?AN_TIM�AYu�ew�R �(�#((�<0.a_aPaP	
Tq>��Q���o�����O�O2/��:	dD/JaR��WY���^���^R^	r � P��� �  8�P�	<�D��G Yk}���������Qp�/@/R//)P;��o\T��Qpg-�t�_DiKT|��[  � l v%������/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OWW�#�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_olO~Od+No`o ro�o�o�o�o�o�o�o &8J\n�������u�  0�"0g�/�-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ����$o��˟ݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�����Do������ ��ҿ�����,�>� P�b�tφϘϪϼ���`������w
�  5 8�J�\�n߀ߒߜկ� ��������	��-�?�Q�c�u����� ��-����� � 2�D�V�h�z��������������������& ��%	�12345678^�" 	��/� `r��������(: L^p����� �� //$/6/H/Z/ l/~/��/�/�/�/�/ �/? ?2?D?V?h?�/ �?�?�?�?�?�?�?
O O.O@Oo?dOvO�O�O �O�O�O�O�O__*_ YON_`_r_�_�_�_�_ �_�_�_ooC_8oJo \ono�o�o�o�o�o�o �oo"4FXj�|������� ��	��s3�E�W��{�Cz  Bp���   ��2����z�$SCR_�GRP 1�(��U8(�\x�^ @ > 	!��	  ׃���"�$� ���-��+��R�w����D~�����#�����O���M-�10iA 890�9905 Ŗ5 M61C >4��J*ׁ
� ����0�����#�1�	�"�z�������¯Ҭ ���c��� O�8�J��������!�����ֿ��B�By���������A��$�  @��<� �R�?��d���Hy�u�O����F@ F�` �§�ʿ�϶������� %��I�4�m��<�l�`�߃ߕߧ߹�B��� \����1��U�@�R� ��v������������;���*<=�
�F���?�d�<�>m󙵎��@�:��� B���ЗЙ����EL_DEFA�ULT  ���_�B��MIPOWERFL  �$1 oWFDO $���ERVENT �1�����"��pL!DUM_�EIP��8��j!AF_INE <�=�!FT����!��4 ���[!RPC�_MAIN\>�8J�nVISw=y���!TP��PU��	d�?/!�
PMON_PR'OXY@/�e./�/�"Y/�fz/�/!RDM_SRV�/r�	g�/#?!R dC?�h?o?!
p�M�/�i^?�?!?RLSYNC�?8��8�?O!ROS�.L�4�?SO" wO�#DOVO�O�O�O�O �O_�O1_�OU__._ @_�_d_v_�_�_�_�_�o�_?oocoiICE_KL ?%y� (%SVCPRG1ho8��e��D�o�m3�o�o�`4 D�`5(-�`6PU�`7x}�`���l9��{�d:?� �a�o��a�oE��a�o m��a���aB���a j叟a���a�5� �a�]��a����a3� ���a[�՟�a�����a ��%��aӏM��a��u� �a#����aK�ů�as� ��a��mob�`�o�` 8�}�w�������ɿ�� �ؿ���5�G�2�k� VϏ�zϳϞ������� ���1��U�@�y�d� �߯ߚ��߾������ �?�*�Q�u�`��� ����������;� &�_�J���n������������sj_DEV� y	�M{C:P�_OUT",?REC 1�Z� �d   	 	�������
 �PJ�%6 (��&�[w�,��*  T �- �- �A�- c |�P����� //B/0/f/x/Z/�/ �/�/�/�/�/�/?�/ ?P?>?t?b?�?�?�? �?�?�?�?OOOLO :OpO�OdO�O�O�O�O �O�O�O$__H_6_X_ ~_l_�_�_�_�_�_�_ �_ ooDo2oTozo\o �o�o�o�o�o�o�o .R@vd�� ��},���� 4�"�X�F�|���p��� ��֏ď����0�� @�f�T���x�����ҟ �Ɵ���,��<�b� P���h�z������ί ��(�:��^�L�n� p�������ܿ�п�  �6�$�Z�H�jϐ�r� �Ϣ����������2� D�&�h�Vߌ�z߰ߞ� ����������
�@�.��d�R��ZjV 1-�w P�m��	�x  P ����
TYPE�VFZN_CF�G ���d7�GRP� 1�A�c ,�B� A� D;�� B���  B�4RB21^HELL:�(
� X����%RSR���� E0iT�x�� ����/S�ew�����%@w�����#�1�������2#�d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he��_ &_8_J_\_��_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}4xcopy �fr:\*.* �virt:\tm�pback�Q=>�192.168.�4�P46:697�6 �R�_�_�_�K}5�Ua�_�_�V�_go�yo�o}9�Ts:o�rderfil.dat.l@oVo�o�o�}0�Rmdb: +o�o�Q�obt�c �_2o?U��
�o ��Sod�v����o�o 6Q���+Ə O`�r����*�<�� ޟ���'���K�\��n����
xyzrate 61 +�@=�O�������>��2848 ��ү c�u�������5�6�ٿ ����"���5�ѿb��tφ��6����em}p:�2392 W�����ύ�.��*.d�������a�s߅ߘ�  +�=�O�������)� ������c�u��� 5����������"Ͻ� ����b�t��������� Q�U�����
����� T���gy����9� T���	��@�� cu���-?��� �/��N_/q/ �/�ߨ�:/L/�/�/?x�&�͐5372?� �/b?t?�?��458 �?�?�?"�?58�?�bOtO�O�ϫ?��͐4016 WO�O�O�O ߹O�I�O`_r_�_�/ ��;_M_�_�_o?'? �T�_�_couo�o�?�? 5O�G�o�o�oO"O�o �H�obt���/�/ IdV���/��6 �g�y����o�o 9T���	���@�ҏc�u������$S�NPX_ASG �1�������� P 0� '%R[?1]@1.1����?���%֟��&� 	��\�?�f���u��� �����ϯ��"��F� )�;�|�_�������ֿ ��˿���B�%�f� I�[Ϝ�Ϧ��ϵ��� ����,��6�b�E߆� i�{߼ߟ�������� ���L�/�V��e�� �����������6� �+�l�O�v������� ��������2V 9K�o���� ���&R5v Yk�����/ ��<//F/r/U/�/ y/�/�/�/�/?�/&? 	??\???f?�?u?�? �?�?�?�?�?"OOFO )O;O|O_O�O�O�O�O �O�O_�O_B_%_f_ I_[_�__�_�_�_�_ �_�_,oo6oboEo�o io{o�o�o�o�o�o �oL/V�e� �������6� �+�l�O�v��������PARAM ������ �	U��P�����OFT_KB_CFG  ヱ����PIN_SIM  ���C�U�g������RVQSTP/_DSB,�򂣟|����SR �/��� & MUL�TIROBOTTgASK������TOP_ON_E_RR  ��~�PTN /��@�A	�RING_PRM�� ��VDT_G�RP 1�ˉ�  	���������� ��Я�����*�Q� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�i�f�x��� �����������/�,� >�P�b�t��������� ������(:L ^p������ � $6HZ� ~������� / /G/D/V/h/z/�/ �/�/�/�/�/?
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8___\_���VPRG_CO7UNT��@��N�RENBU��UM�S���__UPD 1}�/�8  
s_ �oo*oSoNo`oro �o�o�o�o�o�o�o +&8Jsn�� �������"� K�F�X�j��������� ۏ֏���#��0�B� k�f�x���������ҟ ������C�>�P�b� ��������ӯί������UYSDEBSUG�P�P�)�d�Y�H�SP_PASS�UB?Z�LOG� ��U�Sr)�#�0�  ��Q~)�
MC:\��<6���_MPC���UH���Qñ8� �Q~�SAV ������ǲ&�ηS�V;�TEM_TI�ME 1��[ 5(m�=&�::�}Y�T1SVGUNS��P�U'�U���A�SK_OPTIO�N�P�U�Q�Q��BCCFG ��[�u� n�A�a�`a�gZo��߃ߕ��� ��������:�%�^� p�[���������  �����6�!�Z�E�~�@i���������&��� ����&8��nY �}�?��ԫ � �(L:p^ �������/  /6/$/F/l/Z/�/~/ �/�/�/�/�/�/�/2? 8 F?X?v?�?�?? �?�?�?�?�?O*O<O 
O`ONO�OrO�O�O�O �O�O_�O&__J_8_ n_\_~_�_�_�_�_�_ �_o�_ o"o4ojoXo �oD?�o�o�o�o�oxo .TBx�� j������� �,�b�P���t����� Ώ��ޏ��(��L� :�p�^�������ʟ�� o��6�H�Z�؟ ~�l�������د��� ʯ ��D�2�h�V�x� z���¿���Կ
��� .��>�d�Rψ�vϬ� ���Ͼ�������*�� N��f�xߖߨߺ�8� ��������8�J�\� *��n�������� ����"��F�4�j�X� ��|����������� ��0@BT�x �d����� >,Ntb��� ���/�(//8/ :/L/�/p/�/�/�/�/ �/�/�/$??H?6?l? Z?�?~?�?�?�?�?�? O�&O8OVOhOzO�? �O�O�O�O�O�O
__ �O@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<o^o�oro�o�o�o �o�o�o J8 n$O�����X ���4�"�X�B�v���$TBCSG_�GRP 2�B���  ��v� 
 ?�  ������׏����叀��1��U�g�z����~��d, ����?v�	 HC���d�>����e�CL  B���Пܘ���\)>��Y  A�ܟ$�3B�g�B�Bl�i��X�ɼ���X��  �D	J���r�����C ����үܬ���D�@v�=�W�j�}�H�Z� ��ſ����������v�	V3.�00��	m61c�	*X�P�u�Lg�p�>���v�(:��� ��p͟�  O����p������z�JCFG ȖB��� �����������=��=�c�q�K�qߗ� �߻ߦ��������'� �$�]�H��l��� ���������#��G� 2�k�V���z������� �������p*< N���l���� ���#5GY }h����v�b� �>�// /V/D/z/ h/�/�/�/�/�/�/�/ ?
?@?.?d?R?t?v? �?�?�?�?�?O�?*O O:O`ONO�OrO�O�O ��O�O�O_&__J_ 8_n_\_�_�_�_�_�_ �_�_�_�_oFo4ojo |o�o�oZo�o�o�o�o �o�oB0fT� x������� ,��P�>�`�b�t��� ��Ώ�������&� L��Od�v���2����� ȟʟܟ� �6�$�Z� l�~���N�����دƯ �� �2��B�h�V� ��z�����Կ¿�� ��.��R�@�v�dϚ� �Ϫ��Ͼ������� <�*�L�N�`ߖ߄ߺ� �����ߚ������� \�J��n����� �����"���2�X�F� |�j������������� ��.TBxf ������� >,bP�t� ����/�(// 8/:/L/�/�ߚ/�/�/ h/�/�/�/$??H?6? l?Z?�?�?�?�?�?�? �?O�?ODOVOhO"O 4O�O�O�O�O�O�O
_ �O_@_._d_R_�_v_ �_�_�_�_�_o�_*o oNo<oro`o�o�o�o �o�o�o�o&�/> P�/����� ����4�F�X�� (���|�����֏��� �Ə0��@�B�T��� x�����ҟ������ ,��P�>�t�b����� ����������:� (�^�L�n�������2 d�����̿�$�Z� H�~�lϢϐ������� �Ϻ� ��0�2�D�z� �ߞ߰�j��������� �
�,�.�@�v�d�� ������������ <�*�`�N���r����� ��������&J \�t��B�� ����F4j |��^�����/�  2 6#� 6&J/6"�$T�BJOP_GRP� 2���  ?�X,�i#�p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�ق'�!�!>��͘
559>�0+1��33=�CL�� fff?+0?�ffB� J1�%Y?d7z�.��/>��2�\)?0�5���;��hCY� ��  @� �!B�  A�P?�?�3E?C�  D�!�,�0*BOߦ?�3JB���
:���Bl�0��0�$�1�?O~6!Aə�AДC�1D�G6�=q��E6O0�p��B��Q�;�AȾ� ٙ�@L3D�	�@�@__�O�O>�B�\JU�OHH�1t�s�A@33@?1� C�� �@�_�_<&_8_>��D�UV_�0�LP�Q30<{�	�zR� @�0�V�P!o 3o�_<oRifoPo^o�o �o�oRo�o�o�o�o M(�ol�p~���p4�6&�q5	�V3.00�#om61c�$*(��$1!6�A� E�o�E��E���E�F���F!�F�8��FT�F�qe\F�NaF����F�^lF����F�:
F��)F��3G��G��G��G,IR��CH`�C�dT�DU�?D���D��DE(!/�E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[
�F���F��M�;S@;Q��|8��`rz@/&�8��6&<��1�w�^$E�STPARS  �*({ _#HR��A�BLE 1�p+$Z�6#|�Q� � 1�
|�|�|�5'=!|�	|�
|�|�˕6!U|�|�|���'RDI��z!ʟܟ � ��$���O����@��¯ԯ�����S��x# V���˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������U- ����ĜP�9�K�]�o� �-�?�Q�c�u���6ҿNUM  �Uz!� >  Ȑ�����_CFG ������!@b IM?EBF_TT����8x#��a�VER��b�zw�a�R 1�p+O
 (3�6"1 ��  6!�������� �� �9�$�:�H�Z�l� ~���������������H^$��_��@x��
b MI_CHA�Nm� x� kDB'GLV;0o�x�a!�n ETHERADW ?�� �y��$"�\&n RO�UT��!p*!�*�SNMAS�K�x#�255�.h�fx^$OOLOFS_DI���[ՠ	ORQCTRL �p+;/� ��/+/=/O/a/s/ �/�/�/�/�/��/�/��/!?��PE_DE�TAI��PON?_SVOFF�33�P_MON ��H�v�2-9STRT�CHK ����42VTCOMP�ATa8�24:0FP�ROG %�%�MULTIROBOTTO!O06��PLAY��L:_I_NST_MP GL7YDUS���?�2�LCK�LPKQUI�CKMEt �O�2S�CRE�@�
tps��2�A�@�I��@_Y���9�	�SR_GRP 1}�� ���\�l_zZg_�_�_�_�_�_�^�^�oj�Q 'ODo/ohoSe��oo �o�o�o�o�o�o !WE{i�������	1234567��!����X�E1�V[
 �}ipnl/a�gen.htmno���������ȏ~��Panel setup̌}�?��00�B�T�f� ��� ����ԟ���o�� ��@�R�d�v������ #�Я�����*��� ϯůr���������̿ C��g��&�8�J�\� n�����϶������� ��uϣϙ�F�X�j�|� �ߠ����;��������0�B��*NUAL{RMb@G ?�� [�������� ���� ��%�C�I�z��m�������v�SEV7  ����t�ECFG Ձ=�]/BaA$   ;B�/D
 ��/C �Wi{�������� PRֆ�; �To\o�I2�6?K0(%��� �0�����// ;/&/L/q/\/�/�/�/�l�D �Q�/I�_�@HIST 1}ׁ9  ( � ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,?153,1 Ec0�p?�?�?�?/C�� >?P=962n?�?
O`O.O�?�?�136c? |O�O�O�OAOSO�?�O __0_�O�O_Lu_�_ �_�_:_�/�_�_oo )o;o�__oqo�o�o�o �oHo�o�o%7I~��a81�ou�� ����o���)� ;�M��q��������� ˏZ�l���%�7�I� [���������ǟٟ h����!�3�E�W�� ��������ïկ�v� ��/�A�S�e�Pb ������ѿ������ +�=�O�a�s�ϗϩ� ��������ߒ�'�9� K�]�o߁�ߥ߷��� �����ߎ�#�5�G�Y� k�}���������� �����1�C�U�g�y� ��v�����������	 �?Qcu�� (����) �M_q���6 ���//%/�I/ [/m//�/�/�/D/�/ �/�/?!?3?�/W?i? {?�?�?�?�����?�? OO/OAOD?eOwO�O �O�O�ONO`O�O__ +_=_O_�Os_�_�_�_ �_�_\_�_oo'o9o Ko�_�_�o�o�o�o�o �ojo�o#5GY �o}������?���$UI_PA�NEDATA 1�������  	�}��0�B�T�f�x��� )����mt�ۏ��� �#�5���Y�@�}��� v�����ן��������1��U�g�N������ �1��Ïȯگ ����"�u�F���X� |�������Ŀֿ=��� ���0�T�;�x�_� �Ϯϕ��Ϲ������,ߟ�M��j�o߁� �ߥ߷������`�� #�5�G�Y�k��ߏ�� ������������� C�*�g�y�`������� ��F�X�	-?Q c����߫��� �~;"_F ��|����� /�7/I/0/m/���� �/�/�/�/�/�/P/!? 3?�W?i?{?�?�?�? ?�?�?�?O�?/OO SOeOLO�OpO�O�O�O �O�O_z/�/J?O_a_ s_�_�_�_�O�_@?�_ oo'o9oKo�_oo�o ho�o�o�o�o�o�o�o #
GY@}d� �&_8_����1� C��g��_�������� ӏ���^���?�&� c�u�\�������ϟ�� �ڟ�)��M��� ��������˯ݯ0�� ���7�I�[�m���� ������ٿ�ҿ��� 3�E�,�i�Pύϟφ�`�Ϫ���Z�l�}���@1�C�U�g�yߋ�)� ��#������� ��$� 6��Z�A�~�e�w�� ����������2���V�h�O�����v�p���$UI_PANELINK 1�v��  ��  ��}1�234567890����	-?G  ���o����� a��#5G�	�����p&���  R�����Z ��$/6/H/Z/l/~/ /�/�/�/�/�/�/�/ 
?2?D?V?h?z??$? �?�?�?�?�?
O�?.O @OROdOvO�O O�O�O �O�O�O_�O�O<_N_``_r_�_�_�0,�� �_�X�_�_�_ o2oo VohoKo�ooo�o�o�o �o�o�o��,> r}�������� ����/�A�S�e� w��������я��� tv�z����=�O� a�s�������0S��ӟ ���	��-���Q�c� u�������:�ϯ�� ��)���M�_�q��� ������H�ݿ��� %�7�ƿ[�m�ϑϣ� ��D��������!�3� Eߴ_i�{�
�߂��� �߸������/��S� e�H���~��R~'� '�a��:�L�^�p� ��������������  ��6HZl~� ��#�5���  2D��hz��� ��c�
//./@/ R/�v/�/�/�/�/�/ _/�/??*?<?N?`? �/�?�?�?�?�?�?m? OO&O8OJO\O�?�O �O�O�O�O�O�O[�_ ��4_F_)_j_|___�_ �_�_�_�_�_o�_0o oTofo��o��o� �o�o�o,>1 bt����K� ���(�:���� {O������ʏ܏�uO �$�6�H�Z�l����� ����Ɵ؟����� � 2�D�V�h�z�	����� ¯ԯ������.�@� R�d�v��������п ���ϕ�*�<�N�`� rτ��O�Ϻ�Io���� �����8�J�-�n߀� cߤ߇����߽���� o1�oX��o|��� �����������0� B�T�f���������� ����S�e�w�,>P bt��'��� ��:L^p ��#���� / /$/�H/Z/l/~/�/ �/1/�/�/�/�/? ? �/D?V?h?z?�?�?�? ??�?�?�?
OO.O�� ROdO�߈OkO�O�O�O �O�O�O_�O<_N_1_ r_�_g_�_7OM��m�$UI_QU�ICKMEN  }��_�AobRESTOR�E 1�  �|��Rto�o�im�o�o�o �o�o:L^p �%������o ����Z�l�~��� ��E�Ə؏���� � ÏD�V�h�z���7��� ����/���
��.�@� �d�v�������O�Я �����ßͯ7�I� ��m�������̿޿�� ��&�8�J��nπ� �Ϥ϶�a�������Y� "�4�F�X�j�ߎߠ� �������ߋ���0�xB�T�gSCRE`�?#mu1�sco`u2��3���4��5��6��7��8��bUSER�q�v��Tp���ksT����4��5��6���7��8��`NDO_CFG �#k�  n` `PD�ATE ����NonebS�EUFRAME � �TA�n�RTOL_ABRTy��l��ENB����G�RP 1�ci/a?Cz  A�����Q�� $6HRd��`U�����?MSK  ������Nv�%�U�%����bVISCA�ND_MAX��I��FAILO_IMG� �PݗP�#��IMREG�NUM�
,[S�IZ�n`�A��,VONTMOU4��@���2���a��a�����FR:\� � M�C:\�\LOGn�B@F� !��'/!+/O/�Uz �MCV�8#7UD1r&EX{+�S��PPO64_t��0'fn6PO��LIb�*r�#V���,f@�'޻/� =	�(SZ�V�.����'WA�I�/STAT ����P@/�?�?��:$�?�?��2D�WP  ��P� G@+b=���� H�O_JMP�ERR 1�#k
�  �2345678901dF�ψO {O�O�O�O�O�O_�O *__N_A_S_�_
� MLOWc>
 �g_TI�=�'�MPHASE  ���F��PSH�IFT�1 9�]@<�\�Do�U#o Io�oYoko�o�o�o�o �o�o�o6lC U�y������ ��	�V�-�e2�����	VSFT1��2	VM�� S�5�1G� ���%�A�  B8̀�̀�@ pكӁ˂�у��z�ME@�?�q{��!c>&%�a�M1��k�0�{ ��$`0TDINEND��\�O� �z�����S��w��P�{��ϜRELE�Q��Y���\�_AC�TIV��:�R�A ��e���e�:��RD� ���YBO�X �9�د�6���02����190.0.�8�3��254t��QF�	 ��X�j��1�r�obot���   p�૿�5pc��̿������7�����-�f�ZA+BC�����,]@U� �2ʿ�eϢωϛϭ� ������ ���V�=� z�a�s߰�E�Z��1�Ѧ