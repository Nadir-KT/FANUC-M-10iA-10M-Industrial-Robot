��   �S�A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����SBR_T �  | 	$SVMTR_ID $ROBOT9�$GRP_N{UM<AXISQX6K 6NFF3 �_PARAMF	�$�  ,�$MD SPD_L�IT  �$$C�LASS  ������ � � VIRTUAL�\�'  1 �� � 8����ARC Mate� 100iC���aiS8/�4000 40A���	H1 DS�P1-� ��	P�01.14, � 	���
_PCR�� ��C������0��{  ����r���3!M�����  H� � ����?
/m��� �X�� O]]��m��� �R �2.h��>�����7(���h����&���
= �b 	���� �6���b�����g�m 2 � ���y���|�߄�.���Z�B� � �d UG c ��8 :�?�� :
�(/�/�/�/�/��1��/��f?&?x8?J?��2D+��������g�^�2�&���<�"���a?S? �?�"%7�2AMHZl�=P������v��W 5��*�*��r@���? 3!���=��y���p�c5�\��Z r 
���� /$y��?VCd ?'���WB��+"W&�a/s/UD�/ U_g_y_�_�/�_
?�_��_�_	o 4�����<]����W����1�1=��>���� ?�2oVo�T�t�?�22/5�1�223AJ OO�|��r��~!����{���ED�<��9"�R8 �l� �� �&��3 ����� �=w2��(Y5`^�N p�� ��Y���@= � ���� <$��]oVC �}@@'B���Dri��l�W&ic9	`�t # (%Q_� ��/Tq��a���"�4� F��_j��_������ď ֏������8Buo�biS0O.5/6�k=4A�K�o�nq�� ���_�o��H�g��HEAr����	sp 8 ������|�B7~��D
�|�� �� �+$|pL��rB��z?#~ ��n���
l}����s�p2 %Q��x"��b�����
	P�֯� ��U��y�B�T�f�x� ���������:Q)��O�RR�=5BA2F������8���8�p<��͛ m�{�� ��@�������I�[��t�; $���
�/�l��M���� �����ߚ߬����+� ����*�<�N�`�r�&�����76!��?9�Kϥ� ��ym���0�;L���ϹϘ�������ɧ���o l�?#�;���~a��.5صA�S�e�w�@R d�߈�ߙ�����*<|����=GBR�Qgv	v�� p�����	// -/?/Q/c/u/�/�/�/@�/�/�/�/?<�? 9?K?]?o?�?�?�?�? �?�?�?�3oaO� ��qO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_#?�_ �_o!o3oEoWoio{o �o�o�?-OO�oCOUO /ASew�� �������+� =�O�a�s��_������ ͏ߏ���'�9�K� ]��o��u��o۟ ����#�5�G�Y�k� }�������ůׯ��� ��1���U�g�y��� ������ӿ���	�� ����3ϭ���џ�ϫ� ����������)�;� M�_�q߃ߕߧ߹��� ����K��%�7�I�[� m�������#�U� G��k�}�E�W�i�{� �������������� /ASew�� �߭���+ =Oas���� �)�;�//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?� }?�?�?�?�?�?�?�? OO1OCO��[O� ���O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oos?;o Mo_oqo�o�o�o�o�o �o�oKO}OoO8�O�O m������ ��!�3�E�W�i�{� ������ÏoՏ��� �/�A�S�e�w����� ��	ҟş?Qc+� =�O�a�s��������� ͯ߯���'�9�K� ]�o���ݏ����ɿۿ ����#�5�G�Y�k� �ٟ�����!����� ��1�C�U�g�yߋ� �߯���������	�� -�?c�u���� ����������sϥ� ��`����ϕ������� ����%7I[ m������ G��!3EWi{ �����1��� g�y���S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O//�O%/ 7/I/_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogo�?�o �o�o�o�o�o�o	 -?�O�O�O��O�O ������)�;� M�_�q���������ˏ ݏ���oo%�I�[� m��������ǟٟ� ��Y"�����{� ������ïկ���� �/�A�S�e�w����� ����ѿ-�����+� =�O�a�sυϗϩϻ� 7�)���M�_�q�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }��뿳��������� ��1�C�U�g����� �ϰ�������	 -?Qcu��� ����); ��Mq����� ��//%/��J/=/ �������/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?U O/OAOSOeOwO�O�O �O�O�O�O_/Q/�Ou/ �/�/a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�oO�o �o�o#5GYk }��O__�3_E_ ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c��ou����� ��ϟ����)�;� M��r�e����˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�}�E�W�i�{� �ϟϱ���������� ��y�#ߝ������ߛ� �߿���������+� =�O�a�s����� ����;���'�9�K� ]�o����������E� 7� [�m�5GYk }������� 1CUgy� ������	// -/?/Q/c/u/���/�/ +�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO� mOO�O�O�O�O�O�O �O_!_3_�/�/K_�/ �/�/�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�ocO+ =Oas���� ��;_m___(��_�_ ]�o���������ɏۏ ����#�5�G�Y�k� }�������ş��� ��1�C�U�g�y��� ���¯��/�A�S�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�q�͟�ϧϹ��� ������%�7�I�[� ׯɯs��������� ���!�3�E�W�i�{� ������������� �/���S�e�w����� ����������cߕ� ��P�߽߅��� ���'9K ]o������ 7��/#/5/G/Y/k/ }/�/�/�/�/!�/�/ Wi{C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O� �O�O�O�O__)_;_ M___q_�_�/�/�_? '?9?oo%o7oIo[o moo�o�o�o�o�o�o �o!3EW�O{ �������� �/��_�_�_x��_�_ ����я�����+� =�O�a�s��������� ͟ߟ��_�9�K� ]�o���������ɯۯ �I��������k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ��������	�� -�?�Q�c�u߇ߙ߫� '����=�O�a�)�;� M�_�q������� ������%�7�I�[� m���ϣ��������� ��!3EW���� �ߠ������ /ASew�� �����//+/ ��=/a/s/�/�/�/�/ �/�/�/??q:?-? ����?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�OE/ __1_C_U_g_y_�_ �_�_�_�_O?A?�_e? w?�?Qocouo�o�o�o �o�o�o�o); M_q���_� ����%�7�I�[� m���_o�_ȏ#o5o ���!�3�E�W�i�{� ������ß՟���� �/�A�S��e����� ����ѯ�����+� =���b�U�Ϗ�󏻿 Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����m�5�G�Y�k� }ߏߡ߳��������� w�i�����y�� �����������	�� -�?�Q�c�u������� ����+���); M_q����5� '��K�]�%7I[ m������ �/!/3/E/W/i/{/ ���/�/�/�/�/�/? ?/?A?S?e?��?}? �	�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_�/ ]_o_�_�_�_�_�_�_ �_�_o#o�?�?;o�? �?�?�o�o�o�o�o�o 1CUgy� ������S_� -�?�Q�c�u������� ��Ϗ+o]oOo�so�o M�_�q���������˟ ݟ���%�7�I�[� m���������ٯ� ���!�3�E�W�i�{� ��鏲����1�C�� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a߽��ߗߩ߻� ��������'�9�K� ǿ��c�ݿ������ �����#�5�G�Y�k� }��������������� {�CUgy� ������S�� w�@���u��� ����//)/;/ M/_/q/�/�/�/�/�/ '�/??%?7?I?[? m??�?�?�?�?�? GYk3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�/ �_�_�_�_�_oo+o =oOoaoso�?�?�oO O)O�o'9K ]o������ ���#�5�G��_k� }�������ŏ׏��� ��{k