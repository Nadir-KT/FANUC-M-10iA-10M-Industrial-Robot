��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5�AUTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6*_�7_�8_�94F;CO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"YtP_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0��1p�3W >��DC �� Ќ@��hPV���mEX�p� �0g0xۤ�p�r
$TF��2C$MD3i�TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F�"FB�>�@�a2 �@$�PPU�3N�)ύRևAXd�!DU��AI�3�BUF�F=�@1c |pp���pPIT�� PP�M�M��y��F�SIMQSI�"ܢVAڤT�8�A@�w T�`(z�M��P�B�qFAC5Tb�@EW�P1��BTv?�MC�k �$*1JB`p�*1DEC��F��żp�� �H0CHNS_EMP1�G$G��8��@_4��3�p|@P��3�TC c�(r/�0-sx��ܐ�� MBi��!����JR|� i�SEGFR���Iv �aR�TpN�C��PVF��?�bx &��f{u Jc!�Ja��� !28�ץ8�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb��Ӏq�۽�н����Lp�3�B���CRC�e�3CCp����c� �mcҞb�1J�cѿ�.�T���D$ICb�Cq��5r�ե��@v�'���E�V���zF��_��FR,pN��ܫ�?�84�0A�! �r�� �h�Ϩ��p�2�͕a��� �دp�R�Dx Ϗ��o"2�7�!ARV�O`C�$LG�pV�B�1�P��@�t�aA�0'�|�+01Ro�� MEp`"1� CRA 3 A�ZV�g6p�O �FCCb�`�`F�`K������ADI��a� A�bA'�.p��p�`��c�`S4PƑ�a�AMIP��-`Y�3P�M��]pUR��QUA1  ]$@TITO1/S�@S�!����"0�DBOPXWO��B0!5��$SK���2��D�Bq�!"�"�PR�� 
� =����!g# S q1$2�S$z���L�)$�/H���� %�/�$C�!9&?�$ENE�q.c'*?�Ú RE�p�2(H ��O��0#$L|3$$@�#�B[�;���FOs_D��ROSr��#������3RIG7GER�6PApS��>��ETURN�2�c�MR_8�TUw�\�0EWM��M�cGN�P���BLAH��<E���P��&$�P� �'P@�Q3�CkD{��DQ���4�1�1��FGO_AWA�Y�BMO�ѱQ#!��DCS_�)7  �PIS� I  gb {s�C��A��[ �B$�S��AbP�@r�EW-�TNTVճ�BV�Q[C�(c`�UW�r�P�J��P�$0��S�AFE���V_SV>�bEXCLU�砝nONL2��SY��*a&�OT�a'�HI_V�4��B����_ *P0� 9�_�z��p ���ASG�� +nrr�@�6Acc*b��G�#@E�V�.iHb?fANNUNX$0.$fdID�U�2�SC@�`�i�a��jP�fp�z��@I$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6�a�bMS�W�E. 8Q�KE3YI5���TM�10s�qA�vIN��#��"���/ D��HOST_P!�rT��t�a��tn��tsp�pEMXӰV����pLc �ULI�0  �8	=ȳ#�l�D�Tk0�!1 � �$S��ESAMPL���j�۰f璱f���I��0��[ $SUB �k�#0�C��T�r#a�SAVʅ��c����C��P�fP$n0E��w YN_B#2� 0Q�DI{dlpO�(��9#$�R_�I�� �ENC�2_S� 3  5�C߰�f�- �SpU����!4�"g�޲r�1T���5X� j`ȷg��0�0K�4�<AaŔAVER�qĕ�9g�DSP�v��PC��r"��(���ƓoVALUߗHE��ԕM+�IPճ��OkPP ��TH���֤��P�S� �۰F��df�J� �uC1�+6 H�bLL_DUs�~a3@{��3:���OTX"����sȣR_NOAUkTO�!7�p$)�H$�*��c4�(�C`%8�C, �"p�&��L�� 8H *8�LH <6����c "�`, `Ĭ�kª�q���q��sq��~q��7*��8��9��0����U1��1̺1ٺ1�U1�1 �1�1ʥ2(�2����2̺2�ٺ2�2�2 �2��2�3(�3��3T��̺3ٺ3�3�U3 �3�3�4()���?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?�p�@P?9��5�9�E�@A�x��A�z� ;p$TP�?$VARI:�Z�n��UP2�P< ���TDe���K`Q�����Ќ�BAC��"= T�p��e$)�_,�bn�kp+ IFI@G�kp�H  ��P��"F@`�!>t� ;E��sC�ST�D� D���c�<� 	C��{��_����l���R  ���F?ORCEUP?b���FLUS�`H�N�>�F ���RD_CM�@E������ ��@v\MP��REMr F�Q���1k@���7Q
Kr4	NJ�5EFFۓ�:�@IN2Q��OV�O�OVA�	TR3OV���DTՀ�DTMX� ��@ �
ے_PH"p��CL��_TpE�@�p2K	_(�Y_T��v*(��@A;QD� ������!0tܑ0RQ���_�a����M�7�CL�dρR�IV'�{��EAR6ۑIOHPC�@��2��B�B��CM9@����R �GCLF�e!DYk(M�ap#5TuDG��� ̑%��SSD �s? �P�a�!�1���P_(�!�(�!1��E�3�!�3�+5�&�GRA���7�@��;�PW泅ONn��EBU�G_SD2H�P{�_/E A`�=�_�TERM`5Bi5���ORI#:e0C�9SM_�P��Ze0D�9TA�9E�9�UP\�F� -��A{�AdPw3S@B�$SEG�:� EL�{UUSE�@NFIJ�B$�;1젎4�4�C$UFlP=�!$,�|QR@��_G�90Tk�D�~SNST��PAT����AP'THJ��E�p% B`�'EC���A�R$P�I�aSHFT�y�A�A�H_SHOQRР꣦6 �0$�7rPE��E�OVR=���aPI�@�U�b �QAYLOW����IE"�r�A��?���ERV��XQ�Y��mG�>@�BN��U\��Rz2!P.uASYMH��.uAWJ0G�ѡE q�A�Y�R�Ud>@ ��EC���EP;�uP�;�6WOR>@M`�] 0SMT6�G3�cGR��13�aPAL@���`�q�uH � u���TOCA��`P	P�`$OP@����p�ѡ�`0YO��RE�`R4Cb�AO�p낎Be�`�R�Eu�h�A��e$7PWR�IMu�R�R_�c��q=B �I&2H���p_AD�DR��H_LENAG�B�q�q�q$�R��S�JڢSS��SKN��u\��u̳�uٳ�SE�A�����HS��MN�!K������b����O�LX��p����`ACRO3pJ�@��X��+��Q��6�OUP3�b_�IX��a�a1��}򚃳���(�� H��D��ٰ��氋�VIO2S�D�������`�7�L �$d��`Y!_OFF�r�PRM_��~b��HTTP_+��H:�M (|pOB�J]"�p��$��L�E~Cd���N �s ��֑AB_��TqᶔS�`H�L�Vh�KR"uHIoTCOU��BG�LO�q���h��0���`��`SS� ��G�HW�#A:�Oڠ}<`INCPU2VISIOW�͑���n��to��to�ٲ ��IOLN��P 8���R��p$SLzob PUT_n�$p��P& ¢��^Y F_AS�"Q��$L������Q  U�0	P4A��^���ZPHY��-��x��sUOI �#R `� K����$�u�"pPpk���$������/�UJ5�S-���N�E6WJOGKG̲D{IS��pe�Kp�L��#T (�uAVF��+`�CTR�C
�F�LAG2NE�LG�dU ���؜�~13LG_SIZ�����b�4�a��a�FDl�I`�w� m�_�{0 a�^��cg���4������Ǝ���{0��� SC�H_���a �LNT�d�VW���E�"����4��UM�Aљ`�LJ�@�DAUf�E�AU�p��d|�r�GH��b/���BOO��W�L ?�6 ITp��y0�REC��GSCR ܓ�D
�<\���MARGm�!���զ ��d%�����S�����W���U� �J{GM[�MNCHJ���FNKEY\�Kn��PRG��UF���7P��FWD��HL.��STP��V��=@X��А�RS��HO`����C9T��b ��7�[�UL���6�(RD�� ����Gt��@POЛ�������MD�FO{CU��RGEX���TUI��I��4� @�L�����P@����`��P��NE���CANA��Bj�V7AILI�CL !�U?DCS_HII4�D�s�O�(!�S����S���(���_BUFF�!Xj�?PTH$m�@��v`�ěԃ�AtrY�?P��j�3��`WOS1Z2Z3Z�D��� � Z � ���[aEȤ��ȤIKDX�dPSRrO�X��zA�STL�R}��Y&�� Y$E�C���K�&&88�п![ LQ�� +00�	P���`#qdt
��U�dw<���_ \ �`4Г�\��Ѩ#��MC4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#b�D���'B�LD�%�$�%ORGڰ5�2��PVŇVY8�s�T�r �#}d^ ���$6��$�%S�`T� �B0��4�6RCLMC��4]?o?�9세�MI��p}d_ d=њR�Q��DSTB��p� ;F�HHA�X�R JHdLEXGCESr��BM!p
�a`ip/B�T�F�j�`a�p=F_A7J�i��KbOtH�0K�db� \Q���v$MB�C�LI|�)SREQUIR�R�a.\o�AXODEBUZ�ALt M��c�b�{P����2ANDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��XB� N&��aZ���UwPST� ezr7LOC�RIrp�EX<fA�p�9AA�ODAQ��f XfY�OND�rMF,� �Łf�s"��}%�e/�� ���FX3@IGG>�� g ��t"���ܓs#N�s$R�a%��iL��hL�v�@��DATA#?pE��%�tR��Y�Nh t $MD`qI}�)nv� ytq�yt�HP`�Pxu��(�zsANSW)�yt@��yu�D+�)\b���0o�i[ �@CUw�V�p� 0XeRR2��j �Du�{Q��7Bd$C'ALIA@��G���2��RIN��"�<NE�NTE��Ck�r`^�آXb]���_N�q�lk���9�D���Bmn��DIVFDH�@t���qnI$V,���S�$��$Z �X�o�*�����oH �$BE�LT�u!ACCE�L�.�~�=�IR!C�� ���D�T�8��$PS�@�"L  Šp��#^�S�Eы T�PATH3���I�"��3x�p�A_W���ڐ���2nC��4�_{MG�$DD��<T���$FW�Rp`9��I�4��DE7��PPABN��ROTSPEE�[g�� J��[�C@4�x�?$USE_+�VPi��SYY���1- qYN!@A�Ǧ�OFF�qǡMOUf��NG���OL����INC�tMa6���HB��0HBENCS�+�8q9Bp�4�FDm�IN�Ix�]��B���VE��#�y�23_�UP񕋳LOWL����p� B���D�u�9B#P`�x ���BC<v�r�MOSI��B�MOU��@�7PERoCH  ȳOV�� â
ǝ����D��ScF�@MP����� Vݡ�@y�j�LUk��Gj�p�UP=ó���Ķ�TRK��AYLOA�Qe��A��x���p��N`�F�RTI�A$��MOUІ�HB�B S0�p7D5���ë��Z�DUM2ԓS�_BCKLSH_Cx�k����ϣ����=���ޡ �	ACLAL"q��1м@�էCHK� �S�RTY��^�%E1Qq9_�޴_UM�@�9C#��SCL0�r��LMT_J1_LD��9@H�qU�EO��p�b�_�e�k�e�SP�C��u���N�PC��N�Hz \P��C��0~"XT��CN�_:�N9��I�SF!�?�V���U�/����x�T���CB!�SH �:��E�E1T�T��`��y���T��PA �&�_P��_� =�@�����!����J6 1L�@��OG�G��TORQU��ON ֹ��E�R��H�E�g_W2���_郅����I�I�I��Ff`xJ�1�~1�VC3�0BD:B��1�@SBJR�KF9�0DBL�_SM��2M�P_sDL2GRV�`���fH_��8d���COS���LNH��� �����!*,�a1Z���fMY�_(��TH��)THE{T0��NK23��ت"��CB�&CB�CAA�B�"��!�!�&SB� 2�%GTS�Ar�CIMa������,4#97#$DU���H\1� �:B�k62�:AQ(rSf$N	E�D�`I��B+5��$̀�!A�%�5�78���LPH�E�2���2SC%C%@�2-&FC0JM&̀V�8QV�8߀LVJV!KUV/KV=KVKKVYKVgIH�8FRM��T#X!KH/KH=KHKKUHYKHgIO�<O�8�O�YNOJO!KO�/KO=KOKKOYKOM&F�2�!+i%0d�7�SPBALANC�E_o![cLE0H_�%SPc� &�b&|�b&PFULC�h`�b�g�b%p�1k%��UTO_��T13T2�i/�2N��"� {�t#�Ѱ`�0�*��.�T��OÀ<�v I�NSEG"�ͱREqV4vͰl�DIF��f��1lzw��1m�0�OBpq�я?�MI�{���nLCHWA�RY�_�AB��!�$MECH�!o �,�q�AX��P���8�7Ђ�`n 
�d�(�U�ROB��CR�x�H����(�M�SK_f`�p P+ �`_��R/�k�z�����1S�~�|�z��{���z��qINUq��MTCOM_C|� �q  ����pO�$NORE�n����pЂr �8p GRe�uSD��0AB�$XY�Z_DA�1a���D�EBUUq������su z`$��COD��G L���p��$BUFIND�X|�  <�MO�Rm�t $فU A��֐���\�<���rG��u � ?$SIMUL  S��*�Y�̑a�OBJE|�`̖ADJUSꘞݐAY_IS�Dp�3����_FI�=��Tu 7�~�6� '��p} =�C�}p�@bŝD��FRIr��T&��RO@ \�E}��=y�OPWOYq��v0Y�SYSByU/@v�$SOPġ�d���ϪUΫ}pPR�UN����PA��Dp���rɡL�_OUo�顢q�$)�I�MAG��w��0Pf_qIM��L�INv��K�RGOVRDt��X�(�P*�J�|��0L_�`]��0�SRB1�0��M�񦷺ED}��p ��N��PMֲ���c�w�S�L�`q�w x �$OVSL4vSDI��DEX��Đ�#���-�V} *�N 4�\#�B�2�G�B�_ЅM���q�E� �x Hw��p��AWTUSW���C�08o�s���BTM�ǌ�I�k�4��x�԰.q�y Dw�E&�����@E�r��7��ж���EXE��ἱ��p���f q�z @w�f��UP'��$�pQ�XN����������� �PG΅{ h $SUB�����0_���!�MP�WAIv�P7ã�L�OR���F\p˕$�RCVFAIL_9C���BWD΁�v�DEFSP!p | Lw���Я�8\���UNI+������H�R�+�}_L�\pP��x�t���p�} H�> �*�j�(�s`~��N�`KETB�%�RJ�PE Ѓ~��J0SIZE\���X�'�ڡ�S�OR��FORMAT�`��c �,��WrEM�t��%��UX��G��PLI���p�  $>ˀP_SWI�pq��J_PL��AL_� �����A��BԺ�� C��D�$mE��.�C_��U�� � � 1���*�J3K0��^��TIA4��5��6��MOM�����П���ˀB��AD`����������PU� NR��������m��� A$PI�6q��	��� ��K4�)6�U��w|`��SPEEDgPG��������Ի� 4T�� � @��SAMr`��\�]��MOV_�_$�@npt5��5���1���2��������'�2S�Hp�IN�'� @�+����4($<4+T+GAMMWf�1>'�$GET`�p����Da���

pLI�BR>�II2�$H�I=�_g�t��2�&E�;��(A�.� �&LW �-6<�)56�&]��v��p��V��$�PDCK���q��_?�����q�&����7��4���9+� ��$IM_SR��pD�s�rF��r�rL	E���Om0H]��0�-�pq��P~JqUR_SCRN��FA���S_SAV�E_D��dE@�NOa�CAA�b�d@�$q� Z�Iǡs	�I� �J�K � ����H�L��> �"hq������ɢ �� bW^US�A�-M4���a�� )q`��3�WW�I@v�_��q�.MUAo�� �� $PY+�3$W�P�vNG�{� �P:��RA��RH��RO�PL�����q� ��sJ'�X;�OI�&�Zxe8 ���m�� p��ˀ�3s�O�O�O�O�Ot�aa�_т� |�� q�d@��.v��.v��d@��[wFv��E���%sÔt;B�w�|�tPn���PMA�QUa ��Q8��1�wQTH�HOLG�oQHYS��ES�F�qUE�pZB��Oτ�  ـPܐ(�AP����v�!�t�O`�q��u�"���FA��IGROG�����Q2����o�"��p��INFOҁ�׃V����R��H�OI��� (�0SLEQ����@��Y�3����Á��P�0Ow0���!E�0NU��AUT<�A�COPY�=�(/�'��@Mg�N��=��}1������ ��RG4��Á���X_�P�C$;ख�`��W���P��@�������E�XT_CYC b�HᝡRpÁ�r��_NAe!А����ROv`	�� �s ���POR_�1�E2�SRV �)l_�I�DI��T_� k�}�'���dЇ�����U5��6��7��8i��H�SdB���2�$R��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,�0FL`�o@SYN��K�M��Ck��PWR+�9ᘐ���DELA}�dY֟pAD�a"�QSwKIP4� �A�Z$�OB`NT����P_$�M�ƷF@\b Ipݷ�ݷ�ݷd�� ��빸��Š�Ҡ��ߠ�9��J2R�� ��� 4V�EX� TQQ����TQ������� ��`�#�RD�C�V� �`��X)�R�p�����r��~m$RGEAR_� sIOBT�2FLG��LfipER�DTC����Ԍ���2TH2N<S}� 1���uG T\0 ���u�M\Ѫ`I�d"��REF�1Á� yl�h��ENAB��cTPE�04�]�� ��Y�]��ъQn#��*���"�������2�Қ��߼���������3�қ'�9�K�]�o��
�4�Ҝ�������(�����5�ҝ!�3��E�W�i�{��6�Ҟ��������������7�ҟ-?Qcu
�8�Ҡ����x���SMSKÁ%�l��a��EkA��oMOTE6������@�݂TQ�IO�}5�ISTPVONΜ�POW@��� �pJ����p�����E�"$DSB_SIGN�1UQ�x��C\ЖtRS232���R�iDEVI�CEUS�XRSRP�ARIT��4!OP�BIT�QI�OWCONTR+�TQ���?SRCU� MpSU_XTASK�3N�p��0p$TATU�P�E#�0�����p_�XPC)�$FRE?EFROMS	pna��GET�0��UP%D�A�2E#P� :�ߧ� !$USAN�na&�����ERI�0�RpRY$q5*"_j@�Pm1�!N�6WRK9KD����6��QFRIEND�Q�RUFg�҃�0oTOOL�6MY�t�$LENGTHw_VT\�FIR�p�C�@ˀE> +IUF�IN-RM��RGyI�1ÐAITI�b$GXñ3IvFG2v7�G1���p3�B�GP1R�p�1F�O_n 0��!RE��p�53҅�U�TC��3A�A�F ��G(��":��� e1n!��J�8�%���%�]��%�� 74�XS O0�L��T�3�H&��8���%b453G�E�W�0�WsR�TD ����T��M����Q�T�]�$V 2�����1�а91�8�02*�;2k3�;3�:i fa�9-i�aQ��NS���ZR$V��2BVwEVP�	V�B;�����& �S�`��F�"�k�@�2�a�PS�E �$pr1C��_$Aܠ�6wPR��7vMU�cS��t '�/89�� 0�G�aV`��p�d`����50�@��-�
25S^�� ��aRW�����B�&�N�A)X�!�A:@LAh�^�rTHIC�1I�8��X�d1TFEj��q>�uIF_CH�3�qaI܇7�Q�pG1Rx�V���]��:�u�_�JF~�PRԀƱ��RVAT��� ���`���0RҦ�DO�fE��COUԱ��A�XI���OFFS=E׆TRIGNS����c����h�����Hx�Y��IGMA0�PA�pJ�E�ORG�_UNEV�J� ��S�����d ӎ$CА�J�GR3OU����TOށ�!DSP��JOG�Ӑ�#��_Pӱ�"O��q����@�&KEPF�IR��ܔ�@M}R&��AP�Q^�Eh0��K�SYS�q"K�;PG2�BRK�B��߄�pY�=�d�����`AD_�����BS�OC���N��DU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR-���C��ˢΓ�OR٧3N]0ڦF��ڦ��OV��SF��p���F+�r!���CC��1q"LCHD}L��RECOVʤc0��Wq@M������#RO�#��Ȑ_+���� @0�e@VER��$OFSe@CV/ �2WD�}���Z2���TR�!|���E_FDO��MB_CM���B��BL�bܒ#��adt�VQR�$0p���G$�7�AM5��� e����_M;��"'����8$CA��'�E�>8�8$HBK(1���IO<�����QPPA������
���������DVC_DBhC;��#"<Ѝ�r!"S�1[ڤ�S�3[֪�/ATIOq 1q� �ʡU�3���CAB Ő�2�CvP��9P^�B��_� �SUBCPU�ƐS�P � M�)0NS�cM�"r�?$HW_C��U���S@��SA�A�pl$�UNITm�l_�A�T���e�ƐCYC=Lq�NECA����FLTR_2_F�IO�7(��)&B�LPxқ/�.�_SCT�CF_`�Fb�l���|��FS(!E�e�CHA��1��4�D°"3�RS�D��$"}����_Tb�PRO����� KEMi_��a�8!�a !�a��D�IR0�RAILAiCI�)RMr�LO��C���Qq��#q��V��PR=�S�A�C/�c 	��FUsNCq�0rRINP`�Q�0��2�!RAC �B ��[���[gWARn���BL�A�q�A����D�Ak�\���LD@0���Q��qeq�TI"r��K�hPgRIA�!r"AF��Pz!=�;��?,`�R�K���MǀI�!�D�F_@B�%1n�LM��FAq@HRDY4�4_�P@RS�A�0|� �MULSE@x���a ���ưt��m�$�1-$�1$1o������ x*�EaG"p����!AR���Ӧ�09�2,%� 7�wAXE��ROB���WpA��_l-��SY�[�W!‎&S�'WR�U�/-1��@�STRП�����Eb� !	�%��J��AB� ����&9�����OTo0v 	$��ARY�s�#2��Ԓ�	ёFI�@��$LINK(|�qC1�a_�#����%kqj2XYZ@��t;rq�3�C1j2J^8'0B��'�40����+ �3FI���7`�q����'��_Jˑp���O3�QOP_�$2;5���ATBA�2QBC��&�DUβ�&=6��TURN߁"r��E11:�p��9GFL��`_���* �@�5�*7���Ʊ 1�� KŐM��&8���"r��ORQ��a �(@#p=�j�g�#qXUp�����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb��T {�, ��@;�uQ���P \�i��UuQ�We�eL�SERʑe	��!E� O���UdAas���4S�/7����AX��B�'q��E1�e ��i��irp�jJ@�j �@�j�@�jP�j@ �j �!�f��i��i��i ��i��i�y�y��'y�7yTqHyDEBU8�$32����qͲf2G + AB�����رnSVS�7� 
#�d��L�#�L� �1W��1W�JAW��AW� �AW�QW�@!E@?\D2�3LAB�29U�4�Aӏ��C  �o�ERf�5� �� $�@_ A��!�PO��à�0#��
�_MRAt�� �d � T��ٔEcRR����;TY&����I��V�0�cz�TOQ�d�PL[ �d�"ҍ�	��C! � pp`T)0���_V1Vr�aӔ�����2ٛ2�E����@�8H�E���$W���j��V!��$�P@��o�cI��aΣ	 �HELL_CFG�!� 5��Bo_BASq�SR3�\�� a#Sb�T��1�%��2��U3��4��5��6��e7��8���RO�����I0�0NL�\CAqB+�����ACK4� ����,�\@2@�&�?�7_PU�CO. U�OUG�P~ ����m�ذ�����TPհ_KcAR�l�_�RE*��P���|�QUE����uP����CST?OPI_AL7�l��k0��h��]�l0SE�M�4�(�M4�6�T�YN�SO���DI�Z�~�A�����m_T}M�MANRQ���k0E����$KEYSWITCH��ص�m���HE��BE�AT��|�E- LE(~�����U��F!Ĳ�|��B�O_HOM=�OGREFUPPR�&��y!� [�C��O��-ECOC��Ԯ0_IOCMWD
�a���(k��� �# Dh1���UX����M�βgPgCFOR�C�����OM.  �� @�5(�U��#P, 1��, 3���45	�NPXw_ASt�� 0���ADD���$S�IZ��$VAR\���TIP/�.�
�A�ҹM�ǐ��/�H1�+ U"S�U!Cz����FRIF��J�S0���5Ԓ�NF��܍� � xp`SIƗ�TE�C���CSG%L��TQ2�@&���x�� ��STMT��2,�P �&BWuP���SHOW4���S�V�$�� �Q�A00�@Ma}����� �����&���5���6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G�� 0G���0G���@GP��PG��1	1	U1	1+	18	1E	U2��2��2��2��U2��2��2��2��U2��2��2	2	U2	2+	28	2E	U3��3��3��3��U3��3��3��3��U3��3��3	3	U3	3+	38	3E	U4�4��4��4��U4��4��4��4��U4��4��4	4	U4	4+	48	4E	U5�5��5��5��U5��5��5��5��U5��5��5	5	U5	5+	58	5E	U6�6��6��6��U6��6��6��6��U6��6��6	6	U6	6+	68	6E	U7�7��7��7��U7��7��7��7��U7��7��7	7	U7	7+	78	7Ev��VP��UPDs��  �`NЦ��5�YSLOt�� � L��d���A熜aTA�0d��|�AcLU:ed�~�CUѰzjgF!aID_L��֑eHI�jI��$F�ILE_���d���$2�fSA>�� �hO��`E_BLC�K��b$��hD_CPUyM�yA��c�o��d��Y����R ��Đ
PW��!� -oqLA��S=�ts�q~tRUN�qst �q~t���qst�q~tw �T��ACCs��X -$�qLEN;��tH��ph��_�I��ǀLOW_7AXI�F1�q�d2*�MZ���ă��W��Im�ւ�aR�TOR���pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v��������TCV��؁��T ��ي�����t�V��$��V�Jj�R�MA����J��m�u�b����q2j�#�U�{�t�K�JK��VK;���H����3��J0����J�J��JJ��AAL���ڐ��ڐԖ4Օ5���N1���ʋƀJW�LP�_(�g�,��pr�� `�`GGROUw`��B�ПNFLIC��f�R�EQUIRE3�E�BU��qB���w�2�����p���q5�p��� \��APPRҒ�C}�Y�
ްEN�٨CLO7��S_!M��H���u�
�qu�o� ���MC��8���9�_MG��C��Co��`M�в�N�B;RKL�NOL|�N�:[�R��_LINђ�$|�=�J����Pܔ�� ���������������6ɵ�̲8k�+��q>���� ��
���q)��7�PATH3�L�B�L��H�w�ڡ��J�CN�CA��Ғ�ڢB�IN�rU�CV�4a��C!�UMB��Y,���aE�p�����ʴ���PAYwLOA��J2L`OR_AN�q�Lpp����$�M�R_F�2LSHR��N�L�Oԡ�Rׯ�`ׯ�ACRL_G�ŒЛ�� ��Hj`߂$H�M���FLEXܣ��qJ�u� : �������������1�F1�V�j�@�R�d�v�������E ����ȏڏ����"� 4�q���6�M���~�� U�g�y�ယT��o�X��H������藕? �����ǟِݕ�ԕ ����%�7��P��J�� � V�h�z����`AT�採@�EML�� S��J|��Ŝ�JEy�CTR,��~�TN��FQ��HAND_VB-�q��v`�� $���F2M����ebSW��q�'��� '$$MF�:�Rg�(@x�,4�%��0&A�` �=��aM)F�AW�Z`
i�Aw�A��X X�'p�i�Dw�D��Pf�G�p�)STk��!x��!N��DY�pנM�9$ `%Ц�H��H�c�� ����0� ��Pѵڵ����������J��� ���1��Rx�6��QASYMv�����v��J���c���_SH>��ǺĤ��ED����������J��İ%��C�IDِ�_�VI�!X�2PV_UNIX�FThP�J��_R�5_Rc�cTz� pT�V��@���İ�߷�$�U ��������Hqpˢ��aE�N�3�DI����Op4d�`J�� x 
g"IJAA�az�aabp��coc�`a�pdq�a�{ ��OMME��� �b�RqAT(`P�T�@� S��a7�;� Ƞ�@�h�a�iT�@<�� $DUMM�Y9Q�$PS_6��RFC�  S�v� � ���Pa�c XƠ���STE����SBRY�M2�1_VF�8$SV_ERF�O��LsdsWCLRJtA��Odb�`O�p � �D $GLOBj�_LO���u�q�cpAp�r�@aSYS�q�ADR``�`TC}H  � ,��ɩb�W_NA��a�7���SR��?�l ��� 
*?�&Q�0"?�;'?� I)?�Y)��X���h��� x������)��Ռ�Ӷ� ;��Ív�?��O�O�O|�D�XSCRE�j�p����ST�F�s}y`�����/_HA�q� TơgpTYP�b����G�aG���Od0IS_䓀d�;UEMd� ����p�pS�qaRSM_��q*eUNEXCE1P)fW�`S_}pMрx���g�z�����ӑC�OU��S�Ԕ 1-�!�UE&��Ubwr���PROGM�F�L@$CUgpP�O�Q��5�I_�`H>� � 8�� �_HE�PS�#��`?RY ?�qp�b���dp�OUS>�� � @6p�v�$BUTTp�R|pR�COLUMq�<e��SERV5��PANEH�q� w� �@GEU��Fy��)$HE�LPõ)BETERv�)ෆ���A  � ��0��0��0�ҰIN簪c�@N(��IH�1��_�o ֪�LN�r'� �qpձ_ò=��$H��TEX8l����FLA@��/RELV��D`���������M��?,@�ű�m����"�USRVIEW�q�� <6p�`U�`��NFI@;�FOsCU��;�PRI@�m�`�QY�TRI}P�qm�UN<`�Md� #@p�*eW�ARN)e6�SRT+OL%��g��ᴰ�ONCORN��RA�U����T���w�V�IN�Le� =$גPATH9�ג�CACH��LOG�!�LIMKR���x�v���HOST��!�b�R��OgBOT�d�IM>�	 �� ���Zq��Zq;�VCPU_�AVAIL�!�EX	�!AN���q�`�1r��1r��1 ��\��p�  #`C�����@$TOOLz�$��_JMP�� ���e$S�S����VSHI9F��Nc�P�`ג��E�ȐR����OS�UR��Wk`RADILѮ��_�a��:�`9a��`a�r��LULQ�$OUTPUTg_BM����IM��AB �@�rTILNSCO��C7� ������&�� 3��A���q���$m�I�2G�ϑV�pLe9�}��yDJU��N��WAIT֖�h}��{�%! NE�u��YBO�� �� $`�t��SB@TPE��NECp�J^FY�nB_T��R�І�a�$�[YĭcB��dM ���F� �p�$�pvb�OP?�MAS�W_DO�!QT�p�D��ˑ#%��p!"D�ELAY�:`7"JOY�@(�nCE$���3@ �xm��d�pY_ [�!"�`�"��[���P�? ϑZAB�C%��  $��"R��
ϐ�$$�CLAS�������!pϐ� � V�IRT]��/ 0AB�S����1 5�� < �!F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZi{0-�AXL�p��"��63  �{tIN8��qztPRE�����v�p�uLARM�RECOV �9�rwtNG�� �.;	 A   ��.�0PPLIC���?5�p��HandlingTool o�� 
V7.50�P/23-�  ��PB��
��_�SWt� UP�!� x�F0��t����Aϐv� 8[64�� �it��y� N2 �7DA5�� �j� QBy@��o�Noneis�ͅ˰ ��T��]�!LAA+x>�_l�V�uT�:�s9�UTO�"����t�y��HGAPO�N
0g�1��Uh�D� 1581�����̟ޟry����Q 1���p� ,�蘦���;�@��q�_��"�" �3c�.�H����D�HTTHKY X��"�-�?�Q���ɯ ۯ5����#�A�G�Y� k�}�������ſ׿1� ����=�C�U�g�y� �ϝϯ�����-���	� �9�?�Q�c�u߇ߙ� �߽���)�����5� ;�M�_�q����� ��%�����1�7�I� [�m����������! ����-3EWi {������ )/ASew� ���/��/%/ +/=/O/a/s/�/�/�/ �/?�/�/?!?'?9? K?]?o?�?�?�?�?O��?�?�?O#O]���T�O�E�W�DO_C�LEAN��7��CN�M  � ��__/_A_S_�D?SPDRYR�O��HIc��M@�O�_�_ �_�_oo+o=oOoao�so�o�o���pB��v �u���aX�t����|��9�PLUGG����G��U�PRCvPB��@��_�orOxr_7�SEGF}�K[mwxq�O�O������?rqLAP �_�~q�[�m������ ��Ǐُ����!�3�>x�TOTAL�f y�x�USENU�p©� �H���B��RG�_STRING �1u�
��Mn�S5�
ȑ_�ITEM1Җ  n5�� ��$�6�H� Z�l�~�������Ưد����� �2�D��I/O SIGN�AL̕Try�out Mode�ӕInp��Simulatedב�Out��O�VERR�P = �100֒In �cycl��בP�rog Abor���ב��Stat�usՓ	Hear�tbeatїM?H Faul��Aler'�W�E�W� i�{ύϟϱ������� �CΛ�A���� 8�J�\�n߀ߒߤ߶� ���������"�4�F�pX�j�|���WOR{p Λ��(ߎ����� �� $�6�H�Z�l�~����� ���������� 2PƠ�X ��A {������� /ASew������SDEV [�o�#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y?PALTݠ1�� z?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O��O�O�O_�?GRI �`ΛDQ�?_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|�� �������0�xB�T��oPREG�> �� f���Ə؏��� � �2�D�V�h�z��������ԟ���Z���$ARG_��D �?	���;���  w	$Z�	[O��]O��Z�p�.�SB�N_CONFIG� ;��������CII_SAV/E  Z������.�TCELLSE�TUP ;�%�HOME_IO�Z�Z�%MOV_8��
�REP�lU��(�UTOBACK�ܠ��F�RA:\z� X\�z�Ǡ'`�z����ǡi�INI�0�z���n�MESSAG���ǡC���ODE_D�������%�O�4�n�PAU�SX!�;� ((O>��ϞˈϾ� �����������*� `�N߄�rߨ߶�g�l ?TSK  wͥ�<_�q�UPDT+���d!�A�WSM_kCF��;���|'�-�GRP 2:�V?� N�BŰA�߾%�XSCRD1�1�
7� �ĥĢ ����������*��� ����r����������� 7���[�&8J\�n��*�t�GRO�UN�UϩUP_kNA�:�	t�n�_ED�17��
 �%-BCKEDT-�2�'K�`ܵu��z�q�q�z����2t1������q�k�(/��ED3/��/�.a/�/;/M/ED4�/t/)?��/.?p?�/�/ED5`??�?<?.�?O�?�?ED6O�?qO��?.MO�O'O9OED7�O`O_�O.�O\_�O�OED8L_,�_�^-�_ oo_�_�ED9�_�_]o�_	`-9o�oo%oCR _ 9]�oF�o�k�� � NO_DEL���GE_UNU�SE��LAL_?OUT �����WD_ABOR�ﰨ~��pITR_�RTN��|NO�NSk���˥C�AM_PARAM� 1;�!�
 8�
SONY X�C-56 234�567890 �ਡ@���?}��( А\��
���{����^�H�R5q�̹��ŏR5y7ڏ�Aff���KOWA SC�310M
�x��>��d @<�
� ��e�^��П\�� ��*�<��`�r�g��CE_RIA_I��!�=�F���}�z� ��_LeIU�]������<��FB�GP 1.��Ǯ�M�x_�q�0�C*  ��V��C1��9��@��iG���CR�C]��Ud��l��s��R��T���[Դm��v���������� C����(�����=�{HE�`ONFIǰ��B�G_PRI 1�{V���ߖπ�Ϻ����������C�HKPAUS�� ;1K� ,!uD� V�@�z�dߞ߈ߚ��� �������.��R�<�hb���O���������_MOR��� �6��� 	 �����*��N�<��������?��q?$;�;����K��9��P���çaÃ-:���	�

 ��M���pU�ð��<���,~��DB����튒)
mc:c?pmidbg�fF�:���s��p�|/�  �Q��	� �s>��3Q�?�����Yg�/�م�Xf�M/w�O/�
D�EF l��s)��< buf.t�xts/�t/��ާ��)�	`�����=�L���*MC��1�����?43��1���t�īCz � BHH�>'��B�$�9G�<�5@@�C�����1Y
K�@�D���;A�e8��.D�� �1��=B��IE�C�e=�D�<�X�F���1Y	��,�'w�1���s�U��.�p�����1�BDw�M@x8�K��CҨ����g@D��p@�0EYK�EX��EQ�EJ�P F�E�F�� G��=F�^F E�� F�B� H,- Ge��H3Y��:��  >�33 ����~  n48�~@��5Y�E>��ðA��Y<#�
�"Q ���+_�'R_SMOFS�p�.�8��)T1��DE 3��F 
Q��;;�(P  B_<_���R����	op6C�4P�Y
s@ ]A(Q�2s@C�0B3�Ma�C{@@*cw��UT��pFPROG !%�z�o�oigI�q����v��ldKEY_TOBL  �&S�#�� �	
��� !"#$%&'�()*+,-./�01i�:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�����������������������p`LCK�l4�p`�`STAT� ��S_AUTO_�DO���5�IN?DT_ENB!���1R�Q?�1�T2}�^��STOPb���TR�Lr`LETE���Ċ_SCREEN� �Zkc�sc��U��MME�NU 1 �Y  <�l�oR�Y 1�[���v�m���̟�� ���ٟ�8��!�G� ��W�i��������ï կ��4���j�A�S� ��w�����迿�ѿ� ���T�+�=�cϜ�s� ���ϩϻ������� P�'�9߆�]�o߼ߓ� ���������:��#� p�G�Y������� ����$����3�l�C� U���y������������ ��	VY)�_M�ANUAL��t�DwBCO[�RIG>�DBNUM� ���B1 e
�PXW�ORK 1!�[ �_U/4FX�__AWAY�i�/GCP  b=�Pj�_AL� #�j�Yи�܅ `�_�  1}"�[ , 
�@mg�&/~&lMZ��IdPx@P@#ON�TIMه� dɼ`&�
�e�MO�TNEND�o�R�ECORD 1(��[g2�/{�O� �!�/ky"?4?F?X? �(`?�?�/�??�?�? �?�?�?)O�?MO�?qO �O�O�OBO�O:O�O^O _%_7_I_�Om_�O�_  _�_�_�_�_Z_o~_ 3o�_Woio{o�o�_�o  o�oDo�o/�o S�oL�o���� @���+�yV,� c�u��������Ϗ>� P�����;�&���q� ��򏧟��P�ȟ�^� �����I�[�����  ���$�6��������jTOLEREN�CwB���L��͖ CS_CFG� )�/'d�MC:\U�L%0?4d.CSV�� �c��/#A ��CH
��z� //.ɿ���(S�RC_OUT *��1/V�?SGN +��"���#�28-J�AN-20 15�:20027l�2�1:48+ P;��ɞ�/.���f�pa�m���PJPѲ��V�ERSION �Y�V2.0�.�ƲEFLOG�IC 1,� 	:ޠ=�ޠL���PROG_ENqB��"p�ULSk'� ����_WRS�TJNK ��"fE�MO_OPT_S�L ?	�#
 	R575/# =�����0�B����TO  �ݵϗ��V_F EX�d��%��PATH ;AY�A\����\�5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAqU��z�^"MSWX��.�<�4,#�Y�/�
!J�6%Z�I~m��$SBL__FAUL(�0�^9'TDIA[�1<��<� ���1�234567890
��P��HZ l~������ �/ /2/D/V/h/�Z� P� ѩ� yƽ/��6�/�/�/? ?/?A?S?e?w?�?�?��?�?�?�?�?�,/�U3MP���� �A�TR���1OC@PM�El�OOY_TEM=P?�È�3F���G�|DUNI��.�Y�N_BRK 2�_�/�EMGDI_�STA��]��ENC�2_SCR 3�K7(_:_L_^_l& _�_�_�_�_)��C�A14_�/oo/oAo�Ԣ�B�T5�K� ϋo~ol�{_�o�o�o '9K]o� �������� #�5��/V�h�z��л` ~�����ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T���x��������� ү�����,�>�P� b�t���������ο� ���(�f�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������:� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ���*<N` r������� &8J\n� ���������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?��?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O��O__NoETMO�DE 16�5��Q �d�X
�X_j_|Q�PRROR�_PROG %fGZ%�@��_  �U�TABLE  �G[�?oo)oRjR�RSEV_NUM�  �`WP��QQY`�Q_AUT�O_ENB  ��eOS�T_NOna �7G[�QXb W *��`��`��`	��`d`+�`�o�o�o�dHISUc�QOP�k_ALM 18G[� �A��l�P+�ok}����r�o_Nb�`  G[��a�R
�:PTCP_VER !GZ�!�_�$EXTL�OG_REQv9�i\�SIZe�W��TOL  �QD�zr�A W�_BWD�p��xf́t�w_DI�� 9�5��d�T�QsRֆS�TEP��:P�O/P_DOv�f�P�FACTORY_�TUNwdM�EATURE :�5�̀rQHa�ndlingTo�ol �� \sf�mEngli�sh Dicti�onary��ro�duAA V�is�� Mast�er����
EN�̐nalog I�/O����g.fd�̐uto Sof�tware Up�date  F �OR�matic Backup���H596,�g�round Ed�itޒ  1 H�5Camer�a�F��OPLG�X�ell𜩐II�) X�ommՐs�hw���com��c9o���\tp����pane��  o�pl��tyle �select��a�l C��nJ�Ցo�nitor��RD�E��tr��ReOliab𠧒6U�Diagnos(��푥�5528�u���heck Sa�fety UIF���Enhance�d Rob Se�rv%�q ) "�S�r�User F�r[�����a��xt�. DIO �f�iG� sŢ��en]dx�Err�LF�� pȐĳr됮� ܻ���  !��FCTN Menu`��v-�ݡ���TP �Inېfac� � ER JG�C�pבk Exczt�g��H558��igh-Spex��Ski1�  2�
P��?���mmuwnic'�ons���&�l�ur�ې��S�T Ǡ��con�n��2��TXPL��ncr�str�u����"FAT�KAREL C�md. LE�ua�G�545\��Ru�n-Ti��Env��d
!���ؠu++�s)�S/W���[�Licen3seZ��� 4T�0��ogBook(S�yڐm)��H54�O�MACROs,~\�/Offse��7Loa�MH�������r, k�Mec�hStop Pr�ot���� lic�/�MiвShif8����ɒMixx���)���xSPS�Mo�de Switc�h�� R5W�Mo��:�.�� 74 H���g��K�2h�?ulti-T=�M����LN (P{os�Regiڑ�������d�ݐt Fun�ǩ�.������Num~����� l�ne��ᝰ Ad�jup�����  �- W��tatu�w᧒T�RD�Mz�ot��sco+ve U�9����3Ѓ�uest 492�*�o������62;�SNPX yb ���8 J7`���Libr��J�48���ӗ� �Ԅ�
��6O�� Part�s in VCCMt�32���	�{�ޤ�J990��/I�� 2 P��TM/ILIB��H���P�AccD�L�7
TE$TX�ۨ�7ap1S�Te����pkey��wգ��d��Unex�ceptx�mot�nZ���������є�� O���� �90J�єSP CSXC<�f��Ҟ�� Py�We}���P3RI�>vr�t��men�� ��iPɰa�����v�Grid�pla�y��v��0�)�H1��M-10iA(_B201 �2\�� 0\k/�Ascii�l�Т�ɐ/��Col��ԑGuaMr� 
�� /P-��ޠ"K��st{P�at ��!S�Cyqc�҂�orie�v�IF8�ata- quҐ�� ƶ��moH574��RL���am���Pb�HM/I De3�(b����PCϺ�Pas�swo+!��"PE�? Sp$�[���tp\��� ven��Tw��N�p�YELLO�W BOE	k$Ar�c��vis��3�*�n0WeldW�cGial�7�V#tѓOp����1y� �2F�a�portN�(�p�T1�T� ��� ��xy]�&T5X��tw�igj�1�� b� ct\�J�PN ARCPS�U PR��oݲO�L� Sup�2fi�l� &PAɰאcr=o�� "PM(�����O$SS� eвtex�� r���=�=t�ssagT��	P��P@�Ȱ�锱�rtW��H'>r��dpn��n1
�t�!� z ��as�cbin4psy�n��+Aj�M H�EL�NCL V�IS PKGS �PLOA`�MB ��,�4VW�RI�PE GET_V�AR FIE 3�\t��FL[�OO�L: ADD R�729.FD \Kj8'�CsQ�QE���DVvQ�sQNO �WTWTE��}PD�  �^��biRFwOR ��ECTn��`��ALSE A�LAfPCPMO-�130  M" �#h�D: HAN?G FROMmP��AQfr��R709� DRAM AV�AILCHECK�SO!��sQVPCS� SU�@LIMC�HK Q +P~dFF� POS��F�Q �R5938-12 CHARY��0�PROGRA �W�SAVEN`A�ME�P.SV��7��$En*��p?FU��{�TRC|� SH�ADV0UPDAT� KCJўRSTA�TI�`�P MUC�H y�1��IMQ� MOTN-00�3��}�ROBOG�UIDE DAU�GH�a���*�toQu����I� Šhd��ATH�PepMOV�ET�ǔVMXP�ACK MAY ?ASSERT�D���YCLfqTA�rB�E COR vr�*Q3rAN�pRC OPTIONSJ1�vr̐PSH-1k71Z@x�tcǠSU1�1Hp^9R!�Q�`C_T�P��'�j��d{tby app wa 5I�~d�P�HI���p�aTEL��MXSPD TIB5bLu 1��UB6@��qENJ`CE2�6�1��p��s	�ma�y n�0� R6�{�R� �Rtraf�f)�� 40*�p���fr��sysv�ar scr Jq7��cj`DJU���bH V��Q/�PS?ET ERR`J`� 68��PNDA�NT SCREEN UNREA��4'�J`D�pPA���p=R`IO 1���P�FI�pB�pGROUN�PD��G��R�P|�QnRSVIP !p��a�PDIGIT �VERS�r}BLo��UEWϕ P06s  �!��MAGp0�abZV�DI�`� SSUE�ܰ��EPLAN JO�T` DEL�pݡ#�Z�@D͐CALLOb�Q ph��R�Q�IPND��IMGޏR719��MN�T/�PES �pV:L�c��Hol�0Cq����tPG:�`C�M��canΠ��pg�.v�S: 3D �mK�view d2�` �p��ea7У�b� of �Py����ANNOT AC?CESS M��Ɓ�*�t4s a��lyok��Flex/�:�Rw!mo?�P�A?�-�����`n�p�a SNBPJ AUTO-�06f����TB��PIABL�E1q 636��P�LN: RG$�pl�;pNWFMDB�V�I���tWIT 9tx�0@o��Qui#0|�ҺPN RRS?p�USB�� t &� remov�@ �)�_��&AxEPFT�_=� 7<`�pP:��OS-144 ���h s�g��@O�ST� � CRASH DU 9���$P�pW� .}$��LOGIN���8&�J��6b046� issue 6� Jg��: Sl�ow �st��c (Hos`�c��z�`IL`IMPRWtSPOT:Wh:0\�T�STYW ./ЏVMGR�h�T0C�AT��hos��EP�q��� �O�S�:+pRTU' k�-�S� ����E:��ppv@�2�� t\hߐr��m ��all���0�  $�H� WA�͐��3 CNT0s T�� WroU�alarm���0s�d � �0SE1���r: R{�OMEBp����K� 55��RE�àSEst��g  �   �KAN�JI�no���I�NISITALI1Z-p�dn1weρ<�6�dr�� lx`��SCII L�f�ails w�� <��`�YSTEa���8o��Pv� IIH����1W�Gro>Pm 7ol\wpSh@�P���Ϡn cflx�L@АWRI �OF� Lq��p?�F�u�p��de-rel}a�d "APo �SY�ch�Abet�we:0IND t0$gbDO���r�y `�GigE�#�operabilf  PAbHi�H`���c�lead�\e�tf�Ps�r�OS� 030�&: fig��GLA )P ���i��7Np tps�wx�B��If�g�������5aE�a EXCE#dU�_�tP�CLOS��"ro�b�NTdpFaU�c�!���PNIO_ V750�Q1�8�Qa��DB ��P� M�+P�QED�D�ET��-� \rk~��ONLINEhSBUGIQ ߔĠi`�Z�IB�S apA�BC JARKY�Fq� ���0MILT�`� R�pNД �p�0GAR��D*pR8��P�"! jK�0c�T�P�Hl#n�a�Z�E V�� TASK�$VP2(�4`
��!�$�P�`WIBP�K05�!FȐB/���BUSY RUNN�� "�򁐈�2�R-p�LO�N�wDIVY�CUL���fsfoaBW �p���30	V���ˠIT`�a505�.�@OF�UNE�X�P1b�af�@�E���SVEMG� N�MLq� D0pCC_SAFEX 0c�0u8"qD �PET�`9N@�#J87����RsP�A'�M�K��`K�H GUN�CHG۔MECH��pMc� T�  y�, g@�$ ORY LEAKA�;��ޢSPEm�Ja��V�tGRIܱ�@�oCTLN�TRk��FpepR�j50�E�N-`IN�����p `�`�Ǒk!��T3/d\qo�STO�0A�#
�L�p �0�@�Q��АY�&�;pb1TO8pP�s���FB�@YpL`�`DU��aO�sHupk�t4 � P�F� �Bnf�Q�PSVG�N-1��V�SRS	R)J�UP�a2�Qx�#D�q l O��~�QBRKCTR5� ��|"-�r�<pc�j!�INVP�D ZO�� ��T`h#�Q�cHs�et,|D��"DU�AL� w�2*BRV�O117 A]�T�Nѫt�+bTa247`3��q.?��sAUz��i�B�comple�te��604.�� -�`hancZ�U� F��e8�'�  ��npJtPd!�q��`��� 5h596p�!5d�� "p �P�P�Q�0�P2�p�A�� xP��R(}\xPeJ� aʰI���E���1��p� j  �� xSP��^P �A�ApxP�q 5 sig��a��"AC;a��p
�bCexPb_p���.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o�dxPX�b]o2�� �cb�c��ixP�jupfrmp�dxP�o�`exe�ax�oFdxPtped}o���u`�cptlibxzxP�lcr�xrxP�\�blsazEdxP_fm�}gcxP�x���o�|sp�o�mc(��ob_jzop�u6�wQf��t��wms�1q���sld�)��jmc�o\�n��nuhЕ��|cst�e��>�pl�q�p�iwck���uv�f0uߒ��lvisyn�CgaculwQ�
E F  ! �Fc.fd�Qv�� �qw���Data Acquisi���nF�|1�RR631�`��TR�QDMCM� �2�P75H�1��P583xP1��7�1��59`�5�P5�7<PxP�Q����(0���Q��o pxP!/daq\�oA���@�� ge/�etd�ms�"DMER"؟,�pgdD���.��m���-��qaq.<᡾xPmo��h����f{�u�`13��MA�CROs, Sk�saff�@z����03��SR�Q(��Q6��1"�Q9ӡ�R�ZSh��P^xPJ643�@7ؠ�6�P�@�PRS�@����e �Q�UС PI�K�Q52 PTLqC�W��xP3 (��p/O��!�Pn ��xP5��03\s�fmnmc "M�NMCq�<��Q��\$AcX�FM���ci ,Ҥ�X����cdpq+�6
�sk�SK�xP�SH560,P���,�y�refp "GREFp�d�A�jxP6	�of�OFc�<g6y�to�TO_���<�ٺ���+je|�u��caxis2��xPE�\�e�q"IS�DTc��]�prax ��MN��u�b�isde܃h�\��w�xP! isba�sic��B� P�]��QAxes�R�6������.�(Ba�Q�ess��xP����2�D�@�z�atis���(�{����h��~��m��FMc��u�{�
ѩ�MNIS ��ݝ����x����xٺ��x� j75���Devic�� Interfac�R<ȔQJ754��� xP�Ne`��xP��ϐ2�б����d=n� "DNE���~
tpdnui5cUI��ݝ	bd�b�P�q_rsof�Ob
dv_ar�o��u�����stchkc��z	 8�(}onl��G!ffL+H�J(��"l"/�n�b���z�hamp��T�C2�!i�a"�59��S�q��0 (�+P�o��u�!2��xpc_2p�cchm��CHMqP_�|8бpevwsp��2쳌pcsF���#C SenxPa�cro�U·�-�R6�Pd�xPk�����p���gT�L��1d M �2`��8�1c4ԡ�3v qem��GEM,�\i(��Dgesnd��5���H{�}Ha�@s1y���c�Isu�xD��Fmd��I��7�4����u���AccuC�al�P�4� ��ɢ7TޠB0��6+6f�6��99\aFF q�SA(�U��2�
X�p�!�Bd��cb_�SaU=L��  �� ?��ܖto��otplus\tsrnغ(�qb�Wp��t���1���Tool (N. A.)�[K�7�Z�(P�m����bdfcls� k94��"K4p��qtpa=p� "PS9H�>stpswo��p�L7��t\�q���� D�yt5�4�q��w�qк�� �M�uk��rkey����s��}tҾsfeatu6�E!A��� cf)t\Xq��0���d�h5����LRC0�md�!�587���aR�(����d2V��8c?u3l\�pa3}H�&r-�Xu�b��t,�� �q "�q �Ot��~,���{�/��1c�}����y�p�r� �5���S�XAg�-�y����Wj874�-? iRVis���Queu�� Ƒ� -�6�1���(����u���tӑ����
��tpvtsn "VTSN�3C�+�� v\pRDV����*�/prdq\�Q�&�vstk=P����Ƥ�nm&_�դ�cl�rqν���get@�TX��Bd���aoQ8Ͽ�0qstr�D[�� ��t�p'Z����nqpv��@�enlIP�0��D!x�'�|���s1c ߸��tvo/�� 2�q���vb��� �q���!���h]���(� Contr{ol�PRAX�P�5��556�A@5m9�P56.@56@�5A�J69$@9�82 J552 IDVR7�hqA����16�H���La��� ��Xe�frl�parm.f�FRL�am��C9�@(F�����w6{����A��QJ643�� 50�0LSE�
_pVAR $�SGSYSC��R�S_UNITS ��P�2�4tA�TX.�$VNUM_OLD 5�1�xP{��50+�"�` Funct���5tA� }�(�`#@�`3�a0�cڂb��9���@H5נ� �P���(�A���� �۶}����ֻ}���bPRb�߶~ppr4�TPSPI�3�}�r�10�#;A� t��
`���1���96 �����%C�� Aف��=J�bIncr�	�� ��\���1o5q{ni4�MNINp	�xP�`���!��Ho�ur  r� 2�21 �?AAVM����0 ��TUP� ��J545� ��6162��VCAM  (��CLIO ��R6�N2��MSC "P ~�STYL�Cv�28~ 13\��NRE "FHR�M SCH^��DCSU%ORSsR {b�04 ��EIOC�1 �j 542 � o�s| � egis�t�����7�1~�MASK��934"7 ��O�CO ��"3�8Ļ�2���� 0 �HB��� 4�"39�N� Re�� �L�CHK
%OPLG�%��3"%MHCR&.%MC  ; 4? ���6 dPI�54��s� DSW%MDr� pQ�K!637�0Ƚ0p"�1�Р"4 ��6<27 CTNY K � 5 ���"I7��<25�%/�T�%OFRDM� �Sg!<��930 FB( �NBA�P� ( HL�B  Men�S�M$@jB( PVC ���20v��2HT�C�CTMI�L��\@PAC 116U�hAJ`SAI \@�ELN��<29s�?UECK �b�@�FRM �b�OR\���IPL��Rk0�CSXC ���V�VFnaTg@HTTsP �!26 ���G�@obIG{UI"%IPGS�r>� H863 qb�!8�07r�!34 �r�84 \so`! QLx`CC3 Fb�21��!96 rb!51� ���!53R% 1�!s3!��~�.p"9�js VATFUJ7�75"��pLR6^RP�WSMjUCTO��@xT58 F!80����1XY ta3!7�70 ��885&�UOL  GTSo
�<{` LCM �r| gTSS�EfP6 W�>\@CPE `��0cVR� l�QNL"���@001 imrb�c3 =�b�0����0�`6 w�b-P-� R-�b8n@5EW�b9 �Ґa� ����b�`ׁ�b2 20�00��`3��`4*5�`5!�c�#$�`�7.%�`8 h60�5? U0�@B6E�"aRp7� !Pr8� t�a@�tr2 'iB/�1vp3�vp�5 Ȃtr9Σ�a4r@-p�r3 F�Ⴐr5&�re`u��r7� ��r8�U�p9 �\h738�a�R/2D7"�1f���2&�7� �3 7)iC��4>w5Ip�NOr60 C�L�1bE6N�4 I�pyL�uP0��@N�-PJ8�N�8NeN�9 H�r`��E�b7]�|���88�Вࠂ9 2��a�`0�qЂ5�%U0O97 0��@1�0����1 (�q�3 5R���0���@mpU��0�0�7*��H@(q�\P"RB6�q124�b;��@����@06� x�3 pB/x�u ��x��6 H606�a1x� ��7 6 ����p�b155 �����7jUU162� �3 g��4�*�65 2e "_��P�4U1`���B�1���`0'�174� �q��P�E186g R ��P�7 ��P�8&�3 (�9o0 B/�s191�����@202��6� 3���A�RU2x� d��2 b2h`��4�᪂2�4����19v Q�2��u2Jd�Tpt2� ��H�a�2hP�$�5���!U2�p�p
�2�p��@!5�0-@��8 @��9��TX@�� �e5N�`rb26Af�2^R��a�2Kp��1y�b5(Hp�`
�5�0@�gqGA���a52ѐ�Ḳ-6�60ہ5� ׁ�2��8�E��9�EU)5@ٰ\�q5hQ`S*�2ޖ5�p\w�۲��pJ �-P��5�p1i\t�H�4��PCH�7j��phiw�@��P��x��559 ldu� P�D���Q�@������� �`.��P>�:��8�581�"�q�58�!AM۲T�Aw iC�a589��0@�x����5 �a��12׀0.�1���,��2����,�!P\h8���Lp ��,�7��6��0840\��ANRS 0C}A��p���{��ran��FRA��Д�е�� �A%���ѹ�Ҍ��� ��(����Ќ���� ����������ь�����$�G��1��ը���������� sxS�`q�  ������`64��M��iC/50T-H��`����*��)p46���� C��N����m7;5s֐� Sp���b46��v����Г/M-71?�7�З����42������C�2��-�а�70�r�E��/h����`O$��rD���c7c7C�q��Ѕ����L��/��2\imm7c7�g������`���(��e� ����"�������a0 r��c�T,�Ѿ�"��,�� ��x�Ex�m77t����k����5�����)�iC��-HS-�  B
_�>���+�Т�7U�]���Mh7
�s��7�������-9?�/260L�_������Q��������]�9pA/ @���q�S�х����h621��c��92����8��.�)92c0�g $�@�����)$��5$���pylH"O"
��21���t?�350����p��$�0�
�� �350!����0��9�U/0\{m9��M9A3�P��4%� s��3M$���X%u���"him�98J3����� i d �"m4~�103p�� <����h794̂�&R���H�0����\� ��g�5AU��՜��0�� �*2��00��#0�6�АՃ�է!07{r ���������kЙ@����EP �#������?��#!��;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?�ҽCD25L����u0�"l�2BL
#��B��\20�2_�r �re���X��1��N����A@��z��`C��pU��`��04H��DyA�\�`fQ���sU���\�5  ��� p�g�^P��<$85��p�+P=�ab1l��G1LT��lA8�!puDnE(�20T��qJ�1 e�bH85��h�b�Ռ�5[�16B@s��������d2�8�x��m6t!`Q ����bˀ���b#�(�6iB;S�p�!��3 � ��b�s��-`Є_�W8�_����6�I	$�X5�1�U85��R�p6S����/ �/+q�!�q��`�6o���5m[o)�m6s�W��Q�?��setC06p ��3%H�5��10p$����g/��JrH��  9��A�856���d�F�� ���p/2��@h�܅�✐)�5���̑v��(��m6���Y�H�ѝ̑m�6(�Ҝ��a6�DM����#-S�+��H2��� ��Ҽ�� �r̑���✐��l���p1����F���2�\t6h T6H����� ��'Vl���ᜐ�V@7ᜐ/����;3A7��p~S��������4�`圐�V���!3��2�PM[��%�ܖO�chn��ve�l5����Vq���_a�rp#��̑�.���2l_hemq$�.�'�6415���5����?����F�����5 g�L�ј[���1���𙋹1����M7NU�М��eʾ����Euq$D;��-�4��3&H�f�c�Ĝ�h�� ����u���〜���ZS�!ܑ4���M	-����S�$̑�ք �� 0��<�����.07shJ�H�v�� ��sF��S*󜐳����̑���vl�3�A�T��#��QȚ�Te��q�p�r����T@75j�5 �dd�̑1�(UL�&�(� ,���0�\�?���̑�a��� xSP ���a�e�w�2��(�2	�2�C��A/����\�+p�����21 9(ܱ�CL S���� B̺��7F���?�<�lơ1L����c�� ���u9�0����e!/q��O���9�K��r9 (��,�Rs���ז�5�G�m20Ac��i��w�2��:�0`�$��2�2l�0�@k�X�S� ,�ι2��hO���1!41w����2T@� _std ��G�y� �ң�H� jdgm����w0\�  �1L���	�P�~� W*�b��t 5�������3�,���E {������L��5\L��3�L�|# ~���~!���4�#�� O����h�L6A�������2璥����44�����[6\j4s��·���#��ol�E"w�8Pk��� ��?0xj�H1�1Rr��>��]�2a�2AHw�P ��2��|41�8 ��ˡ��{� �%�A<��� +�?�l��0�&�"��|�`Am1�2������3�HqB�� K�R��ˑb�W���Fs ���)�ѐ�!���ah�1����5��16�16C��C����0\imBQ��d���(�b��\B5�-���DiL���O�_�<��PEtL�E�RH�ZǠP8gω�am1l��u� ��̑�b�<����<�$�T�̑�F����I ̑�Dpb��X"��hrް�p� ���^�P��9�0\� j9�71\kckrcfJ�F�s�����c��e "CTME�r����ɛ��a�`mai�n.[��g�`run}�_vc�#0�w��1Oܕ_u����bctme��Ӧ�`ܑ��j735�- K�AREL Use% {�U���J��(1���p� Ȗ�9��B@��L�9��7j�[�atk208 C"K��Kя��\��9��a��̹����c�KRC�a�o ��kc�qJ�&s�����Gr ſ�fsD��:y��s��ˑ1X\j|хrdtdB�, ��`.v�q��� �sǑIf�Wfj�52�TKQuto� Set��J� �H5K536(�9i32���91�58(�i9�BA�1(�74O�,A$�(TCP A@k���/�)Y� ��\tpqtool�.v��v���! �conre;a#�C�ontrol R�e�ble��CNRE(�T�<�4�2���pD�)���S�552��q(g�� (򭂯4X��cOux�\sfu;ts�UTS`�i�栜���t�棂���? 6�T�!�SA OO+D6������ ���,!��6c+� igt�t6i��I0�TW8 ���la��vo58�o�bFå����i�Xh��!Xk�|0Y!8\m6e�!G6EC���v��6��@�������<16�A���A�6s����U�`g�T|ώ���r1�qR��˔Z4�T��� ��,#�eZp)g����<ONO0���uJ��t�CR;��F�a� xS�P�f��prdsuGchk �1��2&&$?���t��*D%$�r (�✑�娟:r��'��s�qO��<scr�c�C�\At�trld J"o�\�V�����Paylo�nf�irm�l�!�87���7��A�3ad �! �?ވI�?plQ��3��3"�q��x pl�`���d7��l�calC�uDu�8��;��mov������initX�:s8�O��a�r4 ��r6�7A4|�e Generatiڲ���q7g2q$��g R�� (Sh��c ,D|�bE��$Ԓ\P�:�"��4��4�4,�. sg��5�F�$d6"e;Qp "�SHAP�TQ n7gcr pGC�a(��&"� ��"GDAL¶��r6�"aW<�/�$dataX:s�"tpad��[q�%tput;a__O7;a��o8�1�yl+s�r �?�:�#�?�5x�?�:	c O�:y O�:�IO�s`O%g�qǒ�?��@0\��"o�j92�;!�Ppl.Col�lis�QSkip #��@5��@J��D��@@\ވ�C@X�7���7�|s2��ptcls�LS�DU�yk?�\_ ets�`�< \�Q��@��d�`dcKqQ�FC;�b�J,�n��` (�D�4eN����T�{ ���'j(�c�����/�IӸaȁ��̠H������зa�e\�mcclmt "�CLM�/��� ma�te\��lmpA�LM�?>p7qmc?����2vm�q��%�3s��_sv90�_x�_msu�2L^v_0� K�o�{in�8(|3r<�c_log8r��rtrcW�E �v_3�~yc롘�d�<�te��d�er$cCe� F	iρ�R��Q�?|�l�enter߄�|��(Sd��1�T�X�+fK�r�a99�sQ9+�5�r\t�q\� "FNDR����STD~n$LANG�Pgui��D⠓�S������sp�!ğ֙uf�ҝ�s����$�����e+�=����������������w�H�r\fn_�ϣ��$`x��tcpma��- �TCP�����R638 R�Ҡ��+38��M7p,���� ��$Ӡ�8p0Р�VS,�6>�tk��99�a�� B3���PզԠ��D�2�����UI��t���hq B���8��������p����re�ȿ��exe@4φ�B���e38�ԡG�rmpWXφ�var@�φ�3N�����vx�!ҡ��qҿRBT $c�OPTN as�k E0��1�R �MAS0�H593>/�96 H50�i�+480�5�H0��Dm�Q�K��7�0�g��Pl�h0ԧ�2�OR�DP��@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`m��b��7Г.f��u�d��r>��splayD�E����1w�UPDT |Ub��887 (��Di{���v�Ӛ�� �⧔��#�B��㟳��o  ����a������60q��B���>��qscan��B���ad@�������q`�䗣�#���8��`2�� vlv�䀃Ù�$�>�b���!y S��Easy/���Util��룙�511 J�����9R7 ��Nor֠��inc),<6Q�� �`c��"4�[���G986FVRx S1o����q�nd6��� �P��4�a\ (��
  �������d��K�b9dZ���men7���o- Me`tyF���Fb�0�TUa�'577?i3R��\�5�u?��!� n���f������l\mh�Ц�űE|hmn�	��<!\O���e�1�� l!��y��Ù�\|p����B�����mh�@��:. aG!���/�t�55�`6�!X�l�.us��|Y/k)ensubL�
��eK�h�� �B \1;5g?y?�?�?D��?�*rm�p�?Ktbox O2K|?�G��C?A%ds���?1ӛ#� �TR��/��P� 4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ă�Q23t.�P׀al��Pr+OP517��#IN0a��Q(}g�N�PESTf3ua�P B�l�ig�h�6�aq���P � xS���`  n�0mb�umpP�Q969�g�69�Qq��P0�b�aAp�@Q� BOqX��,>vche�s�>vetu㒣=w/ffse�3����]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q<t�waǂ tp�Q҄T�aror Rec�ov�b�O�P�642����a�q��a�⁠QErǃ�Qry�з`�P'�T�`�aarൄ����	{'�pak7971��71��m0���>�pjot��P�Xc��C�1�adb -v�ail��nag��<�b�QR629�a�Q���b�P  �
�  �P��$�$CL[q �����������$�PS_DIGI�T��� "�!�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv��������*璬�1:PRODUC�T�Q0\PGST�K�bV,n�9�9�\���$�FEAT_IND�EX��~��� 搠ILECOMP ;���)��"��SETUP2 <����  N� !�_AP2B�CK 1=� � �)}6/E+%,/i/��W/�/~ +/�/O/�/s/�/?�/ >?�/b?t??�?'?�? �?]?�?�?O(O�?LO �?pO�?}O�O5O�OYO �O _�O$_�OH_Z_�O ~__�_�_C_�_g_�_ �_	o2o�_Vo�_zo�o o�o?o�o�ouo
�o .@�od�o�� �M�q���<� �`�r����%���̏ [�������!�J�ُ n�������3�ȟW�� ����"���F�X��|� ���/���֯e����� �0���T��x���� ��=�ҿ�s�ϗ�,Ϡ��9�b�� P/� 2) *.VRiϳ�!�*�����0�����PC�7�>!�FR6:"�c��χ��T��߽߀Lը��ܮx���G*.F��>� �	N��,�k��ߏ��STM �����Qа����!�iPend�ant Pane	l���H��F���4�p�����GIF��������u����JPG&P��<�����	PANELO1.DT���� �����2�Y@�G��
3w������//�
4 �a/�O///�/��
TPEINS.�XML�/���\��/�/�!Custo�m Toolba�r?�PASS�WORD/�F�RS:\R?? %�Passwor�d Config �?��?k?�?OH�6O �?ZOlO�?�OO�O�O UO�OyO_�O�OD_�O h_�Oa_�_-_�_Q_�_ �_�_o�_@oRo�_vo o�o)o;o�o_o�o�o �o*�oN�or� �7��m��&� ��\�����y��� E�ڏi������4�Ï X�j��������A�S� �w�����B�џf� ������+���O���� �����>�ͯ߯t�� ��'���ο]�򿁿� (Ϸ�L�ۿpς�Ϧ� 5���Y�k� ߏ�$߳� �Z���~�ߢߴ�C� ��g�����2���V� ���ߌ���?���� u�
���.�@���d��� ����)���M���q��� ��<��5r� %��[�& �J�n��3 �W���"/�F/ X/�|//�/�/A/�/ e/�/�/�/0?�/T?�/ M?�??�?=?�?�?s? O�?,O>O�?bO�?�O O'O�OKO�OoO�O_ �O:_�O^_p_�O�_#_ �_�_Y_�_}_o�_�_�Ho)f�$FILE�_DGBCK 1�=��5`��� ( ��)
SUMMAR�Y.DGRo�\M�D:�o�o
`D�iag Summ�ary�o�Z
CONSLOG�o�o�a�
J�aConsole logK��[�`MEMCH�ECK@'�o��^qMemory �Data��W��)�qHADO�W���P��sS�hadow Ch�angesS�-c-���)	FTP�=��9����w`qm�ment TBD�׏�W0<�)ETHERNET̏��^�q�Z��aEthernet bp�figurati�on[��P��DCSVRFˏ��Ïܟ�q�%�� verify allߟ�-c1PY���DI�FFԟ��̟a��p{%��diffc���q��1X�?�Q��� ����X��CHGD��¯ԯ�i��px��� ���2p`�G�Y�� ��� �GD��ʿܿq���p���Ϥ�FY3ph�O�a��� ��(�GD������y���p�ϡ�0�UP?DATES.�Ц�~�[FRS:\������aUpdates List����kPSRBWLD'.CM.��\��B���_pPS_ROBOWEL���_���� o��,o!�3���W��� {�
�t���@���d��� ��/��Se��� ��N�r�  =�a�r�& �J���/�9/ K/�o/��/"/�/�/ X/�/|/�/#?�/G?�/ k?}??�?0?�?�?f? �?�?O�?OUO�?yO O�O�O>O�ObO�O	_ �O-_�OQ_c_�O�__ �_:_�_�_p_o�_o ;o�__o�_�o�o$o�o Ho�o�o~o�o7�o 0m�o� ��V �z�!��E��i� {�
���.�ÏR����� �����.�S��w�� ����<�џ`������ +���O�ޟH�������8���߯n����$�FILE_��PR����������� �MDONLY 1=4�~� 
 ��� w�į��诨�ѿ���� ���+Ϻ�O�޿sυ� ϩ�8�����n�ߒ� '߶�4�]��ρ�ߥ� ��F���j�����5� ��Y�k��ߏ���B� ����x����1�C��� g������,���P��� ������?��Lu~�VISBCKR�|<�a�*.VD||�4 FR:\���4 Visi�on VD file� :Lbp Z�#��Y�} /$/�H/�l/�/ �/1/�/�/�/�/�/ ? �/1?V?�/z?	?�?�? ??�?c?�?�?�?.O�? ROdOO�OO�O;O�O �OqO_�O*_<_�O`_��O�__%_�_�MR_GRP 1>4��L�UC4  ;B�P	 ]�o�l`�*u����RHB ���2 ��� �?�� ���He�Y �Q`orkbIh�oJd�o�Sc�o�oE��� L�
~K,t��F�5U�aS%�
�o�o 8��e�B���A��b(�Q6����;o}>)���><�rlq�Q>�:0�xq�o� F�@ �r�d�a}J���NJk�H�9�Hu��F!��IP�s}�?�`�.9�<�9�89�6C'6<,6\b�1�,.��g�R���v�A�PA� ����|�ݏx���%� �I�4�F��j����� ǟ���֟��!��E�X`r�UBH�P�c�������ů�R
6�P;�uP<z�˯`��e�Q cB��P<5���@�33@����4�m�,�@UUU�U�~w�>u.�?!x�^��ֿ����3��=[z��=�̽=V6�<�=�=��=$q��~��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�Ϡ Cώ���C�
�P��P'�6��_V�  m�o��To��xo�ߜo ������A�,�e�P� b���������� ���=�(�a�L���p� ���������������� *��N9r]�� ������8 #\nY�}�� �����/ԭ//A/ �e/P/�/p/�/�/�/ �/�/?�/+??;?a? L?�?p?�?�?�?�?�? �?�?'OOKO6OoO�O HߢOl��ߐߢ��O��  _��G_bOk_V_�_z_ �_�_�_�_�_o�_1o oUo@oyodovo�o�o �o�o�o�oN u����� ����;�&�_�J� ��n�������ݏȏ� �%�7�I�[�"/�� ������ٟ������� 3��W�B�{�f����� ��կ�������A� ,�e�P�b��������O �O�O��O�OL�_ p�:_�����Ϧ����� ���'��7�]�H߁� lߥߐ��ߴ������� #��G�2�k�2��V w�����������1� �U�@�R���v����� ��������-Q �u���r��6 ��)M4q \n������ /�#/I/4/m/X/�/ |/�/�/�/�/�/?ֿ �B?�f?0�BϜ?f� �?���/�?�?�?/OO SO>OwObO�O�O�O�O �O�O�O__=_(_a_ L_^_�_�_�_���_�� o�_o9o$o]oHo�o lo�o�o�o�o�o�o�o #G2kV{� h������� C�.�g�y�`������� ���Џ���?�*� c�N���r�������� ̟��)��M�_�&? H?���?���?�?�?�� ��?@�I�4�m�X�j� ����ǿ���ֿ��� �E�0�i�Tύ�xϱ� ����������_,��_ S���w�b߇߭ߘ��� ��������=�(�:� s�^��������� ��'�9� �]�o��� ��~����������� ��5 YDV�z ������1 U@yd��v� ����/Я*/��
/ �u/��/�/�/�/�/ �/�/??;?&?_?J? �?n?�?�?�?�?�?O �?%OOIO4O"�|OBO �O>O�O�O�O�O�O!_ _E_0_i_T_�_x_�_ �_�_�_�_o�_/o�� ?oeowo�oP��oo�o �o�o�o+=$a L�p����� ��'��K�6�o�Z� �����ɏ��폴�  ��D�/ /z�D/�� h/ş���ԟ���1� �U�@�R���v����� ӯ������-��Q� <�u�`���`O�O�O�� �޿��;�&�_�J� oϕπϹϤ������ ��%��"�[�F��Fo �ߵ����ߠo��d�!� ��W�>�{�b��� ������������A� ,�>�w�b����������������=���$FNO ����\_�
F0l q � FLAG>�(�RRM_CHKT_YP  ] ���d �] ��O=M� _MIN� 	����� �  �XT SSB_CF�G ?\ �����OTP_DEF_OW  	���,IRCOM�� >�$GENO�VRD_DO���<�lTHR� �d�dq_ENB�] qRAVC_GRP 1@�I X(/ %/ 7//[/B//�/x/�/ �/�/�/�/?�/3?? C?i?P?�?t?�?�?�? �?�?OOOAO(OeOpLO^O�OoROU��F\� ��,�B,�8�?����O�O�O	__���  DE_�Hy_�\@@m_B�=�vR/���I�O�SMT�G��SUoo&oRHoOSTC�1H�I�� ��zMS5M�l[bo�	127.0�`=1�o  e�o�o �o#z�oFXj�|�l60s	ano?nymous��0�����=ao�
&�&��o�x��o ������ҏ�3�� ,�>�a�O�������� ��Ο�U%�7�I��]� ���f�x�������� ү����+�i�{�P� b�t���������� ��S�(�:�L�^ϭ� oϔϦϸ������=� �$�6�H�Zߩ���Ϳ s����������� � 2���V�h�z��߰� ��������
��k�}� �ߡߣ���߬����� ����C�*<Nq� _������-� ?�Q�c�eJ��n� ������/ "/E�X/j/|/�/�/ �%'/?[0? B?T?f?x?��?�?�? �?�??E/W/,O>OPO�bO�KDaENT 1=I�K P!�?�O  �P�O�O�O �O�O#_�OG_
_S_._ |_�_d_�_�_�_�_o �_1o�_ogo*o�oNo �oro�o�o�o	�o- �oQu8n�� ������#�� L�q�4���X���|�ݏ ���ď֏7���[����B�QUICCA0��h�z�۟��1ܟ��ʟ+���2,����{�!ROUTE�R|�X�j�˯!P�CJOG̯��!�192.168�.0.10��}GN�AME !�J!?ROBOT�vN�S_CFG 1H��I ��Auto-sta�rted�$FTP�/���/�?޿#? ��&�8�JϏ?nπ� �Ϥ�ǿ��[������"�4�G�#������� �������������� ��&�8�J�\�n��� �����������/�/ �/F���j��ߎ����� ��������0S� T��x����� !�3��G,{�Pb t��C���� /�:/L/^/p/�/ ���	/�/=? $?6?H?Z?)/~?�?�? �?�/�?k?�?O O2O DO�/�/�/�/�?�O�/ �O�O�O
__�?@_R_ d_v_�_�O-_�_�_�_ �_oUOgOyO�O�_ro �O�o�o�o�o�o�_ &8Jmo�o�� ���o)o;oMoO !��oX�j�|�����o ď֏����/���B��T�f�x���^�ST_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
�FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@�G %j%D�F��GI6���MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�a��3Ŀ�
��؇Mr��?�9�4�"}~q�_DCd~�1PL_NAME !<u�� �!Def�ault Per�sonality� (from FwD) �4RR2k!� 1j)TEX)�TH��!�AX d �?>?P?b?t?�?�?�? �?�?�?�?OO(O:O�LO^OpO�O�O�Ox2 -?�O�O�O__0_B_T_f_x_�b<�O�_�_ �_�_�_�_o o2oDo�Voho&xRj" 1o��)&0\�b, ��9��b�a @D7�  �a?��c�a�?�`�a�aA'�6x�ew;�	l�b�	 �x7Jp��`�`�	p �< ��(p� �.r� K��K ��K�=*�J���J?���JV��kq`q�P�x�|� �@j�@T;f�r�f�q�acrs��I�� ��p����p�r�ph}�3���´  � ��>��ph�`z���꜖"�Jm�q� H�N��ac����dw��  _�  P� Q� }�� |  а��m�Əi}	'� �� �I� ��  ����:��È�È=̣��(�ts�a	����I  �n �@H�i~�ab�Ӌ�b��w��urN0�� � 'Ж�q�p@2?��@����r�q�5�C�pC0C�G@ C����`O
�A1]w@B�UV~X�
nwB0"h�A��p�ӊ�p@����aDz���֏����Я	�pv�( �� -���I��-�=��A�a��we_q�`�p �?�ff ��m��>� ����Ƽ�uq@ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`�� <
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC�������� #/*/c/N/wi�6����v/C�`� CCHs/`
=$�p�<!��!��ܼ�'�3A��A�AR1A�O�^?�$�?���5p±
=�ç>����3�W
=�#�]��;e��?������{����<��>(�B��u��=B0�������	�R��zH�F�G����G��H��U`E���C��+��}I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0w/O*OONO9O rO]O�O�O�O�O�O�O �O_�O8_#_\_G_�_ �_}_�_�_�_�_�_�_ "oooXoCo|ogo�o �o�o�o�o�o�o	 B-fQ�u�� �����,��P� b�M���q�����Ώ�� �ݏ�(��L�7�p� [������ʟ���ٟ ���6�!�Z�E�W���:#1($1��9�K����ĥ%��x��Ư!3�8��<�!4Mgs���,�IB+8�J��a?���{�d�d������ȿ���ڼ%P8�P�=:GϚ�`S�6�h�z���R��������������  %�� ��h�Vߌ�z� ��&�g�/9�$�������7����A�S�e�w�  ��������������2 wF�$�&Gb���������!C����@���8�����F�� DzN��� F�P D�������)#B�'9�K]o#?��ͫ@@v
��8��8��8�.
 v���!3 EWi{�����:� ��ۨ��1��$MSKCFMAP  ��� ����(.�ONREoL  �!�9��EXCFEN�BE'
#7%^!FN�Ce/W$JOGOV�LIME'dO S"d��KEYE'�%��RUN�,�%��SFSPDTY�0g&P%9#SIGN|E/W$T1MOT�/�T!�_CE_G�RP 1p��#\x��?p��?�? �?�?�?O�?OBO�? fOO[O�OSO�O�O�O �O�O_,_�OP__I_ �_=_�_�_�_�_�_o�o�_:o�TCO�M_CFG 1qB	-�vo�o�o
Va__ARC_b"��p)UAP_CPL��ot$NOCHEC�K ?	+ �x�%7I[ m���������!�.+NO_WAIT_L 7%S2�NT^ar	+��s�_ERR_12s	)9�� ,ȍޏ���x���&��dT�_MO��t��, �p*oq�9�PA�RAM��u	+���a�ß'g{�� �=?�345678901��,��K� ]�9�i�������ɯۯ��&g�����C���cUM_RSPA�CE/�|����$?ODRDSP�c#6�p(OFFSET_�CART�o��DI�Sƿ��PEN_FILE尨!�ai��`�OPTION_I�O�/��PWORK� ve7s#  ��V�ؤ!!�p�4�p�	 ���p��<����RG_DSBOL  ��P#���ϸ�RIENTT5OD ?�C�� !�l�UT_SIM�_D$�"���V~��LCT w}��h�iĜa[�1�_PEsXE�j�RATv�Ш&p%� ��2^3j)TEX)TH�)�X d3����� ��%�7�I�[�m�� �������������!�3�E���2��u��� ������������c�<d�ASew� ��������썒^0OUa0o(ҿ�(����>u2, ���O ~H @D�  [?�aG?��cc��D][�Z�;��	ls��xoJ���������< ���� ��ڐH�(��H3k7H�SM5G�22G���Gp
͜��'f�/-,ڐC%R�>�D!�M#{|Z/��3�����4y H "�c/u/��/0B_���{�jc��t�!�/ �/�"t32�����/6  ���P%�Q%��%�|�T��S62�q?'e	'�� � �2I�� �  �=�+==��ͳ?�;�	�h	�0�I  ?�n @�2�.��Ov;��ٟ?&g9N�]O  ''�uDt@!� C�C�@F#�H!�/�O�O sb
����@�@�H�@�e0@B�QA�0Yv: �13Uwz$oV_�/z_e_�_�_�	��( �� -�2�1�1ta��Ua�c���:Ar����.  �?�ff ���[o"o�_U�`oDX�0A8���o�j>�1'  Po�V(���e�F0�f�Y���L�?�����xb0@<�
6b<߈;�܍�<�ê<� <�&�,/aA�;r�@Ov0P�?fff?�0?&�ip�T@�.{r�?J<?�`�u#	 �Bdqt�Yc�a� Mw�Bo��7�"�[� F��j�������ُ� ���3����,����(�E�� E�~�3G+� F��a ��ҟ�����,��PP�;���B�pAZ� >��B��6�<OίD��� P��t�=���a�s���<��6j�h��7o��>�S��O��0���Fϑ�A�a�_���C3Ϙ�/�%?��?���������#	�Ę��P �N||CH���Ŀ�������@I�_�'�3�A�A�AR1�AO�^?�$��?�����±
�=ç>�����3�W
=�#�\ U��e���B��@���{����<����(�B��u��=B�0�������	�b�H�F�G����G��H��U`E���C��+��I#��I��HD��F��E��R�C�j=[�
�I��@H�!�H�( E<YD0߻������ ��� �9�$�]�H�Z� ��~������������� #5 YD}h� ������
 C.gR���� ���	/�-//*/ c/N/�/r/�/�/�/�/ �/?�/)??M?8?q? \?�?�?�?�?�?�?�? O�?7O"O[OmOXO�O |O�O�O�O�O�O�O�Ot3_Q(�������b��gUU���W_i_2�3�8�x�_�_2�4Mgs�_��_�RIB+�_�_�a���{�m iGo5okoYo�o}l��%P'rP�nܡݯ�o�=_�o�_�[R�?Q�u���  �p���o��/� �S��z
uүܠ�������ڱ�������8����  /�M��w�e��������l2 �F�$��Gb���t��a�`�p�S�C�y�@p�5�G�Y�۠�F� Dz��� F�P D�!�]����پ��ʯ�ܯ� ��~�?��W�@@�?�K��K���K���
 �|�������Ŀ ֿ�����0�B�TϸfϽ�V� ���{���1��$PAR�AM_MENU �?3���  DE�FPULSEr��	WAITTMO{UT��RCV��� SHELL�_WRK.$CU�R_STYL���	�OPT��P�TB4�.�C�R_DECSN���e�� ߑߣ���������� �!�3�\�W�i�{�����USE_PRO/G %��%����.��CCR���e�����_HOST �!��!��:���T �`�V��/�X��>��_TIME��^���  ��GDE�BUG\�˴�GI�NP_FLMSKĻ���Tfp����PG�A  ����)CyH����TYPE��������� �� -?hc u������� //@/;/M/_/�/�/ �/�/�/�/�/�/??�%?7?`?��WORD� ?	=	R}Sfu	PNSU�Ԝ2JOK�DR�TEy�]TRACECTL 1x3���� �`��`&�?�3�6DT �Qy3�%@�0Do � �c2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�Z� .O|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� �p����� *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o� $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������������(��$PG�TRACELEN�  )�  �_�(��>��_UP z����m�u�Y��n�>�_CFG �{m�W�(�~����PКӂ�DEFS_PD |��'ѶP��>�IN��T_RL }��(��8����PE_CO�NFI��~m�'�mњ��ղ�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�p�ح֚��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P;t _��������  Dz (�
 H�X~i�� ����/�/D/�//h/S/�/��
V�7.10beta�1��  A��E�"ӻ�Ay (�� ?!G��!/>���"����!����!BQ��!A\� �!���!2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?OO :O%O7OpO[O�OO�O �O�O�O�O_�O6_!_ Z_E_~_i_�_�_�_�_ �_�_'o2o�_VoAo So�owo�o�o�o�o�o �o.R=v1�<�/�#F@ �y�} ��{m��y=��1� '�O�a��?�?�?���� ��ߏʏ��'��K� 6�H���l�����ɟ�� �؟�#��G�2�k� V���z��������o ��ίC�.�g�R�d� ���������п	��� -�?�*�cώ���� �������B�;� f�x�������DϹ��� ���������7�"�[� F�X��|������� ����!�3��W�B�{� f��������� ��� ��/S>wbt ������ =OzόϾψ��� �ϼ� /.�'/R�d� v߈߁/0�/�/�/�/ �/�/�/#??G?2?k? V?h?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O���O�O�O_ _?_*_c_N_�_r_�_ �_�_�_�_o�_)oT fx�to���/ �o/>/P/b/t/ mo�|���� ���3��W�B�{� f�x�����Տ����� ��A�S�>�w�b��� �O��џ������+� �O�:�s�^������� ͯ���ܯ�@oRodo �o`��o�o�o��ƿ�o ���*<N�Y�� }�hϡό��ϰ����� ���
�C�.�g�Rߋ� v߈��߬�����	��� -��Q�c�N�ﲟ�� ��l��������;� &�_�J���n������� ����,�>�P�:L ����������� �(�:�3��0iT �x�����/ �///S/>/w/b/�/ �/�/�/�/�/�/?? =?(?a?s?��?�?X? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O*\&_8_r���_�_��$PL�ID_KNOW_�M  ��� Q�TSV ����P��?o"o4o�O�XoCoUo�o R�SM_GRP 1��Z�'0{`�@�`uf�e�`
�5� �g pk'Pe ]o�����������SMR�c�b�mT�EyQ}? yR ����������폯��� ӏ�G�!��-����� ������韫���ϟ� C���)���������`��寧���QST�a�1 1��)��v�P0� A 4� �E2�D�V�h������� ߿¿Կ���9��.� o�R�d�vψ��ϬϾϔ���2�0� Q�<3��3�/�A�S��4l�~ߐߢ��A5���������6
��.�@��7Y�k�}����8���������MAD  �)��PARNU/M  !�}o+���SCHE� S�
���f���S��UPD�f�x��_C�MP_�`H�� �'��UER_CHK-���ZE*�<RSr��_�Q_M�OG���_�X�__RES_G��!� ��D�>1bU �y�����/ �	/����+/ �k�H/g/l/��Ї/ �/�/�	��/�/�/� X�?$?)?���D?c?�h?����?�?�?�V� 1��U�ax�@c�]�@t@(@c�\�@�@D@c�[�*@��THR_INRr�J�b�U�d2FMASS?O �ZSGMN>OqCMO�N_QUEUE ���U�V P~P *X�N$ UhN�FV��@END�A��IEcXE�O�E��BE�@|�O�COPTIO�G���@PROGRAoM %�J%�@��?���BTASK_�IG�6^OCFG ���Oz��_�PDA�TA�c��[@Ц2=�DoVohozo�j 2o�o�o�o�o�o�);M jINFO
[��m��D�� ������1�C� U�g�y���������ӏ����	�dwpt�l �)�QE DIT ���_i��^WER�FLX	C�RGA�DJ �tZAЄ����?נʕFA��I�ORITY�GW�>��MPDSPNQ�����U�GD��OT�OE@1�X� _(!AF:@E� �c�Ч!tcp|n���!ud��>��!icm���?n<�XY_�Q�X�{��Q)� *�1�5��P��]�@� L���p��������ʿ ��+�=�$�a�Hυ�z��*��PORT)Q�H��P�E��_CARTREPP|X��SKSTA�H^�
SSAV�@�tZ�	2500H8�63���_x�
�'��*X�@�swPtS��ߕߧ���URGE��@B��x	WF��DO�F"[W\��������WRUP_DE?LAY �X��ԟR_HOTqX	B%��c���R_NOR�MALq^R��v�S�EMI�����9�Q�SKIP'��tUr�x 	7�1�1� �X�j�|�?�tU���� ����������$ J\n4���� ����4FX |j����� ��/0/B//R/x/�f/�/�/�/tU�$R�CVTM$��D��� DCR'����Ў!>s>.B<� >C^�>���r8�Y7){��:���YF����̮�&�w�:�o?�� <
6�b<߈;܍��>u.�?!<�&�?h?�? �?�@>��?O O2ODO VOhOzO�O�O�O�O�O �?�O�O__@_+_=_ v_Y_�_�_�?�_�_�_ oo*o<oNo`oro�o �o�o�_�o�o�o�o �o8J-n��_� ������"�4� F�X�j�U������ď ���ӏ���B�T� �x���������ҟ� ����,�>�)�b�M� �����������ïկ �Y�:�L�^�p����� ����ʿܿ� ���� 6�!�Z�E�~ϐ�{ϴ� ������-�� �2�D� V�h�zߌߞ߰����� ����
���.��R�=� v��k�������� ��*�<�N�`�r��� ������������� &J\?���� �����"4�FXj|��!GN_ATC 1�	;� AT&�FV0E0��ATDP/6/9�/2/9�AT�A�,AT�%G1%B960��+++�,��H/,�!IO_TYPE  �%��#t�REFP�OS1 1�V+O x�u/�n �/j�/
=�/�/�/Q? <?u??�?4?�?X?�?��?�+2 1�V+ �/�?�?\O�?�O�?�!3 1�O*O<OvO��O�O_�OS4 1��O�O�O_�_t_�_>+_S5 1�B_T_�f_�_o	oBo�_S6 1��_�_�_5o�o��o�oUoS7 1� lo~o�o�oH3l�oS8 1�%�_���SMA�SK 1�V/  q
?�M��XNOS/��r������!MO�TE  n��$��_?CFG ����q����"PL_RAN�G�����POWE/R ������SM_DRYPR/G %o�%�P���TART ���^�UME_PR�O-�?����$_EX�EC_ENB  y���GSPD��pՐݘ��TDB���
�RM�
�MT_�'�T����OB�OT_NAME �o����OB�_ORD_NUM� ?�b!�H863  ��կ���P�C_TIMEOU�T�� x�S23�2Ă1�� L�TEACH ?PENDAN��wƋ�-��M�aintenance Cons�䃌s�"���KC�L/Cm��

����t�ҿ No Use-��Ϝ�0��NPO�򁋁���.�CH_Lf������q	��~s�MAVAIL������糅��SPA�CE1 2��, j�߂�D��s��߂� �{S�8�?�k�v�k�Z߬� �ߤ��ߚ� �2�D� ��hߊ�|��`����� ������ �2�D� ��h��|���`�����P����y���2��� �0�B���f�����@{���3 );M_�������/� /4 4FXj|*/�� �/�/�/?(??=?5Q/c/u/�/�/G?�/ �/�?O�?$OEO,OZO6n?�?�?�?�?dO �?�?_,_�OA_b_I_w_7�O�O�O�O�O �_�O_(oIoo^oofo�o8�_�_�_�_ �_�oo6oEf){���G �No� ���
M� ���*�<�N� `�r�������w���o �収���d.�� %�S�e�w��������� ��Ǐَ���Θ8�+� =�k�}�������ůׯ ͟����%�'�X�K� ]���������ӿ�������#�E�W� `� @����� ��x�����\�e��� ��������R�d߂� 8�j߬߾߈ߒߤ��� �������0�r��� X������������8����
�ύ�_MODE  �{^��S ��{|�2�0�����3��	S|)CWOR�K_AD��WX��+R  �{��`� �� _INT�VAL���d���R_OPTION�� ��H VAT_GRP 2��uwp(N�k|��_ �����/0/B/ ��h�u/T� }/�/�/ �/�/�/�/?!?�/E? W?i?{?�?�?5?�?�? �?�?�?O/OAOOeO wO�O�O�O�OUO�O�O __�O=_O_a_s_5_ �_�_�_�_�_�_�_o 'o9o�_Iooo�o�oUo �o�o�o�o�o�o5 GYk-���u �����1�C�� g�y���M�����ӏ� ��	��-�?�Q�c��� �������������ǟ�;�M�_����$�SCAN_TIM��_%}�R ��(�#((�<}04d %d 
!D�ʣ��u�/�����+U��25���@�d5�P�g��]	���������dd��x�  P���w� ��  8� �ҿ�!���D�� $�M�_�qσϕϧϹπ�������ƿv��F�X��/� �;�ob��p�m��t�_D�iQ̡  � l�|�̡ĥ������ �!�3�E�W�i�{�� ������������� /�A�S�e�]�Ӈ��� ����������) ;M_q���� ���r���j� Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�%�/  0��6��!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O*�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo�O�OJ�o �o�o�o�o�o�o  2DVhz��������
�7?  ;�>�P�b�t����� ����Ǐُ����!� 3�E�W�i�{�������ß �ş3�ܟ� �&�8�J�\�n������������ɯ���;�,� �+��	123456{78�� 	� =5���f�x�������������
�� .�@�R�d�vψϚ�� ����������*�<� N�`�r߄߳Ϩߺ��� ������&�8�J�\� n�ߒ��������� ���"�4�F�u�j�|� �������������� 0_�Tfx�� �����I >Pbt���� ���!/(/:/L/ ^/p/�/�/�/�/�/�/�2�/?�#/9?�K?]?�iCz  �Bp˚   ��h2��*�$SC�R_GRP 1��(�U8(�\x�d�@� � ��'�	 �3�1�2�4(1*� &�I3�F1OOXO}m7��D�@�0�ʛ)���HUK�L�M-10iA 890?�90;��F;�?M61C D�:��CP��1
\&V �1	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^� oOUO>oPo#G�/血��o'o�o�o�o�oB�0�rtA9A�0*  @�BuD&Xw?��ju�bH0�{UzAF@ F�`�r��o��� ��+��O�:�s��m�Bqrr����������B�͏b����7�"�[� F�X���|�����ٟğ ���N���AO�0�B��CU
L���E�jqBq=g��Ҕ�$G@�@pnϯ B���G��I
E�0EL_DE�FAULT  ~�T��E���MIPOWE?RFL  
E*���7�WFDO�� *��1ERVENT 1���`�(�� L!DU�M_EIP��>���j!AF_IN�E�¿C�!FT$������!o:�� ��a�!RPC_MAINb��DȺPϭ�t�VIS�}�Cɻ����!TMP��PU�ϫ�d���E�!
PMON_�PROXYF߮�e 4ߑ��_ߧ�f�����!RDM_SR�V�߫�g��)�!�R�Iﰴh�u�!%
v�M�ߨ�id����!RLSYNC���>�8���!gROS��4��4�� Y�(�}���J�\����� ��������7��[ "4F�j|�� ��!�Eio��ICE_KL ?�%� (%S?VCPRG1n>���3��3���4//�5./3/�6V/[/�7~/�/�H�D�/�9�/�+� @��/��#?��K? ��s?� /�?�H/ �?�p/�?��/O� �/;O��/cO�?�O �9?�O�a?�O��? _��?+_��?S_� O{_�)O�_�QO�_ �yO�_��Os�� ��>o�o}1�o�o�o �o�o�o�o;M 8q\����� ����7�"�[�F� �j�������ُď�� �!��E�0�W�{�f� ����ß���ҟ�� �A�,�e�P���t���������ί�y_D�EV ���MC:�@`]!�OUT���2��REC 1��`e�j� �	 �����˿���8ڿ��
 �`e�� �6�N�<�r�`ϖτ� ���Ϯ�������&�� J�8�n߀�bߤߒ��� ��������"��2�X� F�|�j�������� ������.�T�B�x� Z�l������������� ,P>`bt ������( L:\�d�� ��� /�$/6// Z/H/~/l/�/�/�/�/ .��/?�/2? ?V?D? f?�?n?�?�?�?�?�? 
O�?.O@O"OdORO�O vO�O�O�O�O�O�O_ _<_*_`_N_�_�_x_ �_�_�_�_�_oo8o o,ono\o�o�o�o�o �o�o�o�o "4 jX������ ����B�$�f�T� v������������؏ ��>�,�b�P�r����p�V 1�}� P�
�ܟ� G��T�YPE\��HEL�L_CFG ��.��͟  x	�����RSR�� ����ӯ������� ?�*�<�u�`������������  �%�3�E��Q�\���M�o�p�S�d��2��d]�|K�:�HK 1�H� u������� A�<�N�`߉߄ߖߨ� ����������&�8���=�OMM ��H���9�FTOV_�ENB&�1�OW_REG_UI��~�IMWAIT��a���OUT�������TIM������VAL����_�UNIT��K�1�M�ON_ALIAS� ?ew� ( he�#���������� ����);M��q ����d�� %�I[m� <������!/ 3/E/W//{/�/�/�/ �/n/�/�/??/?�/ S?e?w?�?�?F?�?�? �?�?�?O+O=OOOaO O�O�O�O�O�OxO�O __'_9_�O]_o_�_ �_>_�_�_�_�_�_�_ #o5oGoYokoo�o�o �o�o�o�o�o1 C�ogy��H� ���	��-�?�Q� c�u� �������Ϗ� ����)�;��L�q� ������R�˟ݟ�� ���7�I�[�m��*� ����ǯٯ믖��!� 3�E��i�{������� \�տ�����ȿA� S�e�wω�4ϭϿ��� �ώ����+�=�O��� s߅ߗߩ߻�f����� ��'���K�]�o�� ��>���������� #�5�G�Y��}����������n��$SMO�N_DEFPRO ������ *�SYSTEM* � d=��REC�ALL ?}�� ( �}��>Pbt�� ,�� ���;M_ q��(���� //�7/I/[/m// �/$/�/�/�/�/�/? �/3?E?W?i?{?�? ? �?�?�?�?�?O�?/O AOSOeOwO�OO�O�O �O�O�O__�O=_O_ a_s_�_�_*_�_�_�_ �_oo�_9oKo]ooo �o�o&o�o�o�o�o�o��f&copy �mc:diocf�gsv.io m�d:=>insp�iron:507A2ew��n0.r�frs:orde�rfil.dat� virt:\temp\E���t��a(�v*.d���x�h�z����kx�yzrate 61�}H�Z������h�3��xmpbac�k�b�t����� }-*.sdb6�*C�U� Y������3�=�ڐ2636 ߟp��� ��'�9�S�W�����
�k
�� ��˯ݯn� ��������Z�H�Z�� ���"�4���U�a�s� �ϗϪ�E�T�Y�����lߡi.x.�:\�π8�O���n߀ߒߥe/.�a6�H�ܰ^���� �&�8�����m��� �϶���Z������"� 4���X�i�{����߲� C��������0�B� T�ew����I�� ��,���P�a s����;��`� //(����n/�/��/����4940  H/Z/�/�/?"4� �'a?s?�?�?�E?�(�Y?�?�?O!8�$S�NPX_ASG �1����9A�� P 0� '%R[?1]@1.1O 9?�#3%dO�OsO�O �O�O�O�O�O __D_ '_9_z_]_�_�_�_�_ �_�_
o�_o@o#odo GoYo�o}o�o�o�o�o �o�o*4`C� gy������ �	�J�-�T���c��� ����ڏ�����4� �)�j�M�t�����ğ ������ݟ�0��T� 7�I���m�������� ǯٯ���$�P�3�t� W�i��������ÿ� ���:��D�p�Sϔ� wω��ϭ��� ���$� ��Z�=�dߐ�sߴ� �ߩ������� ��D� '�9�z�]������ ����
����@�#�d� G�Y���}��������� ����*4`C� gy����� �	J-T�c� �����/�4/ /)/j/M/t/�/�/�/ �/�/�/�/?0?4,D�PARAM ��9ECA �	U��:P�4�0$H�OFT_KB_CFG  p3?E�4�PIN_SIM  9K�6�?�?�?��0,@RVQSTP/_DSB�>�21O|n8J0SR ��;� & =O{Op0��6TOP_ON_ERR  p4��9�APTN ��5�@A��BRING_PR�M�O J0VDT_GRP 1�Y9�@  	�7n8_ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2Dk hz������ �
�1�.�@�R�d�v� ��������Џ���� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\����������� ȯگ����"�I�F� X�j�|�������Ŀֿ ����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�tߛ� �ߪ߼��������� (�:�a�^�p���� �������� �'�$�6� H�Z�l�~���������������3VPRG_�COUNT�6�8�A�5ENB�O�M=�4J_UPD� 1��;8  
p2����� � )$6Hql ~�����/� / /I/D/V/h/�/�/ �/�/�/�/�/�/!?? .?@?i?d?v?�?�?�? �?�?�?�?OOAO<O NO`O�O�O�O�O�O�O �O�O__&_8_a_\_�n_�_�_�_YSDOEBUG" � �P�dk	�PSP_PA�SS"B?�[L�OG ���m�P�X�_  ��g�Q
MC:�\d�_b_MPC m��o�o�Qa�o� �vfSAV žm:dUb�U�\gSV�\TEM_TIME 1�� (�P�TNu]�qT1SVGUNYS} #'k�sp�ASK_OPTICON" �gosp�BCCFG ���| �b��z`����4��X�C� |�g�����ď֏���� ��	�B�-�f�Q�c� ���������ϟ�� ,�>�)�b��YR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz��rBr�|�|� ���z� �%��I� 4�m�X���|������� �֏���3��W�B� g���x�����՟���� ����S�>�w�b� ����'2A ��ʯܯ�� ����E�0�i�T��� x���ÿտ翢���� /��?�e�1�/���/ �ϜϮ��������,� �P�>�`߆�tߪߘ� �߼��������L� :�p�^������� ����� �6�H�>/`� r�������������� �� 0Vhz8 ������
 .�R@vd�� �����//</ */L/r/`/�/�/�/�/ �/�/�/�/?8?&?\? J?�?n?�?�?�?�?�� �?OO�?FO4OVOXO jO�O�O�O�O�O�O_ _�OB_0_f_T_v_�_ �_�_z_�_�_�_oo >o,oboPoroto�o�o �o�o�o�o(8 ^L�p���� ���$��H�6�l� ~�(O����f�d��؏ ���2� �B�D�V��� ����n����ԟ
��� .�@�R�d����v��� �����Я���*�� N�<�^�`�r�����̿ ���޿��$�J�8� n�\ϒπ϶Ϥ����� ��ߊ�(�:�L���|� jߌ߲ߠ��������� �0�B�T��x�f�� ������������,� �P�>�t�b������� ��������:( JL^����� � �6$ZH ~l��^���d� � //D/2/h/V/x/ �/�/�/�/�/�/�/? 
?@?.?d?v?�?�?T? �?�?�?�?�?OO<O *O`ONO�OrO�O�O�O �O�O_�O&__6_8_ J_�_n_�_�_�_�_�_ �_�_"ooFo��po �o,oZo�o�o�o�o �o0Tfx�H �������,� >��b�P���t����� ����Ώ��(��L� :�p�^�������ʟ�� �ܟ� �"�$�6�l� Z���~�����دꯔo ��&�ЯV�D�z�h� ������Կ¿��
�� .��R�@�v�dϚτ��  ���� ��������$TBJ�OP_GRP 2�ǌ�� � ?������������_xJBЌ���9� �< ��X���� @����	 �C��} t�b  C��<��>��͘Ր���>̚йѳ33�=�CLj�f�ff?��?�ff�BG��ь�����t��ކ�>�(�\�)�ߖ�E噙�;���hCYj�� � @h��B�  �A����f��C�  Dhъ�1���O�4�N����
:���Bl^���j�i�l�l����A�ə�A�"��D9��֊=qH����нp�h�Q�;�A�j��o��@L��D	2��������$�6�>B��\��T���Q�ts>x�@33@���C���y�1�����>��Dh�����x�����<{�h�@i� ��t ��	���K& �j�n|��� p�/�/:/k/������!��	V�3.00J�m61cI�*� IԿ���/�' Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I�!CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;��;Q�T,8�4`� *�ϴ?�2����3\�X/O��ESTPARS  ���	���HR@ABL/E 1����0�É
H�7 8��9
GB
H
H����
G	
HE

H
HYE��
H�
H
H6FRD	IAO�XOjO|O�O�O�ETO"_4[>_P_�b_t_�^:BS _�  �JGoYoko}o�o�o�o �o�o�o�o1C Ugy����`#o RL�y�_�_�_�_�O�O��O�O�OX:B�rNUoM  ���P��� V@P:B_CFG ˭��Z�h�@��IMEBF_TT%AU��2@��VERS�q���R 1���
 �(�/����b�  ����J�\���j�|��� ǟ��ȟ֟����� 0�B�T���x�������R2�_���@�
��MI_CHAN��� � ��DBGL�V���������E�THERAD ?U��O������h�����ROUT6�!��!����~��SNMASKD�|�U�255.���#�����OOLO_FS_DI%@�u�.�ORQCTRL �����}ϛ3r� �Ϲ���������%� 7�I�[�:���h�z߯��APE_DETA�I"�G�PON_S�VOFF=���P_?MON �֍��2��STRTCH/K �^������VTCOMPAT���O�����FPRO�G %^�%  BCKEDT-Q�<��9�PLAY&H��_INST_Mްe ������US��q��LCK���Q?UICKME�=�ރ�SCREZ�>G�tps� �� �u�z����_��@@�n�.�SR_GRP� 1�^� �O����
��+ O=sa�쀚 �
m������L/ C1gU�y �����	/�-/�/Q/?/a/�/	1?234567�0�/��/@Xt�1���
� �}ipnl�/� gen.htm�? ?2?D?V?`�Panel _setupZ<}P���?�?�?�?�?�?  �??,O>OPObOtO�O �?�O!O�O�O�O__ (_�O�O^_p_�_�_�_ �_/_]_S_ oo$o6o HoZo�_~o�_�o�o�o �o�o�oso�o2DV hz�1'�� �
��.��R��v����������ЏG���U�ALRM��G ?9� �1�#�5� f�Y���}�������џ�ן���,��P��S�EV  �����ECFG ���롽�A�� :��Ƚ�
 Q��� ^����	��-�?�Q��c�u�����������Ԇ� �����I2��?���(%D�6�  �$�]�Hρ�lϥϐ� �ϴ�������#��Gߌ��� �߿U�I�_Y�HIST 1}��  (��� ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1����(�:�� ����962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V