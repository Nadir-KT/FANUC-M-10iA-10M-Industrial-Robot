��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �ET�H_FLTR.�� $�  � �FTP_C�TRL. @ ?$LOG_8	��CMO>$DN�LD_FILTE�� � SUBDIR�CAP�� HOv��NT. 4� �H_NAME �!ADDRT�YPA H_LE�NGTH' ��z +LS �D $ROBO�TIG PEER�^� MASKM�RU~OMGDEyV#���RDM*��DISABLz&�TCPIG�/ 3 $ARP�SIZ&_IP=F'W_MC��oF_IN� FA~�LASSs�HO�_� INFO��wTELK PV�b	 WOR�D  $AC�CESS_LVL�?TIMEOUT�uORT � �I�CEUS= ��$�#  �����!�� � � VIRTUAL�/�!'0 ��%
���F������$�%�v��+ ��F���$�� �-2%;��SHARED �1�)  P!!�!�?���!|?�? �?�?�?O�?%O�?1O OZOOBO�OfO�O�O �O�O_�O�OE__i_ ,_�_P_�_t_�_�_�_ o�_/o�_SooLo�o xo�opo�o�o�o�o �o*Os6�Z �~�����9� �]� ���D�V���z� ۏ����#���Y��H�}�@���)7z _L�IST 1=x/!1.ܒ0��d��ە1�d�2551.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I����o�������O�6���8�`����� �$� ��-� ���-��%P�%��&!Ò�)�0�H!� ���rj3_tpd����! � �!!K�C� e�0ٙ��&W�!Cm ��w߉�S�?!CON� ��z1�=�smon��W�