��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8GW�+0�$Y $DB\� 6COMW!2�MO� H.	 �\rVE�1$F8�RA{$O�UD�cB]CTMP1_FtE2}G1_�3�B�2�FXD�#
 �d $CARD�_EXIST4�$FSSB_TY�P!AHKBD_YSNB�1AGN Gn� $SLOT�_NUM�APR{EV4DEBU� �g1G ;1_EDIT�1 � 1G�=� S�0%$�EP�$OP��U0LETE�_OK�BUS�P7_CR�A$;4AV�� 0LACIw�1�R�@k �1$@ME=N�@$D�V�Q�`PvVA{'��BL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6�_�7_�8_�94:\qO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"YtP_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0��1p�3� >��DC �� Ќ@��hPV���mEX�p� �0g0xۤ�p�r
$TF��2C$MD3i�TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F�"F��40CP@�a2 6�@$�PPU�3N�)ύRևA�X�!DU��AI�3BUF�F=�@1� |pp���pPIZT� PP�M��M�y��F�SIMQSI�"ܢVAڤtT���Px T�`�(zM��P�B�qFAkCTb�@EW�`P1�BTv?�MC�� �$*1JB8`p�*1DEC��F����=�� ��H0CHNS_EMP1�$G��8��@!_4�3�p|@P��3�TCc�(r/�0-sx� �ܐ� MBi��!�����JR� i�SEGF�R��Iv �aR�TrpN�C��PVF4|>�bx &� �f{uJc!�Ja��� !2�8�ץ�AJ���SIZ�3S�c�B�TM���g�|��JaRSINFȑ b���q�۽�н�����L�3�B���CRC�e�3CCp��� �c��mcҞb�1J�c�P��.����D$ICb�Cq�5r�ե��@v�'����EV���zF��_J��F,pN��ܫ��?�4�0A�! � r���h�Ϩ��p�2��͕a�� �د��R>�Dx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�IM�]pUR��QUA1w  $@TITO1�/S@S�!����"0�?DBPXWO��B0=!5�$SK���2M@DBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z���LB�)$�/���� %�/��$C�!&?�$ENE�q.'*?�Ú �RE�p2(H ���O�0#$L|3$$�#�B[�;�К�FO_D��ROSr�#������3�RIGGER�6P�ApS����ETUR�N�2�cMR_8�T�Uw��0EWM��M�GN�P���B#LAH�<E���P��O&$P� �'P@DT�3�CkD{��DQฑ�4�11��FGO_oAWAY�BMO����Q#!�DCS�_�)  �PIS� I gb {s�C��A��[ �B$�S���AbP�@�EW-�TNTVճ�BV�Q[C� (c`�UWr�P�J��P�<$0��SAFE���V�_SV�bEXCL�U��nONL�<зSY�*a&�OT<�a'�HI_V�4�x�B���_ *P0� 9�_z��p 콁�ASG�� + nrr�@6Acc*b��G��#@E�V.iHb?fAN�NUN$0.$fdID�U�2�SC@�`�i��a��j�f��z��@I:$2,O�$FibW$�}�OT9@�1 ?$DUMMYT��d�a��dn�� � �E-o ` ͑HE4�(sg�*b�SAB��SU�FFIW��@CUA=�c5�g6�a�bMSW�E. 8�Q�KEYI5���T�M�10s�qA�vIN䊱��D��/ Dބ�HOST_P! �rT��ta��tn��tsp��pEMӰV��� S�BLc ULI�0  8	=ȳ�ј �Tk0�!1 � �$S��ESAMPL���j�۰f璱f���I��0��[ $SUB �k�#0�C��T�r#a�SAVʅ��c����C��P�fP$n0E��w YN_B#2� 0Q�DI{dlpO�(��9#$�R_�I�� �ENC�2_S� 3  5�C߰�f�- �SpU����!4�"g�޲r�1T���5X� j`ȷg��0�0K�4�<AaŔAVER�qĕ�9g�DSP�v��PC��r"��(���ƓoVALUߗHE��ԕM+�IPճ��OkPP ��TH���֤��P�S� �۰F��df�J� �q�a�C1+6 H�bLL_DUs�~a3@{�0�3:���OTX"����s�"�0NOAUkTO�!7�p$)�H$�*��c4�(�Cy�%8�C, �"p�&��L�� 8H *8�LH <6����c "�`, `Ĭ�kª�q���q��sq��~q��7*��8��9��0����U1��1̺1ٺ1�U1�1 �1�1ʥ2(�2����2̺2�ٺ2�2�2 �2��2�3(�3��3T��̺3ٺ3�3�U3 �3�3�4("'���?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?g �@P?9��5�9�E�@A���A� ;p$T�P�$VARI�:�Z���UP2�P< ���TDe����K`Q���!��BAC�"= T�p��e$�)_,�bn�kp+ IF�IG�kp�H  ��Pİ�rF@`�!>Gt ;E��sC�ST�D� D���c�<� 	C��{�� _���l���R  ���FORCEUP?b^��FLUS�`H��N>�F ���RD_CM�@E������ ��@vMP��REMr F �Q��1k@���7Q
�K4	NJ�5EFF�ۓ:�@IN2Q��O�VO�OVA�	TgROV���DTՀ�DTMX� � �@�
ے_PH"p��CL��_TpE�@d�pK	_(�Y_T��Tv(��@A;QD� ������!0tܑ&0RQ���_�a��2��M�7�CL�dρ�RIV'�{��EAmRۑIOHPC�@d����B�B��CM9@����R �GCLF�e!DYk(M�a6p#5TuDG��8� �%��FSSD �s�? P�a�!�1����P_�!�(�!1��E��3�!3�+5�&�GSRA��7�@��;ᚔPW��ONn��EBUG_SD2H�P�{�_E A ��p�R �TERM�`5Bi6 �OR�I#e0Ci6 �GSM_�P��e0D�9�TA�9Ei5$Z ��UP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1젎4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ3Q�E�p %B`�'EC����AR$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"�r�A��?���ERV��XQ�Y�� mG>@�BN��U\���R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`�0SMT6�G�3�GR��13�aPA�L@���`�q�uH �� ���TOC�A�`P	P�`$O�P����p�ѡ�`�0O��RE�`R�4C�AO�p낎Be��`R�Eu�h�A��eo$PWR�IMu��RR_�cN��q=B �I&2H���p_A�DDR��H_LE�NG�B�q�q�q$�Rj��S�JڢSS��SKN��u\��u̳�uFٳSE�A�jrS��[MN�!K���0��b����OLX���p����`ACRO 3pJ�@��X�+��Q���6�OUP3�b_"�IX��a�a1��}� ������(��H��D���ٰ��氋�IO
2S�D�����	�7�L $d��`Y!�_OFFr�PR�M_��"�HTT�P_+�H:�M (�|pOBJ]"�p��-$��LE~Cd����N � ��֑AKB_�TqᶔS�`lH�LVh�KR"~uHITCOU��[BG�LO�q����h�����`��`S9S� ���HW�#A�:�Oڠ<`INC�PU2VISIO W�͑��n��to��to�~ٲ �IOLN��P 8��R��p�$SLob PU�T_n�$p��P�& ¢��Y F_AS:�"Q��$L�������Q  U�0	P4A0��^���ZPHY��-���x��UOI �#R `�K����$�u�"pPpk����$�����q1UJ5�S�-���NE6WJOG�KG̲DIS�� c�Kp���#T (��uAVF�+`�CTR<�C
�FLAG2�;LG�dU �������13LG_SIZ�����b�4�a��a�FDl�I`�w� m�_� {0a�^��cg���4��ƀ��Ǝ���{0��� S�CH_���aR�L�N�d�VW���E �"����4��UM�A�r�`LJ�@�DAUfՃEAU�p��d|�r�GqH�b����BOO��WL ?�6 I�T��y0�REC���SCR ܓ�Dx
�\���MARGm� !��զ ��d%�����	S����W���U� ��JGM[�MNCH|J���FNKEY\��K��PRG��UF���7P��FWD��H]L��STP��V��=@��А�RS��HO`����C9T��b ��7�[�UL���6�(R�D� ����Gt��@P�O��������MD�F�OCU��RGEX.��TUI��I��4�@�L�����P����`��P��NE��CANA��Bj�oVAILI�CL !~�UDCS_HII4���s�O�(!�SH���S����__BUFF�!X�5?PTH$m����v`��D���AtrY��?P��j�3��`O+S1Z2Z3Z8|�� Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�AC���K�&&z�� [ LQ��+0 0�	P���`#qdt
�U��dw<���_ \ ?�4Г�\��Ѩ#\0�C4�] ��CL�DPL��UTRQL�I��dڰ�)�$FLAG&�� 1�#�D����'B�LD�%�$�%ORGڰ5�2�PVŇV�Y8�s�T�r�$}d^ A���$6��$�%S�`�T� �B0�4�6RCLMC�4]?o?�9�세�MI�p}d_ Yd=њRQ���DSTB�p� �;F�HHAX�R |JHdLEXCESr�7�CM!p�a`� /B�T�B��`5a�p=F_A7Ji���KbOtH� K�db q\Q���v$MBC��LI|�)SREQU�IR�R�a.\o�AXD�EBUZ�ALt M��c�b�{P����2�ANDRѧ`�`d0;�2�ȺSDC��N�INl�K�x`��X� �N&��aZ���UP�ST� ezrL�OC�RIrp�E�X<fA�p�9AAOwDAQ��f XY�3OND�rMF,� �f�s"��}%�e/� �v�FX3@IGG�� g ��t"���ܓs#N�s$R�a% ��iL��hL�v�@�ODATA#?pE��%�tR��Y�Nh �t $MD`qI�}�)nv� ytq�ytH�P`�Pxu��(�zsAN�SW)�yt@��yuD�+�)\b���0o�i -�@CUw�V�p 0�XeRR2��j D�u�{Q��7Bd$CA�LIA@��G��2N��RIN��"�<E�'NTE��Ck�r^��آXb]���_N�ql@k���9�D���Bm��7DIVFDH�@��:�qnI$V,��Sv�$��$Z��X�o�*����o�H �$BEL�T�u!ACCEL��.�~�=�IRC��� ���D�T�8��$PS�@�"L�� �r��#^�S�Eы T�PATH3���I���3x�p�A_W��ڐ����2nC��4�_M=G�$DD��T���$FW�Rp9���I�4��DE7�P�PABN��ROTSPEE�[g�� �J��[�C@4����$USE_+�VP�i��SYY���1 �qYN!@A�ǦOsFF�qǡMOU��3NG���OL����INC�tMa6��HBx��0HBENCS+��8q9Bp�4�FDm�IN��Ix�]��B��V�E��#�y�23_UyP񕋳LOWL�A��p� B���Du�@9B#P`�x ���BCv��r�MOSI��BM�OU��@�7PERC7H  ȳOV��â 
ǝ����D�Sc@F�@MP����� Vݡ�@y�j�LUk��GjĆp�UP=ó���ĶT�RK��AYLOA�Qe��A��Ԓ����8N`�F�RTI�A$��MOUІ�HB�BS0�p7D5���ë�Z��DUM2ԓS_�BCKLSH_C Ԓk����ϣ����=���ޡ �	ACLA�L"q��1м@��C�HK� �S�RT�Y��^�%E1Qq_��޴_UM�@�C�#��SCL0�r�LMT_J1_L��"9@H�qU�EO�p��b�_�e�k�e�SPC`��u���N�PC�BN�Hz \P��C�0�~"XT��CN_b:�N9��I�SF!�?�V���U�/���ԒdT���CB!�SH� :��E�E1T�T����0y���T��PA ��_P��_� =��Ơ���!����J6 L��@��OG�G�ToORQU��ONֹ���E�R��H�E�g_	W2���_郅T���I�I�I��	Ff`xJ�1�~1��VC3�0BD:B�1��@SBJRK�F9�0DBL_�SM��2M�P_D9L2GRV��0��fH_��d���COS���LNH���������!*,�aZ���fMY�_(��TH��)THET=0��NK23���"l��CB�&CB�CAA�B�"��!��!Ư&SB� 2�%GT	S�Ar�CIMa������,4#97#$DU���H\1� �:Bk6�2�:AQ(rSf$NE�D�`I��B+5��	$̀�!A�%�5�7���LPH�E�2���2SC%C%�2�-&FC0JM&̀V�8V��8߀LVJV!KV�/KV=KVKKVYKVgIH�8FRM��#X�!KH/KH=KHKKH�YKHgIO�<O�8OT�YNOJO!KO/KUO=KOKKOYKOM&�F�2�!+i%0d�7S�PBALANCE�_o![cLE0H_�%SPc� &�b&�b>&PFULC�h�b��g�b%p�1k%�U�TO_��T1T2�i/�2N��"�{� t#�Ѱ`�0�*�.��T��OÀ<�v IN�SEG"�ͱREV84vͰl�DIF�ŕ��1lzw��1m�0OaBpq�я?�MI{����nLCHWAR�Y�_�AB��!�$MECH�!o ��q�AX��P����7Ђ�`n 
�d(�nU�ROB��CRԒ�H���'�MS�K_f`�p P �`_��R/�k�z�����1S�~�|�z�{�ؔ�z��qINUq�MTCOM_C� >�q  ���p~O�$NOREn�����pЂr 8fp GRe�uSD�0�AB�$XYZ�_DA�1a���DE�BUUq������s �z`$��COD��� L���p��$BUFINDX�|�  <�MOR^m�t $فUA� �֐���Ԑ<��r�G��u � $SIMUL  S�*�xY�̑a�OBJE�`>̖ADJUS�ݐOAY_IS�D��3����_FI�=��Tu 7�~�6�'���p} =�C�}p�@b�DN��FRIr��T��RO@ \�E}�����OPWOYq�v}0Y�SYSBU/@v�$SOPġd����ϪUΫ}pPRUN,����PA��D���r\ɡL�_OUo��q�$)�IMA�G��w��0P_qIM��L�INv�K�?RGOVRDt�梄X�(�P*�J�|��0L�_�`]��0�RB�1�0��M��E�D}��p ��N�PMdֲ��c�w�SL�`�q�w x $OwVSL4vSDI��DEX����#�$��-�V} *�N4�\@#�B�2�G�B�_�M��y�q�E� �x Hw��p��AT+USW���C�0o��s���BTM�ǌ�I
�k�4��x�԰q�y Dw�E&���@E�r��7��жЗ�EXE��ἱ���8��f q�z @w���3UP'��$�pQ�XN����������� �PG΅{ h? $SUB�����0_���!�MPW�AIv�P7ã�LO�R���F\p˕$R�CVFAIL_C���BWD΁�v��DEFSP!p | Lw���Я�\���UNI+�����bH�R�+�}_L\pAP��x�t���p�}H��> �*�j�(�s`~�NN�`KETB�%�J�PE Ѓ~��J0SIZE	 ��X�'����S�OR��FORMAT�`��c ��WrEM�t��%�U1X��G�G�LI��p��  $ˀP�_SWI�p��J_�PL��AL_ )�����A��B��� uC��D�$E�[�.�C_�U�� � � ����*�J3K0����TWIA4��5��6��MOM�������4��ˀB��AD����؟�����PU� NR ������u��m���� A$PI �6q��	����� K4�)6�U��w`��_SPEEDgPG� �������Ի�4T��� � @��SAMr`��\�]��MOV_�_$�npt5���5���1���2���������'�S�Hp�IN�'�@� +����4($4+T+�GAMMWf�1'��$GET`�p���D�a���

pLIBRt>�II2�$HI=�!_g�t��2�&E;��(1A�.� �&LW�-6 <�)56�&]��v�p���V��$PD#CK���q��_?�����q�&���7����4���9+� ��$IM_SR�pD`�s�rF��r�rLE��¹Om0H]��0����pq��PJqUR_SCRN�FA����S_SAVE_�D��dE@�NOa�C AA�b�d@�$q�Z�I ǡs	�I� �J�K� �� ��H�L��>�"hq ������ɢ��@ bW^US�A���M4���a��)q`� �3�WW�I@v�_�q����MUAo�� � �$PY+�$W�P�vNG�{��P:���RA��RH��RO�PL������q� ��s'�X;�OI�&�Zxe ����m�� p��ˀ�3 s�O�O�O�O�O�aa�_т� |��q�d@ ��.v��.v��d@��[wFv��E���%w�c�tJ;B�w�|�tP���PMA�QUa ���Q8��1�Q�TH�HOLW�Q7HYS��ES��q�UE�pZB��Oτ�  ـPܐ(�A��(��v�!�t�O`�q���u�"���FA��IR#OG�����Q2����o�"��p��INF�Oҁ�׃V����R�vH�OI��� (�0SLEQ������ Y�3����Á��P0QOw0���!E0sNU��AUT�A�COPY�=�/�'��@Mg�N��=�}1h������ ��RG���Á���X_�P��$;ख�`��W��P���@�������EX_T_CYC bH�ȝ�RpÁ�r��_N�Ae!А���R�Ov`	�� � 9���POR_�1�\E2�SRV �)_�6I�DI��T_�k��}�'���dЇ�����5*��6��7��8i�H�iSdB���2�$��)F�p��GPLeAdA
�TAR�Б@����P�2�裔d� �,�0FL`�o@Y�N��K�M��Ck��GPWR+�9ᘐ��ODELA}�dY�p�AD�a�qQSK;IP4� �A�$�-OB`NT����P_$�M�ƷF@\bIp ݷ�ݷ�ݷd���� 빸��Š�Ҡ�ߠz�9��J2R� n��� 4V�EX� TQQ����TQ������� ��`�#�RDCN�V� �`��X)�R�p�����r��m$�RGEAR_� I9OBT�2FLG��fi&pER�DTC����|����2TH2NS�}� 1� ��G T\0 �$��u�M\Ѫ`I�d���EF�1Á�� l�h��ENAB��cTPE�04�]� ���Y�]��ъQn#��@*��"�������2����߼���������3�қ'�9�K�]�o����4�Ҝ����������� N��5�ҝ!�3�E�W�i�{��P��6�Ҟ������P�������7�ҟ@-?Qcu�8�����������SMSKÁ� ��p�0��EkA�QR�EMOTE6������@�݂TQ�IIO}5�ISTP���POW@��� ��pJ����p�����E�"$DSB_S�IGN�1UQ�x�Cx\�TP�S232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+�TQ��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�PHE#�0�����p_XP�C)�$FREEFROMS	pna��GET�0��UPD2�A�2��SP� :�ߧ� !$USAN�na&�����ERI�0�RpRY$q5*"_j@�Pm1�!N�6WRK9KD����6��QFRIEND�Q�RUFg�҃�0oTOOL�6MY�t�$LENGTHw_VT\�FIR�p�C�@ˀE> +IUF�IN-RM��RGyI�1ÐAITI�b$GXñ3IvFG2v7�G1���p3�B�GP1R�p�1F�O_n 0��!RE��p�53҅�U�TC��3A�A�F ��G(��":��� e1n!��J�8�%���%�]��%�� 74�XS O0�L��T�3�H&��8���%b453G�E�W�0�WsR�TD ����T��M����Q�T�]�$V 2�����1�а91�8�02*�;2k3�;3�:i fa�9-i�aQ��NS���ZR$V��2BVwEVP�	V�B;�����& �S�`��F�"�k�@�2�a�PS�E��$pr1C��_$Aܠ�6wPR��7vMU�cS��t '�/89�� 0�G�aV`��p�d`����50�@��-�
25S^�� ��aRW�����B�&�N�A)X�!�A:@LAh�^�rTHIC�1I�8��X�d1TFEj��q>�uIF_CH�3�qaI܇7�Q�pG1Rx�V���]��:�u�_�JF~�PRԀƱ��RVAT��� ���`���0RҦ�DO�fE��COUԱ��A�XI���OFFS=E׆TRIGNS����c����h�����Hx�Y��IGMA0�PA�pJ�E�ORG�_UNEV�J� ��S�����d ӎ$CА�J�GR3OU����TOށ�!DSP��JOG�Ӑ�#��_Pӱ�"O��q����@�&KEPF�IR��ܔ�@M}R&��AP�Q^�Eh0��K�SYS�q"K�;PG2�BRK�B��߄�pY�=�d�����`AD_�����BS�OC���N��DU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR-���C��ˢΓ�OR٧3N]0ڦF��ڦ��OV��SF��p���F+�r!���CC��1q"LCHD}L��RECOVʤc0��Wq@M������#RO�#��Ȑ_+���� @0�e@VER��$OFSe@CV/ �2WD�}���Z2���TR�!|���E_FDO��MB_CM���B��BL�bܒ#��adt�VQR�$0p���G$�7�AM5��� e����_M;��"'����8$CA��'�E�>8�8$HBK(1���IO<�����QPPA������
���������DVC_DBhC;��#"<Ѝ�r!"S�1[ڤ�S�3[֪�/ATIOq 1q� �ʡU�3���CAB Ő�2�CvP��9P^�B��_� �SUBCPU�ƐS�P � M�)0NS�cM�"r�?$HW_C��U���S@��SA�A�pl$�UNITm�l_�A�T���e�ƐCYC=Lq�NECA����FLTR_2_F�IO�7(��)&B�LPxқ/�.�_SCT�CF_`�Fb�l���|��FS(!E�e�CHA��1��4�D°"3�RS�D��$"}����_Tb�PRO����� KEMi_��a�8!�a !�a��D�IR0�RAILAiCI���Mr�LO��C���Qq��#q��V��PR=�S�A�p�C/�c 	��FUsNCq�0rRINP`�Q�0��2�!RAC �B ��[���[gWARn���BL�A�q�A����D�Ak�\���LD@0���Q��qeq�TI"r��K�hPgRIA�!r"AF��Pz!=�;��?,`�R�K���MǀI�!�D�F_@B�%1n�LM��FAq@HRDY4�4_�P@RS�A�0|� �MULSE@x���a ���ưt��m�$�1-$�1$1o������ x*�EaG"p����!AR���Ӧ�09�2,%� 7�wAXE��ROB���WpA��_l-��SY�[�W!‎&S�'WR�U�/-1��@�STRП�����Eb� !	�%��J��AB� ����&9�����OTo0v 	$��ARY�s�#2��Ԓ�	ёFI�@��$LINK(|�qC1�a_�#����%kqj2XYZ@��t;rq�3�C1j2J^8'0B��'�40����+ �3FI���7`�q����'��_Jˑp���O3�QOP_�$2;5���ATBA�2QBC��&�DUβ�&=6��TURN߁"r��E11:�p��9GFL��`_���* �@�5�*7���Ʊ 1�� KŐM��&8���"r��ORQ��a �(@#p=�j�g�#qXUp�����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb��T {�, ��@;�uQ���P \�i��UuQ�We�eL�SERʑe	��!E� O���UdAas���4S�/7����AX��B�'q��E1�e ��i��irp�jJ@�j �@�j�@�jP�j@ �j �!�f��i��i��i ��i��i�y�y��'y�7yTqHyDEBU8�$32����qͲf2G + AB�����رnSVS�7� 
#�d��L�#�L� �1W��1W�JAW��AW� �AW�QW�@!E@?\D2�3LAB�29U�4�Aӏ��C  �o�ERf�5� �� $�@_ A��!�PO��à�0#��
�_MRAt�� �d � T��ٔEcRR����;TY&����I��V�0�cz�TOQ�d�PL[ �d�"ҍ�	��C! � pp`T)0���_V1Vr�aӔ�����2ٛ2�E����@�8H�E���$W���j��V!��$�P@��o�cI��aΣ	 �HELL_CFG�!� 5��Bo_BASq�SR3�\�� a#Sb�T��1�%��2��U3��4��5��6��e7��8���RO�����I0�0NL�\CAqB+�����ACK4� ����,�\@2@�&�?�7_PU�CO. U�OUG�P~ ����m�ذ�����TPհ_KcAR�l�_�RE*��P���|�QUE����uP����CST?OPI_AL7�l��k0��h��]�l0SE�M�4�(�M4�6�T�YN�SO���DI�Z�~�A�����m_T}M�MANRQ���k0E����$KEYSWITCH��ص�m���HE��BE�AT��|�E- LE(~�����U��F!Ĳ�|��B�O_HOM=�OGREFUPPR�&��y!� [�C��O��-ECOC��Ԯ0_IOCMWD
�a���&k��� �# Dh1���UX����M�βgPgCFOR�C�����OM.  �� @�5(�U��#P, 1��, 3���45`P�SNP�X_ASt�� 0Κ�ADD���$�SIZ��$VA�R���TIP/�.��A�ҹM�ǐ���/�1�+ U"S�U!C<z���FRIF��J�aS���5Ԓ�NF�¸�Ѝ� � xp`S�I��TE�C���CSKGL��TQ2�@&������ ��STMTd��,�P �&BWuP���SHOW4����SV�$�� �Q�A00�@Ma}� ��� �����&���U5��6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G ��0G���0G���@�G��PG��1	1�	1	1+	18	1�E	2��2��2��2���2��2��2��2���2��2��2	2�	2	2+	28	2�E	3��3��3��3���3��3��3��3���3��3��3	3�	3	3+	38	3�E	4�4��4��4���4��4��4��4���4��4��4	4�	4	4+	48	4�E	5�5��5��5���5��5��5��5���5��5��5	5�	5	5+	58	5�E	6�6��6��6���6��6��6��6���6��6��6	6�	6	6+	68	6�E	7�7��7��7���7��7��7��7���7��7��7	7�	7	7+	78	7�E��VP��UPD>s�  �`Nм��5�YSLOt�� � L��d���A�aTA�0d��|��ALU:ed�~�CU�ѰjgF!aID_L��ÑeHI�jI��$FILE_���d���$2�fSA>��� hO��`E_BL�CK��b$��hD_CPUyM�yA��cȿo�d��Y����R ;�Đ
PW��!�[ oqLA��S=�8ts�q~tRUN�q st�q~t���qst�q�~t �T��ACC�s��X -$�qLEN;��tH��p�h�_�I��ǀLOWo_AXI�F1�q
�d2*�MZ���ă���W�Im�ւ�aR�TOR��pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v�������TCV��؁��T��ي�����t�V�H���V�Jj�R�MA�"��J��m�u�b����q2j�#�U�{�t�6K�JK��VK;���4H���3��J0�����JJ��JJ��AAAL��ڐ��ڐԖ4Օ5���N1���ʋ�ƀW�LP�_(�g�x,��pr�� `�`�GROUw`��B>��NFLIC��f�REQUIRE3�EBU��qB���w�2����p���q5�p��� \��APP�R��C}�Y�
ްE�N٨CLO7��SC_M��H���u�
�q�u�� ���MCp�����9�_MG��C�Co��`M�в�N�wBRKL�NOL|�tN�[�R��_LIN�H��|�=�J����Pܔ ������������������6ɵ�̲8k�|D����� ���
��q)��7�PATH3�L�B�L��Hôwࡠ�J�CN�CaA�Ғ�ڢB�IN�r�UCV�4a��C!�U�M��Y,���aE��p����ʴ���PA�YLOA��J2L�`R_AN�q�L�pp���$�M�R_?F2LSHR��N�LOԡ�Rׯ�`ׯ�ACRL_G�Œ�ț� ��Hj`߂$yHM���FLEXܣ��qJ�u� :���������0����1�F1�V� j�@�R�d�v�������E����ȏڏ���� "�4�q���6�M���~�@��U�g�y�ယT��o�X��H������藕 ?�����ǟِݕ� ԕ����%�7��P��>J�� � V�h�z���`AT�採@��EL�� S��J�|�Ŝ�JEy�CTYR��~�TN��FQ���HAND_VB�-���v`�� $���F2M����ebS�W�q�'��� '$$MF�:�Rg�(@x�,4�%��0&A�` �=��aM)F�AW�Z`
i�Aw�A��X X�'p�i�Dw�D��Pf�G�p�)STk��!x��!N��DY�pנM�9$ `%Ц�H��H�c�� ����0� ��Pѵڵ����������J��� ���1��Rx�6��QASYMv�����v��J���c���_SH>��ǺĤ��ED����������J��İ%��C�IDِ�_�VI�!X�2PV_UNIX�FThP�J��_R�5_Rc�cTz� pT�V��@���İ�߷�$�U ���������Hqpˢ��aE�N��`DI����O�4d �`J�� x g"IJAA�az�aa bp�coc�`a�pdq�a�� ��OMMEB��� �b�RqAT(`PT�@� S��a7�;�AȠ�@�h�a�iT�@�<� $DUM�MY9Q�$PS�_��RFC�E`$v � ���Pa�� XƠ���ST�E���SBRY�M�21_VF�8$S/V_ERF�O��Ls�dsCLRJtA��O�db`O�p �� D $GLOBj�_LO���u�q��cAp�r�@aSYS��qADR``�`T�CH  � ,x��ɩb�W_NA����7�Ac�TS�R���l  ���
*?�&Q�0"?� ;'?�I)?�Y)��X��� h���x������)��Ռ �Ӷ�;��Ív�?��O�O�O�D�XSCR�E栘p����ST��s}y`����Ea/_HA�q�s TơgpTYP�b����G�aG��Z�Od0IS_��d�UEMd� �Ȁ��ppS�qaRS�M_�q*eUNEX�CEP)fW�`S_ }pM�x���g�z����ÎӑCOU��S�Ԕ �1�!�UE&���Ubwr��PROGM��FL@$CU�gpPO�Q��5�I_��`H� � 8\�� �_HE�PS��#��`RY ?��qp�b��dp�O�US�� � @�6p�v$BUTT�p�RpR�COLU�Mq�e��SERV<5�PANEH�q�� � �@GE�U���Fy��)$�HELPõ)BETERv�)ෆ���A  � ��0��0���0ҰIN簪c��@N��IH�1���_� ֪�L�N�r� �qpձ_�ò=�$H��T�EXl����FLA�@��RELV��DP`��������M��?,�ű�m����"��USRVIE�W�q� <6p�`U:�`�NFI@;��FOCU��;�PR�I@m�`�QY�T�RIP�qm�U9N<`Md� #@pҞ*eWARN)e6�S�RTOL%��g�t�ᴰONCORN��'RAU����T���w��VIN�Le�� $גPATH�9�גCACH��LsOG�!�LIMKR�����v���HOS�T�!�b�R���OBOT�d�I%M>� d�� ����Zq�Zq;�VCPU_AVAIL�V!�EX	�!AN����q��1r��1r��1q �ѡ�p�  #`�C����@$TO�OL�$��_JM�P� ���e�$SS����VS�HIF��Nc�P �`ג�E�ȐR����OSUR��Wk`RGADILѮ��_�a���:�9a��`a�r��L�ULQ$OUTP�UT_BM����I�M�AB �@�rT;ILSCO��C7������� &��3��A���q���m�I�2G�n�y@rMd�}��yDJU��~N�WAIT֖��}��{�%! NE޿u�YBO�� ?�� $`�tv�SB@TPE��NECp�J^FY�.nB_T��R�І �a$�[YĭcB��dM���F� �p�$�pb�OP?�MAS��_DO�!QT�pD��ˑ#%��p!"DELAY�:`7"JOY�@(�nCE$���3@ �xm��d�pY_[�!"�`�"��[����P? АZ�ABC%��  �$�"R��
E`��$$CLAS������!E`4�� � VIRT]��/ 0gABS����1 5�� < �!F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6HpZi{0-�AXL�pt��"�63  �{t�IN��qztPRE������v�p�uLA�RMRECOV c9�rwtNG��� .;	 A �  �.�0PPL�IC��?5�p��Hand�lingTool� o� 
V7.�50P/23-� � �PB��
���_SWt� UPn�!� x�F0���t���A� v�o 864�� �ity�y� N2� 7DA5 j� Q�B@ϐo�Non�eisͅ˰ ���T�]�!LA�Ax>�_l�V��uT��s9�UTO��"�Њt�y��HGA�PON
0g�1��U�h�D 1581����̟ޟry��^��Q 1��� �p�,�蘦���;�p@��q_��"�"� �c�.�H����D�HTTHKYX��"�-�?�Q� ��ɯۯ5����#�A� G�Y�k�}�������ſ ׿1�����=�C�U� g�yϋϝϯ�����-� ��	��9�?�Q�c�u� �ߙ߽߫���)���� �5�;�M�_�q��� �����%�����1� 7�I�[�m�������� ��!����-3E Wi{���� ��)/ASe w����/�� /%/+/=/O/a/s/�/ �/�/�/?�/�/?!? '?9?K?]?o?�?�?�? �?O�?�?�?O#O]����TO�E�W�DO?_CLEAN��7���CNM  � �__/_A_S_��DSPDRYRL�O��HIc��M@�O �_�_�_�_oo+o=o Ooaoso�o�o���pB�F�v �u���aX�t�������9�PLUG�G���G��U�PRC*vPB�@��_�o�rOr_7�SEGF}�K[mwxq�O�O������?rqLAP�_�~q�[�m�� ������Ǐُ�����!�3�x�TOTAL��f yx�USENU
�p�� �H���B���RG_STRIN�G 1u�
��Mn�S5�
~ȑ_ITEM1Җ  n5�� ��$� 6�H�Z�l�~������� Ưد���� �2�D��I/O SI�GNAL̕T�ryout Mo{deӕInp���Simulate�dבOut���OVERR�P �= 100֒I?n cycl��ב�Prog Ab�or��ב��St�atusՓ	Heartbeatї�MH Faul<��Aler'�W� E�W�i�{ύϟϱ������� �CΛ�A ����8�J�\�n߀ߒ� �߶����������"��4�F�X�j�|���WOR{pΛ��(ߎ�����  ��$�6�H�Z�l�~� �������������� 2PƠ�X  ��A{����� ��/ASe�w�����SDEV[�o�#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U?|g?y?PALT� �1��z?�?�?�?�?O "O4OFOXOjO|O�O�O��O�O�O�O�O_�?GRI�`ΛDQ�?_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o�o�o2_l�R��a\_ �o"4FXj| ����������0�B�T��oPREG�>�� f���Ə؏ ���� �2�D�V�h� z�������ԟ���~Z��$ARG_���D ?	����;�� � 	$Z�	[O�]O��Z�p�.��SBN_CONF�IG ;��������CII_S�AVE  Z������.�TCELL�SETUP �;�%HOME_�IOZ�Z�%MO�V_��
�REP��lU�(�UTOBA�CKܠ���FRA:\z�c \�z�Ǡ'`��z���ǡi�INI��0z���n�MESSAG���ǡ|C���ODE_D�������%�O�4�n�P�AUSX!�;� ((O>��Ϟ� �ϾϬ��������� �*�`�N߄�rߨ߶��g�l TSK  �wͥ�_�q�UPDT�+��d!�A�WS�M_CF��;����'�-�GRP Y2:�?� N�BŰ�A��%�XSCRDv1�1
7� �ĥĢ���������� *�������r������� ����7���[�&8�J\n��*�t�G�ROUN�UϩU�P_NA�:�	�t��_ED�1�7�
 �%-BCKEDT-�02�'K�`���Q-t�z�q�q�z���2t1�����q�k�(/��ED3/��/��.a/�/;/M/ED4 �/t/)?�/.?p?�/�/ED5`??�?<?�.�?O�?�?ED6 O�?qO�?.MO�O'O9OED7�O`O_�O�.�O\_�O�OED80L_,�_�^-�_8 oo_�_ED9�_�_]o�_	-9o�oo%oCR_ 9]�o�F�o�k� � NO_�DEL��GE_�UNUSE��L�AL_OUT �����WD_A�BORﰨ~��pI�TR_RTN𷀞�|NONSk����˥CAM_PA?RAM 1;�!��
 8
SON�Y XC-56 �23456789�0 ਡ@����?��( CА\�
���{����^�HR5q�̹���ŏR57ڏ�A�ff��KOWA SC310M
��x�̆�d @<�
���e�^�� П\����*�<���`�r�g�CE_RIWA_I�!�=��F��}�z� .��_LIU�]�����<��FB�GwP 1��Ǯ��M�_�q�0�C*�  ����C1��9J��@��G���CR��C]��d��l��s���R�����[Դm���v���������� C����(��؂��=�HE�`ON�FIǰ�B�G_P_RI 1�{V� ��ߖϨϺ�����������CHKPAU�S�� 1K� ,!uD�V�@�z�dߞ� �ߚ��߾������.�@�R�<�b���O���������_MO5R�� �6��� 	 �����*�@�N�<�������$?��q?;�;����)K��9�P���ça�-:���	�

��M���pU��ð��<��,~��D�B���튒)
m�c:cpmidb�g�f�:�  M#��¥�p�T/���������� �s>ܑ2�3U�V?��p'�p(U�g�/� �����Uf�M/w�O/�
D�EF l��s)��< buf.t�xts/�t/��ާ��)�	`�����=�L���*MC��1�����?43��1���t�īCz � BHH�B�^�B�$�B5��5@@�C����>'�Y
K�D\�nD��C��|@8��.D��� @��=F��&�E�CeE��d�<�X�F��B��IY	X���'w�1����s���.�p���b���BDw�M@x8��K�CҨ����g@D��p@�0EYK�E�X�EQ�E�JP F�E�F� G��>�^F E�� F�B� H,- Ge��H3Y��:��  >�33 ����~  n48�~@��5Y�E>��ðA��Y<#�
�"Q ���+_�'R_SMOFS�p�.�8��)T1��DE 3��F 
Q��;;�(P  B_<_���R����	op6C�4P�Y
s@ ]A(Q�2s@C�0B3�Ma�C{@@*cw��UT��pFPROG !%�z�o�oigI�q����v��ldKEY_TOBL  �&S�#�� �	
��� !"#$%&'�()*+,-./�01i�:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�����������������������p`LCK�l4�p`�`STAT� ��S_AUTO_�DO���5�IN?DT_ENB!���1R�Q?�1�T2}�^��STOPb���TR�Lr`LETE���Ċ_SCREEN� �Zkc�sc��U��MME�NU 1 �Y  <�l�oR�Y 1�[���v�m���̟�� ���ٟ�8��!�G� ��W�i��������ï կ��4���j�A�S� ��w�����迿�ѿ� ���T�+�=�cϜ�s� ���ϩϻ������� P�'�9߆�]�o߼ߓ� ���������:��#� p�G�Y������� ����$����3�l�C� U���y������������ ��	VY)�_M�ANUAL��t�DwBCO[�RIGڇ>
�DBNUM� ���B1 e
�PXW�ORK 1!�[ �_U/4FX�__AWAY�i�/GCP  b=�Pj�_AL� #�j�Yи�܅ `�_�  1}"�[ , 
�@mg�&/~&lMZ��IdPx@P@#ON�TIMه� dɼ`&�
�e�MO�TNEND�o�R�ECORD 1(��[g2�/{�O� �!�/ky"?4?F?X? �(`?�?�/�??�?�? �?�?�?)O�?MO�?qO �O�O�OBO�O:O�O^O _%_7_I_�Om_�O�_  _�_�_�_�_Z_o~_ 3o�_Woio{o�o�_�o  o�oDo�o/�o S�oL�o���� @���+�yV,� c�u��������Ϗ>� P�����;�&���q� ��򏧟��P�ȟ�^� �����I�[�����  ���$�6���������"TOLEREN�CwB���L��Ϳ CS_CFG� )�/'d�MC:\U�L%0?4d.CSV�� �c��/#A ��CH
��z� //.ɿ���(S�RC_OUT *��1/V�?SGN +��"���#�29-J�AN-20 23�:09027l�1�:48+ P;��ɞ�/.��f��pa�m��P�JPѲ��VE�RSION �Y�V2.0.��ƲEFLOGI�C 1,� 	:ޠ=�ޠL���PROG_ENB���"p�ULSk' �����_WRST�JNK ��"fEM�O_OPT_SL� ?	�#
 ?	R575/#=ـ����0�B����TO  �ݵϗ��[V_F EX�d�%���PATH AY�A\������5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAU���z�^"MSWX�.D�<�4,#�Y�/�
!J�6%ZI�~m��$SBL_/FAUL(�0�9'/TDIA[�1<�<�� ���12�34567890
��P��HZl ~������� / /2/D/V/h/�� -P� ѩ�y� �/��6�/�/�/?? /?A?S?e?w?�?�?�?��?�?�?�?�,/�UM�P���� �AT�R���1OC@PME�l�OOY_TEMP?�È�3F���G��|DUNI��.�YN_BRK 2_��/�EMGDI_S�TA��]��ENC2_SCR 3�K7(_:_L_^_l&_��_�_�_�_)��C�A14_�/oo/oAoԢt�B�T5�K�� �o~ol�{_�o�o�o '9K]o�� �������#� 5��/V�h�z��л`~� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T���x���������ү �����,�>�P�b� t���������ο�� ��(�f�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������:� �2� D�V�h�z������ ������
��.�@�R� d�v������������ ��*<N`r ������� &8J\n�� ��������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?��?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O�__NoETMODoE 16�5�QW �d�X
X_�j_|Q�PRROR_PROG %GZ�%�@��_  �UTABLE  G[��?oo)oRjRR�SEV_NUM � �`WP��QQY`�Q_AUTO_ENB  �e�OS�T_NOna �7G[�QXb  �*��`��`��`��`d`+�`�o�o�o�d�HISUc�aOP�k_�ALM 18G[� �A��l�P+ �ok}�����o�_Nb�`  G[�a�R
�:PTCP_�VER !GZ!��_�$EXTLO�G_REQv蜁i\�SIZe�W�T�OL  �aDz�r�A W�_B�WD�p��xf́t�_�DI�� 9�5��d�T�asRֆST�EP��:P�OP�_DOv�f�PF�ACTORY_T�UNwdM�EAT?URE :�5̀�rQHan�dlingToo�l �� \sfm�Englis�h Dictio�nary��rod�uAA Vi�s�� Masteyr����
EN̐�nalog I/yO����g.fd̐�uto Soft�ware Upd�ate  F O�R�matic �Backup��H�596,�gr�ound Edi�tޒ  1 H5�Cameraz�F��OPLGX��ell𜩐II)� X�ommՐsh�w���com��co����\tp���p�ane��  op�l��tyle s�elect��al� C��nJ�Ցon�itor��RDE���tr��Rel�iab𠧒6U�D?iagnos(��^��5528�u���heck Safety UIF���Enhanced� Rob Ser}v%�q ) "S��r�User Fr�[�����a��xt.� DIO �fi�G� sŢ��end�x�Err�LF� IpȐĳr됮� ��  !��FCT�N Menu`�v�-�ݡ���TP I�nېfac�  ER JGC�}pבk Exct��g��H558��i�gh-Spex�S�ki1�  2
�P��?���mmun;ic'�ons��&��l�ur�ې��ST� Ǡ��connz��2��TXPL���ncr�stru�����"FAT�KAREL Cmod. LE�uaG��545\��Runw-Ti��Env���d
!���ؠ+:+�s)�S/W��[��Licens�eZ��� 4T�0�o�gBook(Syvڐm)��H54O�MACROs,\¿/Offse��Loa�MH�������r, k�Mech�Stop Proyt���� lic/�{MiвShif����ɒMixx��)�xSPS�Mod�e Switchn�� R5W�Mo�z:�.�� 74 ����g��K�2h�ulti-T=�M����LN (Po=s�Regiڑ�������d�ݐt Fu�n�ǩ�.�����N�um~����� ln�e��ᝰ Adj�up�����  -{ W��tatuw����T�RDM�z�ot��scove U�9����3Ѓ�uest 4�92�*�o�����6�2;�SNPX b< ���8 J7`����Libr��J�48����ӗ� �Ԅ�
�6�O�� Parts� in VCCMt�32���	�{Ѥ�oJ990��/I�� 2 P��TMI�LIB��H���P��AccD�L�
�TE$TX�ۨ�a�p1S�Te����p�key��wգ�d���Unexc�eptx�motn`Z��������єƉ� O���� 9�0J�єSP CS�XC<�f��Ҟ� �Py�We}���PR�I�>vr�t�m�en�� ��i�Pɰa�����vG�rid�play`��v��0�)�H1��M-10iA(B�201 �2\� �0\k/�Asci�i�l�Т�ɐ/�C�ol��ԑGuar&� 
�� /P-�ޠ�"K��st{Pa�t ��!S�Cyc8�҂�orie�⑻IF8�ata- q�uҐ�� ƶ��mH�574��RL��a�m���Pb�HMI De3�(b�����PCϺ�Passswo+!��"PE? cSp$�[���tp��.� ven��Tw�N��p�YELLOW� BOE	k$ArcN��vis��3*��n0WeldW�ci�al�7�V#t�O�p����1y� 2zF�a�portN�(�p�T1�T� ��� ��xy]�&TX��tw�igj�1� �b� ct\�JP�N ARCPSU� PR��oݲOL�� Sup�2fil� &PAɰאcro�� "PM(�����O$SS� eвte�x�� r���=�t��ssagT��P��P@�Ȱ�锱��rtW��H'>r�dspn��n1
t��!� z ��asc�bin4psyn���+Aj�M HE�L�NCL VI�S PKGS PwLOA`�MB ��,�4VW�RIP�E GET_VA�R FIE 3\�t��FL[�OOL�: ADD R7�29.FD \j�8'�CsQ�QE��D�VvQ�sQNO W�TWTE��}PD � �^��biRFO;R ��ECTn�`���ALSE AL�AfPCPMO-1�30  M" #�h�D: HANG FROMmP�AQ�fr��R709 �DRAM AVA�ILCHECKS�O!��sQVPCS �SU�@LIMCH�K Q +P~dFF �POS��F�Q R�5938-1?2 CHARY�0�PROGRA �W�SAVEN`AM]E�P.SV��7��$En*��p?FU�{��TRC|� SHA�DV0UPDAT �KCJўRSTAT�I�`�P MUCH� y�1��IMQ �MOTN-003���}�ROBOGU�IDE DAUG�H�a���*�tou�����I� Šhd�A�TH�PepMOVE�T�ǔVMXPA�CK MAY A�SSERT�D��Y�CLfqTA�rBE COR vr*Q�3rAN�pRC O�PTIONSJ1v�r̐PSH-17�1Z@x�tcǠS�U1�1Hp^9R!�Q�`_�T�P��'�j�d�{tby app �wa 5I�~d�PHqI���p�aTEL��MXSPD TB$5bLu 1��UB6@�q�ENJ`CE2�61ꏠp��s	�mayc n�0� R6{��R� �Rtraff\)�� 40*�p���fr��sysva�r scr J78��cj`DJU��b�H V��Q/�PSE�T ERR`J` �68��PNDAN�T SCREEN? UNREA��'�J`D�pPA���pR�`IO 1���PF�I�pB�pGROUN�PD��G��R�P�Q>nRSVIP !p�a��PDIGIT VgERS�r}BLo�U�EWϕ P06 9 �!��MAGp�abZV�DI�`� �SSUE�ܰ�EPLAN JOT`O DEL�pݡ#Zz�@D͐CALLOb��Q ph��R�QIwPND��IMG��R719��MNT]/�PES �pVL�c��Hol�0Cq��N�tPG:�`C�M��canΠ��pg.�v�S: 3D m~K�view d�`� �p��ea7У�b�� of �Py���A�NNOT ACCESS M��Ɓ*��t4s a��lo�k��Flex/:ڈRw!mo?�PA�?�-�����`n�pa� SNBPJ AUTO-�06f�����TB��PIABLE�1q 636��PLgN: RG$�pl;p�NWFMDB�VI|���tWIT 9x�:0@o��Qui#0�Ҿ�PN RRS?pU�SB�� t & _remov�@ )��_��&AxEPFT_f=� 7<`�pP:�OS-144 ���h s�g��@OS�T� � CRAS�H DU 9���$P�pW� .$���LOGIN��8�&�J��6b046 �issue 6 �Jg��: Slo�w �st��c (Hos`�c���`�IL`IMPRWtS?POT:Wh:0�T�STYW ./�V�MGR�h�T0CA]T��hos��E�q���� �O�S:N+pRTU' k�-S�Y ����E:��pv@8�2�� t\hߐ��9m ��all��0�s  $�H� WA͐���3 CNT0 �T�� WroU�a�larm���0s�d � �0SE1���r R{�OMEBp���nK� 55��REà�SEst��g   �  �KANJ�I�no���IN�ISITALIZ-p�dn1weρ<���dr�� lx`�S�CII L�fa_ils w�� ��`�YSTEa���o���Pv� IIH���1�W�Gro>Pm ol\wpSh@�P��~Ϡn cflxL@�АWRI �OF �Lq��p?�F�up���de-rela��d "APo S�Y�ch�Abetw}e:0IND t0�$gbDO���r� �`�GigE�#operabilf  PAbHi�H`��c��lead�\et�f�Ps�r�OS p030�&: fig��GLA )P ��i����7Np tpswZx�B��If�g�������5aE�a E�XCE#dU�_�tPC�LOS��"robV�NTdpFaU�c��!���PNIO /V750�Q1��Q�a��DB ��P �M�+P�QED�DEyT��-� \rk���ONLINEhSBUGIQ ߔĠi`Z��IB�S apABC JARKYFqr� ���0MIL�`*� R�pNД �p0WGAR��D*pRМ�P�"! jK�0cT��P�Hl#n�a�ZE� V�� TASK�$VP2(�4`
�!p�$�P�`WIBPKk05�!FȐB/���BUSY RUNN�� "�򁐈���R-p�LO�N�D;IVY�CUL��gfsfoaBW� p���30	V��ˠ�IT`�a505.��@OF�UNEXH�P1b�af�@�E���SVEMG� NM�Lq� D0pCC_�SAFEX 0c�08�"qD �PET�`N�@�#J87����RPsP�A'�M�K�`�K�H GUNC{HG۔MECH�p�Mc� T�  y,� g@�$ ORY LEAKA�;�ޢGSPEm�Ja��V�t�GRIܱ�@�C7TLN�TRk�Fp�epR�j50�ENF-`IN�����p �`0�Ǒk!��T3/dq.o�STO�0A�#�L�p �0�@�Q�АaY�&�;pb1TO8pP�s���FB�@Yp`&�`DU��aO�sup$k�t4 � P�F� B�nf�Q�PSVGN�-1��V�SRSR)J�UP�a2�Q�#<D�q l O��Q?BRKCTR5Ұ��|"-�r�<pc�j!I{NVP�D ZO� ���T`h#�Q�cHse�t,|D��"DUA�L� w�2*BRVO_117 A]�TN�p�t�+bTa2473�0�q.?��sAUz�i��B�complet�e��604.�{ -�`hanc�U� F��e8��  ��npJtPd!q�ܱ`��� 5h59	6p�!5d�� "p�P�P�Q�0�P2�p�A� HxP��R(}\xPe� %aʰI���E��1���p� j  �� xSPO�^P �A�AxP��q 5 sig��a��"AC;a��
��bCexPb_p��.�pc]l<bHbcb_�circ~h<n�`tl1�~`xP`o�dxP�b,]o2�� �cb�c�i|xP�jupfrm�d8xP�o�`exe�a�o<FdxPtped}o��|u`�cptlibxzxP�lcr�xrxP\blsazEdxP_fm�}gcxP�x���o|�sp�o�mc(��ob_�jzop�u6�wf(��t��wms�1q��csld�)��jmc�o�\�n��nuhЕ��|s1t�e��>�pl�qp��iwck���uvf�0uߒ��lvisn��CgaculwQ
}E F  ! Fc�.fd�Qv�� q�w���Data A�cquisi��nxF�|1�RR631`���TR�QDMCM Z�2�P75H�1�P�583xP1��71֫�59`�5�P57@<PxP�Q����(����Q��o pxP!daq\�oA��@��� ge/�etdm~s�"DMER"؟�,�pgdD���.�mp���-��qaq.<ጡ�xPmo��h���f�{�u�`13��MACROs, SksaCff�@z����03�SQR�Q(��Q6��1�Q9ӡ�R�ZSh��PxP�J643�@7ؠ6X�P�@�PRS�@����e �Q�UС PIK��Q52 PTLC��W��xP3 (��p/O��!�Pn ��xP5��03\sf�mnmc "MNCMCq�<��Q��\$AcX�FM���ci,� ��X����cdpq+�
�sk�SK�xP�SH560,P��,��y�refp "R#EFp�d�A�jxP	�of�OFc�<gy�to�TO_���������+je�u>��caxis2�xP�E�\�e�q"ISD�Tc��]�prax ��MN��u�b�isde܃h�\�w��xP! isbaskic��B� P]�ޔQAxes�R6p������.�(Ba�Q�ess��xP����2�D�@�z�atis���(�{�����4~��m��FMc�u�x{�
ѩ�MNIS�� ݝ����x����ٺ���x� j75��D�evic�� In?terfac�R��QJ754��� xP�Ne`��xP����2�б����dn� "DNE���
�tpdnui5U1I��ݝ	bd�bP|�q_rsofO�b
dv_aro���u�����stchkc��z	 �(}onl��G!ffL+H�J(��"l"/�n�b��z�Ohamp��T�C�!i�a"�59��S�q��0 (�+P�o�u��!2��xpc_2pc�chm��CHMP8_�|8бpevws��8�2쳌pcsF��#�C SenxPac�ro�U·�-�R6 �Pd�xPk�����p��qgT�L��1d M�2 `��8�1c4ԡ�3 q;em��GEM,\i|(��Dgesnd�5����H{�}Ha�@sy���c�Isu�xD��Fmd��I��7�4����u���AccuCaAl�P�4� ��ɢ7ޠ�B0��6+6f�6���99\aFF q�S( �U��2�
X�p�!�Bd��cb_�SaUL��  �� ?�ܖ�to��otplu?s\tsrnغ�qb�Wp��t���1���Tool (N. A.)�[K�7�Z�(P�m����b�fcls� k94�"�K4p��qtpap� "PS9H�stpswo��p�L7��t\�q����D� yt5�4�q��w�q���� �M�uk��rkey����s��}t�s�featu6�EA��� cf)t\Xq������d�h5���LaRC0�md�!�587���aR�(����2V���8c?u3l\�pa3}H�&r-�Xu���1t,�� �q "�q�O t��~,���{�/��1c�}����y�p�r�� 5���S�XAg�-�y��ށWj874�- �iRVis���Queu�� Ƒ�-�6�1���(����u����tӑ����
�t�pvtsn "V�TSN�3C�+�� v�\pRDV����*�p�rdq\�Q�&�vstk=P�������nm&_�դ�clrqqν���get� TX��Bd���aoQϿ�0qstr�D[� ¡�t�p'Z����np8v��@�enlIP0���D!x�'�|���sc ߸��tvo/��2�q���vb���� q���!���h]��(�� Contro�l�PRAX�P5ξ�556�A@59��P56.@56@5�A�J69$@98�2 J552 IDVR7�hqA���16��H���La��� ��Xe�frlp�arm.f�FRL�am��C9�@(F�����w6{��x�A��QJ643��� 50�0LSE�
_pVAR $S�GSYSC��RS_UNITS �P�2�4tA�TX.$�VNUM_OLD� 5�1�xP{�5�0+�"�` Funct���5tA� }��`#@�`3�a0�cڂ��19���@H5נ� �P���(�A���� ۶}����ֻ}��bcPRb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`d���1���96������%C�� Aف��J�bIncr�	�����\���1o5qn=i4�MNINp	xP��`���!��Hour  �� 2�21 �AAVM����0 ��TUP ���J545 ���6162�VCAM  (�CLIO ��R6�N2�MgSC "P �?STYL�C��28~ 13\�N�RE "FHRM� SCH^�D�CSU%ORSR� {b�04 ��EIOC�1 j� 542 � os�| � egistP�����7�1��MASK�9�34"7 ��OCSO ��"3�8�b�2���� 0 HBh��� 4�"39N�� Re�� �LC{HK
%OPLG%z��3"%MHCR.%�MC  ; 4? ��6m dPI�54�sn� DSW%MD� 9pQ�K!637�0�0dp"�1�Р"4 ��6<27 CTN �K � 5 ���"7���<25�%/�T�%F'RDM� �Sg!��930 FB( N�BA�P� ( HLB�  Men�SMx$@jB( PVC ���20v��2HTC��CTMIL���\@PAC 16�U�hAJ`SAI \@E�LN��<29s��UECK �b�@FgRM �b�OR����IPL��Rk0C�SXC ���VV�FnaTg@HTTP9 �!26 ���G�@obIGU=I"%IPGS�r� H863 qb�!�0�7r�!34 �r�84 \so`! Qx`&CC3 Fb�21�!�96 rb!51 L���!53R% 1!Qs3!��~�.p"9js� VATFUJ77Q5"��pLR6^RP�wWSMjUCTO�@bxT58 F!80����1XY ta3!77s0 ��885�UOL  GTSo
�{`� LCM �r| T3SS�EfP6 W�\@�CPE `��0V1R� l�QNL"��@�001 imrb�c3 =�b�0���0ƒ`6 w�b-P- �R-�b8n@5EW�b9 �Ґa� ���b��`ׁ�b2 200I0��`3��`4*5��`5!�c�#$�`7�.%�`8 h605v? U0�@B6E"a�Rp7� !Pr8 �t�a@�tr2 i�B/�1vp3�vp5I Ȃtr9Σ�a4@9-p�r3 F��r�5&�re`u��r7 ���r8�U�p9 \�h738�a�R2�D7"�1f��2�&�7� �3 7iC��4>w5Ip�Or'60 C�L�1bEN�4 I�pyL�uPИ�@N�-PJ8�N�8NeN�9 H�r`�EE�b7]�|���8���ࠂ9 2��a`�0�qЂ5�%U09'7 0��@1�0����1 (�q�3 5R���0���mp U��0�0�7*��H@(q�\P"RB6�q124�b;��@����@06� x�3 �pB/x�u ��x�6_ H606�a1� <��7 6 ��x�p�b155 �����7jUU162 L�3 g��4*�65 2e "_���P�4U1`���B1����`0'�174 �q��P�E186 3R ��P�7 ��P��8&�3 (�907 B/�s191���Θ@202��6 a3���A�RU2� <d��2 b2h`���4�᪂2�4���1I9v Q�2��u2d��Tpt2� ��H�a2�hP�$�5���!U2��p�p
�2�p��@5��0-@��8 @�9F��TX@�� �e5�`'rb26Af�2^R�a@�2Kp��1y�b5Hp�`
�5�0@�gqGA����a52ѐ�Ḳ6��60ہ5� ׁ2Ҹ�8�E��9�EU5@ٰ\�q5hQ`S�2ޖ5�p\w�۲�p�J �-P��5�p1\�t�H�4��PCH�7j��phiw�@��P��x��559 ld u� P�D���Q�@������� �`.��P>�8�581�"�q5�8�!AM۲T�A ;iC�a589��@�x����5 �a��1�2׀0.�1���,�2p����,�!P\h8��RLp ��,�7��6�0�840\��ANRS 0C}A��p���{��ran��FRA��Д�е���A %���ѹ�Ҍ����� (����Ќ���З� ��������ь����B$�G��1��ը���������� x9S�`q�  ������`64��M��iC?/50T-H����0��*��)p46��� �C��N����m75s֐� Sp��b�46��v����ГM-71?�7�З����42������C��-�а�70�r�	E��/h����O�$��rD���c7c7�C�q��Ѕ���L���/��2\imm7c7�g������`���(��e��� ��"�������a �r��c�T,�Ѿ�" ��,�� ��x�Ex�m77t����k����5�����)�iC��-HS-� B
�_�>���+�Т�7@U�]���Mh7��s��7������-�9?�/260L_@������Q����h���]�9pA/@����q�S�хx���h621��c��92������.�)92c0�g$ �@�����)$��5$���pylH"O"
�2�1���t?�350 ����p��$�
�� �350!����0��9�U/0\m=9��M9A3��(4%� s��3M$���X%u���"him9@8J3����� i d�"m4~�103p�� ����h794̂�&R���H�0����\��� g�5AU��՜��0���*2��00��#06��АՃ�է!07{r ��������k�@�@����EP�# ������?��#!��;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?�ҽCD�25L����0:�"l�2BL
#��B��\20�2_�r�r e���X��1��N���H�A@��z��`C�p`U��`��04��$DyA�\�`fQ���sU���\�5  ���� p�3^P��<$85����+P=�ab1l��1#LT��lA8�!uD�nE(�20T��J8�1 e�bH85���b4�Ռ�5[�16Bs ��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3�  ��b�s��-`�_W8�_����6Id	$�X5�1�U85��R�p6S����/�/ +q�!�q��`�6o��q5m[o)�m6sW���Q�?��set0�6p ��3%H�5��10p$����g/�Jr�H��  ��A�856����F2�� ���p/2��h� ��܅�✐)�5��̑`v��(��m6��BY�H�ѝ̑m�6�Ҕ���a6�DM����-S�+��H2���� �Ҽ�� �r̑���`����l���p1����F���2�\t6h T6H����Ҝ� 'Vl���ᜐ�V7᠜�/����;3A7���p~S��������4��`圐�V���!3
��2�PM[��%ܖnO�chn��vel5�����Vq���_ar�p#��̑�.���2l_hemq$�.�'�6415���5���?�@���F�����5g�L�ј[���1����1����M7NU��М��eʾ����u"q$D;��-�4��3&H�f�c�Ĝ�h���� ��u���㜐���ZS�!ܑ4���M-����S�$̑�ք �� 0��<�����07shJ�H�v�À� sF��S*󜐳���̑@���vl�3�A�T�#���QȚ�Te��q�prX����T@75j�5�d d�̑1�(UL�&�(�,����0�\�?���̑�a�� xSP���a�e�w�2��(�	�2�C��A/���\��+p�����21 (ܱ�CL S���� B̺��7F���?�<�lơ1L����c� Č��u9�0����e/q��O���9�K��r9 (��,�Rs����5�G�m20c ��i��w�2��:�0`�$��2�2l�0�k� X�S� ,�ι2��O�4��1!41w���y2T@� _std��G�y� �ң�H� jdgm����w0\�  �1L���	�P�~�W*�b��t 5�����J�3�,���E{�������L��5	\L��3�L�|#~���~!���4�#��O����h�L6A��������2璥���4�4�����[6\j4s��·���#��ol�E"w�8Pk����� ?0xj�H1�1Rr�>�l�]�2a�2Aw�$P ��2��|41�8�� ˡ��{� �%�A<��� +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K� R��ˑb�W���Fs� ��)�ѐ�!���a�1�����5��16�1�6C��C����0\imBQ��d����b���\B5�-���DiL���O�_�<ѠPEtL�E�RH�ZǠPg���am1l��u��� ̑�b�<����<�$�T�̑�F����Ȋ�Dpb��X"��hr���p� ���^P��9�0\� j97�1\kckrcf�J�F�s�����c��e? "CTME�r����ɛ��a�`main�.[��g�`run}�_vc�#0�w�1�Oܕ_u����bct�me��Ӧ�`ܑ�j�735�- KA�REL Use {�U���J��1���p� Ȗ�9�B@@��L�9��7j[��atk208 "�K��Kя��\��9���a��̹����cK�RC�a�o ��kc �qJ�&s�����Grſ �fsD��:y��s�ˑf1X\j|хrdtB�2, ��`.v�q��� �sǑIf�Wfj5�2�TKQuto �Set��J� H�5K536(�93�2���91�58(�94�BA�1(�74O,A~$�(TCP Ak����/�)Y� �\�tpqtool.�v��v���! c�onre;a#�Co�ntrol Re�ble��CNRE(�T�<�4�2���D�8)���S�552��q(g�� (򭂯4X��cOux�\sfuts�UTS`�i������t�棂��? q6�T�!�SA OO+D6���������,!��6c+� i\gt�t6i��I0�TW8 ���la��vo58�o�bFå��i�Xh��!Xk�0Y�!8\m6e�!6#EC���v��6���� �����<16�A���A�6s����U�g˰T|ώ���r1�qR��˔Z4�T�����,#�eZp)g����@<ONO0���uJ��tCR�;��F�a� xSP��f��prdsuc#hk �1��2&&?���t��*D%$�r(��✑�娟:r��'�sp�qO��<scrc�xC�\At�trldJ�"o�\�V����P�aylo�nficrm�l�!�87��@7��A�3ad� ! �?ވI�?plQ��3��3"�q��x pl�`���d7��l�calC�uDu���;��mov�����OinitX�:s8O���a�r4 ��r67�A4|�e Gene�ratiڲ���7�g2q$��g R� G(Sh��c ,|�"bE��$Ԓ\�(:�"��4��4�4�. sg��5�F$d�6"e;Qp "S�HAP�TQ ngcr pGC�a(�&x"� ��"GDA¶&��r6�"aW�/�$dataX:s�"�tpad��[q�%tput;a__O7;a�Po8�1�yl+s�r�?��:�#�?�5x�?�:c O�:y O�:�IO�	s`O%g�qǒ�?�@p0\��"o�j92;!��Ppl.Coll{is�QSkip#� �@5��@J��D��@\�ވ�C@X�7��7��|s2��ptcl�s�LS�DU�k<?�\_ ets�`�< \�Q��@���`2dcKqQ�FC;��1J,�n��` (��"4eN����T�{�� �'j(�c�����/I��aȁ��̠H������зa�e\m�cclmt "C�LM�/��� mat�e\��lmpALaM�?>p7qmc?����2vm�q��%�3s���_sv90�_x_Gmsu�2L^v_� K�o�{in�8(3r><�c_logr���rtrcW� "�v_3�~yc���d�<�te��de�r$cCe� Fiρ�R��Q�?�>l�enter߄|���(Sd��1�TXj�+fK�r�a99sQ�9+�5�r\tq~\� "FNDR�}��STDn$�LANG�Pgui��D⠓�S�������sp�!ğ֙uf�ҝ�s����$�����e+�=����������������w�H�r\�fn_�ϣ��$`x�t�cpma��- T�CP�����R63�8 R�Ҡ��38��M7p,���Ӡ� $Ӡ�8p0Р�VS,�>�tk��99�a��B3 ���PզԠ��D�2�����UI��t���hqB� ��8��������p����re�ȿ��exe @4φ�B���e38�ԡ�G�rmpWXφ�var@�φ�3N��ψ��vx�!ҡ��q��RBT $c�OPTN ask� E0��1�R M{AS0�H593/՟96 H50�i�480�5�H0��mԢQ�K��7�0�g�P�l�h0ԧ�2�OR�DP��@"��t\mas��0�a��"��������k�գR�����ӹ`m��b��7�.If��u�d��r��splayD�E���|1w�UPDT Ub���887 (��D	i{���v�Ӛ�Ԛ‧���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q`�䗣�#��К�`2�� vlv������$�>�b���! <S��Easy/К�Util��룙�5�11 J�����R�7 ��Nor֠��i�nc),<6Q�� ��`c��"4�[���9�86FVRx So����q�nd6����P ��4�a\ (��
  ��������d��K�bd�Z���men7���-7 Me`tyFњ�Fb�0�TUa�577?i3R��\�5�u?��!� �n���f������l\mh�Ц�űE|�hmn�	��<\�O���e�1�� �l!��y��Ù�\|p����B���Ћmh�@��:.a G!���/�t�55�6�0�!X�l�.us��Y/>k)ensubL���eK�h�� �B\1 ;5g?y?�?�?D��?*�rm�p�?Ktbox O2K|?�G��C?�A%ds���?1ӛ#� �TR��/��P�4B �`�U�P�V�P"�Q�P�0�U�PO��P�"�T3��U�P�f�Pk"�2}�4��T�P�f�P2�"�Q5 �S�Q���R?Ă�Q3t.�P׀al��P+�OP517��IN0a��Q(}g��P'ESTf3ua�PB�l�ig�h�6�aq��P � xS�΅`  n�0mbusmpP�Q969g�C69�Qq��P0�ba�Ap�@Q� BOX8��,>vche�s��>vetu㒣=wffse�3���]�`;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q<twaNǂ tp�Q҄Ta�ror Reco�v�b�O�P�642����a�q��a�f�QErǃ�Qry���`�P'�T�`�aar�������	{'�pak971��71��m���>�pjot��PXch��C�1�adb -�a;il��nag���b�QR629�a�Q����b�P  �
�  �P��$$�CL[q ����������$��PS_DIGIT\���"� !�4�F�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv�����@��*璬1�:PRODUCT��Q0\PGSTK�bV,n�99��\���$F�EAT_INDE�X��~��� 搠ILEC�OMP ;���)��"��SET�UP2 <����  N �!�_AP2BC�K 1=� G �)}6/E+%,/i/��W/�/~+/ �/O/�/s/�/?�/>? �/b?t??�?'?�?�? ]?�?�?O(O�?LO�? pO�?}O�O5O�OYO�O  _�O$_�OH_Z_�O~_ _�_�_C_�_g_�_�_ 	o2o�_Vo�_zo�oo �o?o�o�ouo
�o. @�od�o��� M�q���<�� `�r����%���̏[� ������!�J�ُn� ������3�ȟW���� ��"���F�X��|�� ��/���֯e������ 0���T��x������ =�ҿ�s�ϗ�,ϻ��9�b�� P/ }2) *.VRi���!�*����������PC�7�!��FR6:"�c��χ��T��߽�L�����ܮx���*#.F��>� �	N�,��k��ߏ��STM� �����Qа����!�iPenda�nt Panel���H��F���4���8���GIF��������u����JPG&P��<�����	PANEL1'.DT��������2�Y� G��
3w�@����//�
4��a/�O///�/�
�TPEINS.XSML�/���\�/��/�!Custom� Toolbar�?�PASSW�ORD/�FR�S:\R?? %�Password Config�? ��?k?�?OH�6O�? ZOlO�?�OO�O�OUO �OyO_�O�OD_�Oh_ �Oa_�_-_�_Q_�_�_ �_o�_@oRo�_voo �o)o;o�o_o�o�o�o *�oN�or�� 7��m��&�� �\�����y���E� ڏi������4�ÏX� j��������A�S�� w�����B�џf��� ����+���O������ ���>�ͯ߯t���� '���ο]�򿁿�(� ��L�ۿpς�Ϧ�5� ��Y�k� ߏ�$߳�� Z���~�ߢߴ�C��� g�����2���V��� �ߌ���?����u� 
���.�@���d���� ��)���M���q��� ��<��5r�% ��[�&� J�n��3� W���"/�F/X/ �|//�/�/A/�/e/ �/�/�/0?�/T?�/M? �??�?=?�?�?s?O �?,O>O�?bO�?�OO 'O�OKO�OoO�O_�O :_�O^_p_�O�_#_�_ �_Y_�_}_o�_�_Ho�)f�$FILE_�DGBCK 1=���5`��� ( �)�
SUMMARY�.DGRo�\MD�:�o�o
`Di�ag Summa�ry�o�Z
CONSLOG�o�o�a
�J�aConso?le logK�[��`MEMCHECCK@'�o�^q�Memory D�ata��W��)�qHADOW����P��sSh�adow Cha�ngesS�-c-��)	FTP=Ъ�9����w`qmment TBD׏��W0<�)ET?HERNET̏�^��q�Z��aEth�ernet bpf�iguratio�n[��P��DCSV�RFˏ��Ïܟ�q�%�� veri?fy allߟ-c�1PY���DIF�Fԟ��̟a��p%=��diffc����q��1X�?�Q��c ����X��CHGD��¯ԯi�B�px��� ���2`�8G�Y�� ��� �GD��ʿܿq��pq���Ϥ�FY3h�8O�a��� ��(�GD������y��p��ϡ�0�UPDATES.�Ц��[?FRS:\������aUpdate?s List���k�PSRBWLD.CM.��\��B���_pPS_ROBOWEL���_����o ��,o!�3���W���{� 
�t���@���d��� ��/��Se��� ��N�r�  =�a�r�&� J���/�9/K/ �o/��/"/�/�/X/ �/|/�/#?�/G?�/k? }??�?0?�?�?f?�? �?O�?OUO�?yOO �O�O>O�ObO�O	_�O -_�OQ_c_�O�__�_ :_�_�_p_o�_o;o �__o�_�o�o$o�oHo �o�o~o�o7�o0 m�o� ��V� z�!��E��i�{� 
���.�ÏR������� ���.�S��w���� ��<�џ`������+� ��O�ޟH������8�ຯ߯n����$FoILE_��PR����������� �MDO?NLY 1=4��? 
 ���w� į��诨�ѿ������ �+Ϻ�O�޿sυ�� ��8�����n�ߒ�'� ��4�]��ρ�ߥ߷� F���j�����5��� Y�k��ߏ���B��� ��x����1�C���g� �����,���P����� ����?��Lu�?VISBCKR�<�>a�*.VD|�>4 FR:\���4 Visio�n VD file� :LbpZ �#��Y�}/ $/�H/�l/�/�/ 1/�/�/�/�/�/ ?�/ 1?V?�/z?	?�?�??? �?c?�?�?�?.O�?RO dOO�OO�O;O�O�O qO_�O*_<_�O`_�O��__%_�_�MR_�GRP 1>4��L�UC4  B�P	 ]�ol�`�*u����RHB ���2 ��� ��� ���He�Y�Q `orkbIh�oJd�o�S�c�o�oO\ ��M��7L[��F�5U�aT>��x�o�o A��B�-\A��.�Q6���;�o%F}?RU\�?W�lq�Q?V�o<xq}E�� F@ �r�d�a}�J��NJk��H9�Hu���F!��IP�s�X~�`�.9�<�9�89�6C'6<,�6\b�  A�/�-BHr!Aw�a�0���� ��  @�6�%&]�Ay;0���� H���,>p1������ |�ݏx���%��vp��A6Β@U��{�v�a����� ��П����ߟ��<��'�hzBH�P ��a`�Q��Q= �K���ï�T
6�P;�uP=�f˯`�o�e�Q cB��P<5���@�33@����4�m�,�@UUU�U�~w�>u.�?!x�^��ֿ����3��=[z��=�̽=V6�<�=�=��=$q��~��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�Ϡ Cϫo��C�
�P��P'�6��_V�  m�o��To��xo�ߜo ������A�,�e�P� b���������� ���=�(�a�L���p� ��������>p������ *��N9r]�� ������8 #\nY�}�� �����/ԭ//A/ �e/P/�/p/�/�/�/ �/�/?�/+??;?a? L?�?p?�?�?�?�?�? �?�?'OOKO6OoO�O HߢOl��ߐߢ��O��  _��G_bOk_V_�_z_ �_�_�_�_�_o�_1o oUo@oyodovo�o�o �o�o�o�oN u����� ����;�&�_�J� ��n�������ݏȏ� �%�7�I�[�"/�� ������ٟ������� 3��W�B�{�f����� ��կ�������A� ,�e�P�b��������O �O�O��O�OL�_ p�:_�����Ϧ����� ���'��7�]�H߁� lߥߐ��ߴ������� #��G�2�k�2��V w�����������1� �U�@�R���v����� ��������-Q �u���r��6 ��)M4q \n������ /�#/I/4/m/X/�/ |/�/�/�/�/�/?ֿ �B?�f?0�BϜ?f� �?���/�?�?�?/OO SO>OwObO�O�O�O�O �O�O�O__=_(_a_ L_^_�_�_�_���_�� o�_o9o$o]oHo�o lo�o�o�o�o�o�o�o #G2kV{� h������� C�.�g�y�`������� ���Џ���?�*� c�N���r�������� ̟��)��M�_�&? H?���?���?�?�?�� ��?@�I�4�m�X�j� ����ǿ���ֿ��� �E�0�i�Tύ�xϱ� ����������_,��_ S���w�b߇߭ߘ��� ��������=�(�:� s�^��������� ��'�9� �]�o��� ��~����������� ��5 YDV�z ������1 U@yd��v� ����/Я*/��
/ �u/��/�/�/�/�/ �/�/??;?&?_?J? �?n?�?�?�?�?�?O �?%OOIO4O"�|OBO �O>O�O�O�O�O�O!_ _E_0_i_T_�_x_�_ �_�_�_�_o�_/o�� ?oeowo�oP��oo�o �o�o�o+=$a L�p����� ��'��K�6�o�Z� �����ɏ��폴�  ��D�/ /z�D/�� h/ş���ԟ���1� �U�@�R���v����� ӯ������-��Q� <�u�`���`O�O�O�� �޿��;�&�_�J� oϕπϹϤ������ ��%��"�[�F��Fo �ߵ����ߠo��d�!� ��W�>�{�b��� ������������A� ,�>�w�b����������������=���$FNO ����\_�
F0l q � FLAG>�(�RRM_CHKT_YP  ] ���d �] ��O=M� _MIN� 	����� �  �XT SSB_CF�G ?\ �����OTP_DEF_OW  	���,IRCOM�� >�$GENO�VRD_DO���<�lTHR� �d�dq_ENB�] qRAVC_GRP 1@�I X(/ %/ 7//[/B//�/x/�/ �/�/�/�/?�/3?? C?i?P?�?t?�?�?�? �?�?OOOAO(OeOpLO^O�OoROU��F\� ��,�B,�8�?����O�O�O	__���  DE_�Hy_�\@@m_B�=�vR/���I�O�SMT�G��SUoo&oRHoOSTC�1H�I�� ��zMS5M�l[bo�	127.0�`=1�o  e�o�o �o#z�oFXj�|�l60s	ano?nymous��0�����iao�
&�&��o�x��o ������ҏ�3�� ,�>�a�O�������� ��Ο�U%�7�I��]� ���f�x�������� ү����+�i�{�P� b�t���������� ��S�(�:�L�^ϭ� oϔϦϸ������=� �$�6�H�Zߩ���Ϳ s����������� � 2���V�h�z��߰� ��������
��k�}� �ߡߣ���߬����� ����C�*<Nq� _������-� ?�Q�c�eJ��n� ������/ "/E�X/j/|/�/�/ �%'/?[0? B?T?f?x?��?�?�? �?�??E/W/,O>OPO�bO�KDaENT 1=I�K P!�?�O  �P�O�O�O �O�O#_�OG_
_S_._ |_�_d_�_�_�_�_o �_1o�_ogo*o�oNo �oro�o�o�o	�o- �oQu8n�� ������#�� L�q�4���X���|�ݏ ���ď֏7���[����B�QUICCA0��h�z�۟��1ܟ��ʟ+���2,����{�!ROUTE�R|�X�j�˯!P�CJOG̯��!�192.168�.0.10��}GN�AME !�J!?ROBOT�vN�S_CFG 1H��I ��Auto-sta�rted�$FTP�/���/�?޿#? ��&�8�JϏ?nπ� �Ϥ�ǿ��[������"�4�G�#������� �������������� ��&�8�J�\�n��� �����������/�/ �/F���j��ߎ����� ��������0S� T��x����� !�3��G,{�Pb t��C���� /�:/L/^/p/�/ ���	/�/=? $?6?H?Z?)/~?�?�? �?�/�?k?�?O O2O DO�/�/�/�/�?�O�/ �O�O�O
__�?@_R_ d_v_�_�O-_�_�_�_ �_oUOgOyO�O�_ro �O�o�o�o�o�o�_ &8Jmo�o�� ���o)o;oMoO !��oX�j�|�����o ď֏����/���B��T�f�x���^�ST_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
�FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@oG %j%@�_MOV�u����MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�5�
��5���۵MO~q_�DCd~�1PL_N�AME !<u�� �!Defa�ult Pers�onality �(from FD�) �4RR2k! �1j)TEX)TsH��!�AX d�? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO@^OpO�O�O�Ox2-? �O�O�O__0_B_T_f_x_�b<�O�_�_�_ �_�_�_o o2oDoVotho&xRj" 1o�)�&0\�b, ��9��b�a @D��  �a?��c�a?x�`�a�aA'�6�e�w;�	l�b	� �xJp��`�`	p� �< ��(p� �.r� K��K ��K=�*�J���J���JV��kq`�q�P�x�|� @j�@T;f�r��f�q�acrs��I�� ��p���p�r�ph}�3���´  ��>���ph�`z��w꜖"�Jm�q� H�N��ac��$��dw��  ��  P� Q� �>� |  а�m��Əi}	'� �� �I� ��  ����:��È�È=����(��#�a	���I�  �n @@H�i~�ab�Ӌ�b�$�w���"N0��  �'Ж�q�p@2��@����r�q5��C�pC0C�@� C����`
��A1q �  @B�V~JX�
nwB0h�A���p�ӊ�p�`���aDz���֏���Я	��pv�( �� -��I��-��=��A�a�we_q��`�p �?�ff� ��m��� ����Ƽ�!@ݿ:�>1�  P�apv(�`ţ� �=�qs�t��?���`x�`�� <
6b<�߈;܍�<��ê<� <�#&P�ό�AO��c�1��ƍ�?fff?�O�?&��qt@�.��J<?�`��wi4����dly�e ߾g;ߪ�t��p�[� ��߸ߣ����� ��0��6�wh�F0%� r�!��߷�1ى���~�E�� E�O�?G+� F�!��� /���?�e�P���t���lyBL�cB��Enw 4�������+��R�� s����������h�Ô�>��I�mXj���A�y�we�C�������A�#/*/c/N/wi������v/C�`� C!Hs/`
=$�p�<!�!���ܼ�'�3A��A�AR1AO��^?�$�?����±
=���>����3�?W
=�#�]�;�e�׬a@�����{����<��>(�B��u��=B0�������	�R��zH�F�G����G��H��U`E���C��+��}I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0w/O*OONO9O rO]O�O�O�O�O�O�O �O_�O8_#_\_G_�_ �_}_�_�_�_�_�_�_ "oooXoCo|ogo�o �o�o�o�o�o�o	 B-fQ�u�� �����,��P� b�M���q�����Ώ�� �ݏ�(��L�7�p� [������ʟ���ٟ ���6�!�Z�E�W���:#1( ��9�K����ĥ ���x��Ư!3�8��<�!4Mgs���,�IB+8�J��a?���{�d�d������ȿ���ڼ%P8�P�=:GϚ�`S�6�h�z���R��������������  %�� ��h�Vߌ�z� ��&�g�/9�$�������7����A�S�e�w�  ��������������2 wF�$�&Gb���������!C����@���8�����F�� DzN��� F�P D�������)#B�'9�K]o#?��ͫ@@v
4$8��8��8�.
 v���!3 EWi{�����:� ��ۨ��1��$MSKCFMAP  ��� ����(.�ONREoL  �!�9��EXCFEN�BE'
#7%^!FN�Ce/W$JOGOV�LIME'dO S"d��KEYE'�%��RUN�,�%��SFSPDTY�0g&P%9#SIGN|E/W$T1MOT�/�T!�_CE_G�RP 1p��#\x��?p��?�? �?�?�?O�?OBO�? fOO[O�OSO�O�O�O �O�O_,_�OP__I_ �_=_�_�_�_�_�_o�o�_:o�TCO�M_CFG 1qB	-�vo�o�o
Va__ARC_b"��p)UAP_CPL��ot$NOCHEC�K ?	+ �x�%7I[ m���������!�.+NO_WAIT_L 7%S2�NT^ar	+��s�_ERR_12s	)9�� ,ȍޏ���x���&��dT�_MO��t��, �/�*oq�9�PA�RAM��u	+���a�ß'g{�� �=?�345678901��,��K� ]�9�i�������ɯۯ��&g�����C���cUM_RSPA�CE/�|����$?ODRDSP�c#6�p(OFFSET_�CART�o��DI�Sƿ��PEN_FILE尨!�ai��`�OPTION_I�O�/��PWORK� ve7s#  ��V�ؤ��p�4�p�	 ���p��<����RG_DSBOL  ��P#���ϸ�RIENTT5OD ?�C�� !�l�UT_SIM�_D$�"���V~��LCT w}��h�iĜa[�1�_PEsXE�j�RATv�Ш&p%� ��2^3j)TEX)TH�)�X d3����� ��%�7�I�[�m�� �������������!�3�E���2��u��� ������������c�<d�ASew� ��������썒^0OUa0o(ҿ�(����>u2, ���O ~H @D�  [?�aG?��cc��D][�Z�;��	ls��xoJ���������< ���� ��2�H�(��H3k7H�SM5G�22G���Gp
͜��'f�/-,2�C%R�>�D!�M#{|Z/��3�����4y H "�c/u/��/0B_���{�jc��t�!�/ �/�"t32�����/6  ���P%�Q%��%�|�T��S62�q?'e	'�� � �2I�� �  �=�+==��ͳ?�;�	�h	�0�I  ?�n @�2�.��Ov;��ٟ?&g9N�]O  ''�uDt@!� C�C�@F#�H!�/�O�O sb
����@�@�H�@�e`0B�QA�0Yv: �13Uwz$oV_�/z_e_�_�_�	��( �� -�2�1�1ta��Ua�c���:A-����.  �?�ff ���[o"o�_U�`oDXÜQ8���o�j>�1'  Po�V(���e�F0�f�Y���L�?�����xb�P<�
6b<߈;�܍�<�ê<� <�&�,/aA�;r�@Ov0P�?fff?�0?&�ip�T@�.{r�?J<?�`�u#	 �Bdqt�Yc�a� Mw�Bo��7�"�[� F��j�������ُ� ���3����,����(�E�� E�~�3G+� F��a ��ҟ�����,��PP�;���B�pAZ� >��B��6�<OίD��� P��t�=���a�s���<��6j�h��7o��>�S��O��0���Fϑ�A�a�_���C3Ϙ�/�%?��?���������#	�Ę��P �N||CH���Ŀ�������@I�_�'�3�A�A�AR1�AO�^?�$��?��� �±
�=ç>�����3�W
=�#�\ U��e���B��@���{����<����(�B��u��=B�0�������	�b�H�F�G����G��H��U`E���C��+��I#��I��HD��F��E��R�C�j=[�
�I��@H�!�H�( E<YD0߻������ ��� �9�$�]�H�Z� ��~������������� #5 YD}h� ������
 C.gR���� ���	/�-//*/ c/N/�/r/�/�/�/�/ �/?�/)??M?8?q? \?�?�?�?�?�?�?�? O�?7O"O[OmOXO�O |O�O�O�O�O�O�O�Ot3_Q(�������b��gUU���W_i_2�3�8�x�_�_2�4Mgs�_��_�RIB+�_�_�a���{�m iGo5okoYo�o}l��%P'rP�nܡݯ�o�=_�o�_�[R�?Q�u���  �p���o��/� �S��z
uүܠ�������ڱ�������8����  /�M��w�e��������l2 �F�$��Gb���t��a�`�p�S�C�y�@p�5�G�Y�۠�F� Dz��� F�P D�!�]����پ��ʯ�ܯ� ��~�?��W�@@�?�K��K���K���
 �|�������Ŀ ֿ�����0�B�TϸfϽ�V� ���{���1��$PAR�AM_MENU �?3���  DE�FPULSEr��	WAITTMO{UT��RCV��� SHELL�_WRK.$CU�R_STYL���	�OPT��P�TB4�.�C�R_DECSN���e�� ߑߣ���������� �!�3�\�W�i�{�����USE_PRO/G %��%����.��CCR���e�����_HOST �!��!��:���T �`�V��/�X��>��_TIME��^���  ��GDE�BUG\�˴�GI�NP_FLMSKĻ���Tfp����PG�A  ����)CyH����TYPE��������� �� -?hc u������� //@/;/M/_/�/�/ �/�/�/�/�/�/??�%?7?`?��WORD� ?	=	R}Sfu	PNSU�Ԝ2JOK�DR�TEy�]TRACECTL 1x3���� �`/ &�`�`�>��6DT Qy3��%@�0D � ޱc�a0:@V�@BR�2ODO VOhO�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟���`� �2�D�V�.I v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� j����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o��o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ����������*��$PGT�RACELEN � )�  ���(��>�_�UP z��e�m�u�Y�n��>�_CFG {Fm�W�(�~����PКӂ�DEFSP/D |��'�P���>�IN��TR�L }��(�8�����PE_CON�FI��~m���mњ��ղ�L�ID����=�G�RP 1��W���)�A ����&ff(�A+33�D�� D]� ?CÀ A@1����(�d�Ԭ��0�0�?� 	 1��8�֚��� ´�����B�9����O��9�s�(�>�T?��
5�������� �=��=#�
 ����P;t_�������� G Dz (�
 H�X~i��� ���/�/D///�h/S/�/��
V7�.10beta1���  A��E�"ӻ�A �(�� ?!G��!>����"����!{���!BQ��!�A\� �!���!2p
����Ț/8?J?\?�n?};� ���/� �/�?}/�?�?OO:O %O7OpO[O�OO�O�O �O�O�O_�O6_!_Z_ E_~_i_�_�_�_�_�_ �_'o2o�_VoAoSo �owo�o�o�o�o�o�o .R=v1�/�#F@ �y�}� �{m��y=��1�'� O�a��?�?�?������ ߏʏ��'��K�6� H���l�����ɟ��� ؟�#��G�2�k�V� ��z��������o� �ίC�.�g�R�d��� �������п	���-� ?�*�cώ���Ϯ� �����B�;�f� x�������DϹ��߶� �������7�"�[�F� X��|��������� ��!�3��W�B�{�f� �������� ����� /S>wbt� �����= OzόϾψ����� �� /.�'/R�d�v� �߁/0�/�/�/�/�/ �/�/#??G?2?k?V? h?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O���O�O�O__ ?_*_c_N_�_r_�_�_ �_�_�_o�_)oTf x�to���/�o />/P/b/t/m o�|����� ��3��W�B�{�f� x�����Տ������ �A�S�>�w�b����O ��џ������+�� O�:�s�^�������ͯ ���ܯ�@oRodo�o `��o�o�o��ƿ�o� ��*<N�Y��}� hϡό��ϰ������� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�c�N�ﲟ��� l��������;�&� _�J���n��������� ��,�>�P�:L�� ���������� (�:�3��0iT� x�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?a?s?��?�?X?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O *\&_8_r����_�_��$PLI�D_KNOW_M�  ��� Q�TSV ���P��?o"o4o�OXo�CoUo�o R�SM_?GRP 1��Z'U0{`�@�`uf
�e�`
�5� �gpk 'Pe] o�������X���SMR�c��m1T�EyQ}? yR�� ��������폯���ӏ �G�!��-������� ����韫���ϟ�C� ��)������������寧���QST�a1W 1��)���P;0� A 4��E 2�D�V�h�������߿ ¿Կ���9��.�o� R�d�vψ��ϬϾ�����2�0� Q�	<3��3�/�A�S߂�4l�~ߐߢ��5 ���������6
��.�@��7Y�k�}���8��������M_AD  )���PARNUM  !�}o+��WSCHE� S�
��pf���S��UPDf��x��_CM�P_�`H�� �'��UER_CHK-���ZE*<�RSr��_�Q_MO�G���_�X�_R/ES_G��!��� D�>1bU� y�����/�	/����+/� k�H/g/l/��Ї/�/ �/�	��/�/�/�X� ?$?)?���D?c?h?�����?�?�?�V �1��U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_�INRr�J�b�Ud�2FMASS?O Z�SGMN>OqCMON�_QUEUE a��U�V P~P X�N$ UhN�FV�@�END�A��IEX1E�O�E��BE�@�O>�COPTIO�G���@PROGRAM7 %�J%�@�?����BTASK_I�G�6^OCFG ኤOz��_�PDATuA�c��[@Ц2=�DoVohozo�j2o �o�o�o�o�o)x;M jINFO[��m��D��� �����1�C�U� g�y���������ӏ����	�dwpt�l �)�QE DIT ��_i��^WERF�LX	C�RGADoJ �tZA���¿�?נʕFA��IOORITY�GW���MPDSPNQ�����U�GD��OTO�E@1�X� (/!AF:@E� c�~Ч!tcpn�>��!ud����!icm���?<��XY_�Q�X�=��Q)� *�1�5��P��]�@�L� ��p��������ʿ� �+�=�$�a�Hυϗ�=*��PORT)QH���P�E��_C?ARTREPPX�>�SKSTA�H�
�SSAV�@�tZ	�2500H86A3���_x�
�'��X�@�swPtS��x�ߧ���URGE�@�B��x	WF��DO�F"[W\��������WRUP_DEL�AY �X���RO_HOTqX	B%��c���R_NORM�ALq^R��v�SE�MI�����9�QS�KIP'��tUr�x 	7�1�1�� X�j�|�?�tU������ ��������$J \n4����� ���4FX |j������ �/0/B//R/x/f/�/�/�/tU�$RCgVTM$��D�� �DCR'������!?��LB�'��CE�>�x��=��8.�(gC����e���ߠ�������:�o?�� �<
6b<߈�;܍�>u.��?!<�& �?h?�?�?�@>��?O  O2ODOVOhOzO�O�O �O�O�O�?�O�O__ @_+_=_v_Y_�_�_�? �_�_�_oo*o<oNo `oro�o�o�o�_�o�o �o�o�o8J-n ��_������ �"�4�F�X�j�U�� ����ď���ӏ�� �B�T��x������� ��ҟ�����,�>� )�b�M����������� �ïկ�Y�:�L�^� p���������ʿܿ�  ����6�!�Z�E�~� ��{ϴϗ�����-��  �2�D�V�h�zߌߞ� ����������
���.� �R�=�v��k��� �������*�<�N� `�r������������ ����&J\? �������� "4FXj|���!GN_ATC �1�	; �AT&FV0E0��ATDP/6/9/2/9��ATA�,�AT%G1%B�960�++U+�,�H/,�!�IO_TYPE � �%�#t�R�EFPOS1 1}�V+ x�u/�n�/j�/
=�/ �/�/Q?<?u??�?4?�?X?�?�?�+2 1�V+�/�?�?\O�?x�O�?�!3 1�O�*O<OvO�O�O_�OS4 1��O�O�O_��_t_�_+_S5 1�B_T_f_�_o	oBo>�_S6 1��_�_��_5o�o�o�oUoS7 1�lo~o�o�oH�3l�oS8 1� %_����SMASK 1��V/  
?�M��XNOS/�r�����~�!MOTE  n���$��_CFG ᢫��q���"PL_�RANG�����POWER ������SM_DRYPRG %o��%�P��TART� ��^�UME_PRO-�?����$�_EXEC_EN�B  ���GS�PD��Րݘ��T3DB��
�RM�
��MT_'�T�����OBOT_NA_ME o�����OB_ORD_�NUM ?��b!H863�  �կ����PC_TIMoEOUT�� x�oS232Ă1��� LTEA�CH PENDA1N��w��-���Mainte�nance Co#ns���s�"���?KCL/Cm��
�
���t�ҿ ?No Use-��8Ϝ�0�NPO�򁮋���.�C7H_L������q�	��s�MAVA#IL�����糅���SPACE1 2��, j�߂�D��s�߂� �{S�?8�?�k�v� k�Z߬��ߤ��ߚ�  �2�D���hߊ�|�� `����������  �2�D��h��|����`���������y���2����0�B���f� ����{���3);M_ ������/� /44FXj| */���/�/�/?(??=?5Q/c/u/�/ �/G?�/�/�?O�?$OEO,OZO6n?�?�? �?�?dO�?�?_,_�O A_b_I_w_7�O�O �O�O�O�_�O_(oIo@o^oofo�o8�_ �_�_�_�_�oo6oE�f){���Gw �o� �:��
M� ��� *�<�N�`�r������� w���o�収���d.��%�S�e�w��� ��������Ǐَ��� Θ8�+�=�k�}����� ��ůׯ͟����%� '�X�K�]��������� ӿ������#�E��W� `� @ �������x�����\�e����������� R�d߂�8�j߬߾߈� �ߤ����������0� r���X�������@������8����
�����_MODE � �{��S �"�{|�2�0��ψ��3�	S|)CWORK_AD���R�+R  ��{�`� �� _?INTVAL���d����R_OPTI[ON� ��H �VAT_GRP �2��up#(N�k| ��_����� /0/B/��h�u/T�  }/�/�/�/�/�/�/? !?�/E?W?i?{?�?�? 5?�?�?�?�?�?O/O AOOeOwO�O�O�O�O UO�O�O__�O=_O_ a_s_5_�_�_�_�_�_ �_�_o'o9o�_Iooo �o�oUo�o�o�o�o�o �o5GYk-� ��u����� 1�C��g�y���M��� ��ӏ叧�	��-�?� Q�c������������ ���ǟ�;�M�_�����$SCAN_GTIM��_%}��R �(�#(�(�<04+d d 
!AD�ʣ��u�/X�����U���25���@�d5�P�g��]	�������p��dd�x�  P����� �� � 8� ҿ�!���D��$�M�_�qσ� �ϧϹ��������ƿv��F�X�x�/� ;�ob���pm��t�_DiQ̡  � l�|�̡ĥ �������!�3�E�W� i�{���������� ����/�A�S�e�] �Ӈ������������� );M_q� ������ r���j�Tfx�� �����//,/ >/P/b/t/�/�/�/�/8�/�%�/  0��6 ��!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O* �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo�O �OJ�o�o�o�o�o�o �o 2DVhz �������
�7?  ;�>�P�b� t���������Ǐُ� ���!�3�E�W�i�{�p������ß �ş 3�ܟ��&�8�J�\�@n�������������ɯ����,� ��+�	123�45678�� +	� =5���f� x����������� ��
��.�@�R�d�v� �Ϛ�៾�������� �*�<�N�`�r߄߳� �ߺ���������&� 8�J�\�n�ߒ��� ���������"�4�F� u�j�|����������� ����0_�Tf x������� I>Pbt� ������!/ (/:/L/^/p/�/�/�/�/�/�/�2�/?��#/9?K?]?�iC�z  Bp˚  � ��h2��*��$SCR_GRP� 1�(�U8(�\xd��@ � ��'�	 �3�1�2 �4(1*�&�I3�F1O�OXO}m��D!�@�0ʛ)���HUK��LM-10i�A 890?�90�;��F;�M61CA D�:�CP��1
\&V�1	�6F��CW�9)A7Y	(R�_�_Ф_�_�_�\�� �0i^�oOUO>oPo #G�/���o'o�o�o\�o�oB�0��rtAA�0*  !@�Bu&Xw?��ju��bH0{UzAF@ F�`�r��o �����+��O� :�s��mBqrr����������B�͏b���� 7�"�[�F�X���|��� ��ٟğ���N���AO�0�B�CU
L���E�<jqBq=��Ҕ�$Gs@�@pϯ B����G�I
E�0EL�_DEFAULT�  �T���E��MIP�OWERFL  �
E*��7�WFD�O� *��1ER�VENT 1����`(�� L!�DUM_EIP���>��j!AF�_INE�¿C�!'FT������9!o:� ��a��!RPC_MAINb�DȺPϭ�t�'VIS}�Cɻ����o!TP��PU���d��E�!
PM�ON_PROXYF߮�e4ߑ��_ߧ��f����!RDMO_SRV�߫�g�ߎ)�!R�Iﰴh,�u�!
v�M�ߨ��id���!RLSgYNC��>�8��>�!ROS��4��4��Y�(�}���J� \������������� 7��["4F�j |����!�E�io�ICE_K�L ?%� (�%SVCPRG�1n>���3��3����4//�5�./3/�6V/[/�7@~/�/��D�/�9�/�+�@��/��#? ��K?��s?� / �?�H/�?�p/�?� �/O��/;O��/cO �?�O�9?�O�a? �O��?_��?+_� �?S_�O{_�)O�_ �QO�_�yO�_��O s����>o�o}1 �o�o�o�o�o�o�o ;M8q\�� �������7� "�[�F��j������� ُď���!��E�0� W�{�f�����ß��� ҟ���A�,�e�P� ��t��������ί��y_DEV ~��MC:��@`!�OUT���2��REC� 1�`e�j�= �� 	 ������˿���ڿ��
 �`e���6�N�<� r�`ϖτϦ��Ϯ��� ����&��J�8�n߀� bߤߒ��߶������� "��2�X�F�|�j�� ������������� .�T�B�x�Z�l����� ��������,P >`bt���� ��(L:\ �d����� / �$/6//Z/H/~/l/ �/�/�/�/.��/?�/ 2? ?V?D?f?�?n?�? �?�?�?�?
O�?.O@O "OdORO�OvO�O�O�O �O�O�O__<_*_`_ N_�_�_x_�_�_�_�_ �_oo8oo,ono\o �o�o�o�o�o�o�o �o "4jX�� �������� B�$�f�T�v������� �����؏��>�,��b�P�r���p�V 1��}� P
�ܟ� y���TYPE\���HELL_CFOG �.��͟�  	�����RSR������ӯ�� �����?�*�<�u� `�����������ο�  �%@�3�E��Q�\���1M�o�p��d���2��d]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&��1�OW_REG�_UI��8�IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he�#�� ������������) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������o���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( ��}(copy f�rs:*.dt �virt:\te�mp\=>ins�piron:5072 O^p���o�}xyzrate 61GHZ����3.or�derfil.d�a:mpback@Fas��� *.mdb6 *C�
Y��/�	0.@C2636 �p/�/ �/�-G/Y#W/�/�/?�
� �/�/�/ n?�?�?��	Z2H?Z? �?�?O"4/�U'aO sO�O�O�EOT(YO�O��O_�9.x�$:\ �O8PO-�On_�_�_�5/.Ua6_H_�0^_�_ oo&O8O�O�Omoo �o�O�O�OZo�o�o "_4_�_X_i{��_ �_C�_���o0o BoToe�w����o�oI� �o�����,�P a�s������;��`� ���(>��˟ݟn�������?�	4940 H�Z�����"�4� ����a�s�������E� ��Y�����!�3�F� £ݿnπϒϥ�6�H� Š^�����&�8������m�ߑߤ��
8124ǯY������!� 33������n�����:488G�Y����� �!�3�����a�s��� ����E���Y����� !�3�F�����n�� ��6H��^� &�8�����m��� ����Z��/"4 �Xi/{/�/��C/ ��/�/?0BT e?w?�?��I?��?��?OO�$SNP�X_ASG 1�����9A�� P 0 �'%R[1]�@1.1O 9?�$3%dO�OsO�O�O�O �O�O�O __D_'_9_ z_]_�_�_�_�_�_�_ 
o�_o@o#odoGoYo �o}o�o�o�o�o�o�o *4`C�gy �������	� J�-�T���c������� ڏ�����4��)� j�M�t�����ğ���� ��ݟ�0��T�7�I� ��m��������ǯٯ ���$�P�3�t�W�i� �������ÿ���� :��D�p�Sϔ�wω� �ϭ��� ���$��� Z�=�dߐ�sߴߗߩ� ������ ��D�'�9� z�]��������� 
����@�#�d�G�Y� ��}������������� *4`C�gy ������	 J-T�c��� ���/�4//)/ j/M/t/�/�/�/�/�/��/�/?0?4,DPA�RAM �9E}CA �	��:�P�4�0$HOF�T_KB_CFG�  q3?E�4PI�N_SIM  9K�6�?�?�?�0,@�RVQSTP_DSB�>�21On8J0�SR ��;� G& =O{Oq0�6�TOP_ON_E_RR  q4�9~�APTN �5��@A�BRING_PRM�O� J0VDT_G�RP 1�Y9�@  	�7n8_(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2Dkhz �������
� 1�.�@�R�d�v����� ����Џ�����*� <�N�`�r��������� ̟ޟ���&�8�J� \�����������ȯگ ����"�I�F�X�j� |�������Ŀֿ�� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�tߛߘߪ� ����������(�:� a�^�p������� ���� �'�$�6�H�Z� l�~���������������3VPRG_CO7UNT�6��A�5NENB�OM=��4J_UPD 1}��;8  
 q2������  )$6Hql~� ����/�/ / I/D/V/h/�/�/�/�/ �/�/�/�/!??.?@? i?d?v?�?�?�?�?�? �?�?OOAO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_��_�_YSDEBSUG" � �Pdk	��PSP_PASS�"B?�[LOG� ��mr�P�X�_  �g~�Q
MC:\d<�_b_MPCm�H�o�o�Qa�o �~vfSAV �m�:dUb�U\gS�V�\TEM_TI�ME 1�� �(�P4�T3�o	T1SVGUNS} �#'k�spAS�K_OPTION�" �gospBC?CFG ��|c �b��z`� ���4��X�C�|�g� ����ď֏������ 	�B�-�f�Q�c����� �����ϟ��,�>�)�b��YR���S��� ƯA������ ��D� �nd��t9�l������� ��ڿȿ�����"� X�F�|�jϠώ��ϲ� ��������B�0�f� T�v�xߊ��ߦؑ��� ����(��L�:�\� ��p���������� � �6�$�F�H�Z��� ~������������� 2 VDzh�� �������4 Fdv���� ��//*/�N/</ r/`/�/�/�/�/�/�/ �/??8?&?\?J?l? �?�?�?�?�?�?�?�? OO"OXOFO|O2�O �O�O�O�OfO_�O_ B_0_f_x_�_X_�_�_ �_�_�_�_oooPo >otobo�o�o�o�o�o �o�o:(^L np�����O� �$�6�H��l�Z�|� ����Ə؏ꏸ���� 2� �V�D�f�h�z��� ��ԟ����
�,� R�@�v�d��������� ίЯ���<��T� f�������&�̿��ܿ ��&�8�J��n�\� �π϶Ϥ�������� ��4�"�X�F�|�jߌ� �ߠ����������� .�0�B�x�f��R��� ���������,��<� b�P�������x����� ����&(:p ^�������  6$ZH~l ��������/ &/D/V/h/��/z/�/��/�/�/�&0�$T�BCSG_GRP� 2��%��  �1 
? ?�  /?A? +?e?O?�?s?�?�?�?��?�;23�<d�, �$A?1	� HC���6>�@E�5CL  �B�'2^OjH4Jݸ�B\)LFY g A�jO�MB��?F�IBl�O�O�@�JG|_�@�  D	�15_ __$YC-P{_F_$`_j\��_�]@0�> �X�Uo�_�_6oSoo�0o~o�o�k�h�0	V3.00'2�	m61c�c	�*�`�d2�o�e>əJC0(�a�i �,p�m-  �0�����omvu1JC�FG ��%� 1 #0vz��r8Br�|�|��� �z� �%��I�4�m� X���|��������֏ ���3��W�B�g��� x�����՟������ ��S�>�w�b����� '2A ��ʯܯ����� �E�0�i�T���x��� ÿտ翢����/�� ?�e�1�/���/�Ϝ� ���������,��P� >�`߆�tߪߘ��߼� �������L�:�p� ^����������� � �6�H�>/`�r�� ��������������  0Vhz8�� ����
.� R@vd���� ���//</*/L/ r/`/�/�/�/�/�/�/ �/�/?8?&?\?J?�? n?�?�?�?�?���?O O�?FO4OVOXOjO�O �O�O�O�O�O__�O B_0_f_T_v_�_�_�_ z_�_�_�_oo>o,o boPoroto�o�o�o�o �o�o(8^L �p������ �$��H�6�l�~�(O ����f�d��؏��� 2� �B�D�V������� n����ԟ
���.�@� R�d����v������� �Я���*��N�<� ^�`�r�����̿��� ޿��$�J�8�n�\� �π϶Ϥ�������� ��(�:�L���|�jߌ� �ߠ����������0� B�T��x�f���� ���������,��P� >�t�b����������� ����:(JL ^������  �6$ZH~l ��^���dߚ / /D/2/h/V/x/�/�/ �/�/�/�/�/?
?@? .?d?v?�?�?T?�?�? �?�?�?OO<O*O`O NO�OrO�O�O�O�O�O _�O&__6_8_J_�_ n_�_�_�_�_�_�_�_ "ooFo��po�o,o Zo�o�o�o�o�o0 Tfx�H�� �����,�>�� b�P���t��������� Ώ��(��L�:�p� ^�������ʟ���ܟ � �"�$�6�l�Z��� ~�����دꯔo�� &�ЯV�D�z�h����� ��Կ¿��
��.���R�@�v�dϚτ�  9���� ��������$TBJOP_GRP 2ǌ���  �?������������x�JBЌ��9� �< �X�=��� @���	 �C�� t�b  C���я>��͘Րդ�>�̚йѳ33=�CLj�fff}?��?�ffBGР�ь�����t�ц�>w�(�\)�����E噙�;���hCYj��  @�h��B�  A�����f��C�  �Dhъ�1��O��4�N����
:_���Bl^��j��i�l�l����Aəg�A�"��D���֊=qH���н�p�h�Q�;��A�j�ٙ�@L��D	2�����x��$�6�>B�\���T���Q�tsx�@�33@���C����y�1����>�#�Dh�����������<{�h�@ i� ��t��	 ���K&�j �n|���p�@/�/:/k/�ԇ����!��	V3.�00J�m61cI�*� IԿ��/�'� Eo�E���E��E��F��F�!�F8��F�T�Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G�,I�!CH`��C�dTDU�?�D��D��D�E(!/E\��E��E�h��E�ME��s�F`F+'\�FD��F`=�F}'�F���F�[
F����F��M;��;Q��T,8�4` *(�ϴ?�2���3\��X/O��ESTPARS  ��	����HR@ABLE K1����0��
H��7 8��9
G
HP
H����
G	
H

HQ
HYE��
H
Hu
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_$�^:BS _� �JGo Yoko}o�o�o�o�o�o �o�o1CUg y����`#oRL�y �_�_�_�_�O�O�O�O��OX:B�rNUM [ ���P���� V@P:B_CFG ˭�Z�h��@��IMEBF_�TT%AU��2@�V�ERS�q��R� 1���
 ($�/����b� ���� J�\���j�|���ǟ�� ȟ֟�����0�B��T���x�������2�_ԧ��@�
��MI__CHAN�� �} ��DBGLV����������ETHERAD ?��O�������h������ROUT��!��!������SNMASKD��U�255.���#������OOLOFS�_DI%@�u.�O�RQCTRL �����}ϛ3rϧϹ� ��������%�7�I߀[�:���h�z߯�APE_DETAI"��G�PON_SVO�FF=���P_MOON �֍�2���STRTCHK ��^�����VT?COMPAT��O������FPROG �%^�%GET�DAT����9�P�LAY&H��_IN�ST_Mް �������US�q��L�CK���QUIC�KME�=���SC�REZ�G�tps� ���u�z�����_��@@n�.�S�R_GRP 1о^� �O� ���
��+O=sa�쀚�
m�� ����L/C 1gU�y��� ��	/�-//Q/?/�a/�/	1234�567�0�/�/@X�t�1���
 �}�ipnl/� g?en.htm�?� ?2?D?V?`P�anel setupZ<}P�?�?�?�?�?�? �??,O >OPObOtO�O�?�O!O �O�O�O__(_�O�O ^_p_�_�_�_�_/_]_ S_ oo$o6oHoZo�_ ~o�_�o�o�o�o�o�o so�o2DVhz� 1'���
�� .��R��v��������ЏG���UALR�M��G ?9� �1�#�5�f�Y��� }�������џן����,��P��SEV � ����E?CFG ������A��   BȽ�
 Q���^� ���	��-�?�Q�c�@u�������������C �����I��?���(%D�6� � $�]�Hρ�lϥϐ��� ��������#��G����� �߿U�I_�Y�HIST 1վ�  (��� ��,/SOF�TPART/GE�NLINK?cu�rrent=editpage,��,1����,�;��� ����menu��962�߆���0��K�]�o�36u�
� �.�@���W�i�{��� ������R����� /A��ew��� �N��+= O�s��������f��f//'/ 9/K/]/`�/�/�/�/ �/�/j/�/?#?5?G? Y?�/�/�?�?�?�?�? �?x?OO1OCOUOgO �?�O�O�O�O�O�OtO �O_-_?_Q_c_u__ �_�_�_�_�_�_�� )o;oMo_oqo�o�_�o �o�o�o�o�o%7 I[m� �� �����3�E�W� i�{������ÏՏ� ������A�S�e�w� ����*���џ���� �ooO�a�s����� ����ͯ߯���'� ��K�]�o��������� F�ۿ����#�5�Ŀ Y�k�}Ϗϡϳ�B��� ������1�C���g� yߋߝ߯���P����� 	��-�?�*�<�u�� ������������ )�;�M���������� ������l�%7 I[������ �hz!3EW i������� v////A/S/e/P����$UI_PA�NEDATA 1������!�  	�}�w/�/�/�/�/?? )?>?��/i?{?�? �?�?�?*?�?�?OO OAO(OeOLO�O�O�O��O�O�O�O�O_&Y� b�>RQ?V_h_ z_�_�_�__�_G?�_ 
oo.o@oRodo�_�o oo�o�o�o�o�o�o *<#`G��}�-\�v�#�_�� !�3�E�W��{��_�� ��ÏՏ���`��/� �S�:�w���p����� џ������+��O� a���������ͯ߯ �D����9�K�]�o� �������ɿ���Կ �#�
�G�.�k�}�d� �ψ����Ͼ���n��� 1�C�U�g�yߋ��ϯ� ��4�����	��-�?� ��c�J������ ���������;�M�4� q�X����������� %7��[�� �����@� �3WiP�t �����/�// A/����w/�/�/�/�/ �/$/�/h?+?=?O? a?s?�?�/�?�?�?�? �?O�?'OOKO]ODO �OhO�O�O�O�ON/`/ _#_5_G_Y_k_�O�_ �_?�_�_�_�_oo �_Co*ogoyo`o�o�o �o�o�o�o�o-`Q8u�O�O}��@������)� >��U-�j�|������� ď+��Ϗ���B� )�f�M���������������ݟ�&�S�K��$UI_PANELINK 1�U�  ��  ��}1�234567890s���������ͯդ �Rq����!�3�E�W� �{�������ÿտm��m�&����Qo�  �0�B�T�f�x�� v�&ϲ���������� ��0�B�T�f�xߊ�"� �����������߲� >�P�b�t���0�� ����������$�L� ^�p�����,�>�����`�� $�0,&� [gI�m��� ����>P3 t�i��Ϻ�  -n��'/9/K/]/o/ �/t�/�/�/�/�/�/ ?�/)?;?M?_?q?�? �UQ�=�2"��?�? �?OO%O7O��OOaO sO�O�O�O�OJO�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5oGo�_ko}o�o�o �o�oTo�o�o1 C�ogy���� �B�	��-��Q� c�F�����|������ �֏�)��M���= �?��?/ȟڟ��� �"�?F�X�j�|��� ��/�į֯����� 0��?�?�?x������� ��ҿY����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z���� -���������
��. RdG��}� ���c���<�� `r������� �//&/8/J/�n/ �/�/�/�/�/7�I�[� 	�"?4?F?X?j?|?� �?�?�?�?�?�?�?O 0OBOTOfOxO�OO�O �O�O�O�O_�O,_>_ P_b_t_�__�_�_�_ �_�_oo�_:oLo^o po�o�o#o�o�o�o�o  ��6H�l~ a������� �2��V�h�K����� ��1�U
��.� @�R�d�W/�������� П������*�<�N� `�r��/�/?��̯ޯ ���&���J�\�n� ������3�ȿڿ��� �"ϱ�F�X�j�|ώ� �ϲ�A��������� 0߿�T�f�xߊߜ߮� =���������,�>� ��b�t�����+ ������:�L�/� p���e�����������  ��6���ۏ���$UI_QU�ICKMEN  }���}���RESTOR�E 1٩�  �
�8m3\n ���G���� /�4/F/X/j/|/' �/�/�//�/�/?? 0?�/T?f?x?�?�?�? Q?�?�?�?OO�/'O 9OKO�?�O�O�O�O�O qO�O__(_:_�O^_ p_�_�_�_QO[_�_�_ I_�_$o6oHoZoloo �o�o�o�o�o{o�o  2D�_Qcu�o �������.� @�R�d�v��������xЏ⏜SCRE� �?�u1�sc� u2�3��4�5�6�7��8��USER�����T���ksT'���4��5��6���7��8��� NDO_CFG ڱ�  �  � PD�ATE h���None�S�EUFRAME � ϖ��RTOL_ABRT�����ENB(��G�RP 1��	�?Cz  A�~�|��%|�������į֦��X�� UH�X�7�?MSK  K�S��7�N�%uT�%������VISCA�ND_MAXI��I�3���FAILO_IMGI�z �% �#S���IMREG�NUMI�
���S�IZI�� �ϔ�,�ONTMOU4'�K�Ε�&�����a��a���s�FR:\��� � M�C:\(�\LOGnh�B@Ԕ !{��Ϡ�����z �MCV����7UD1 �EX	��z ��PO64_t�Q��n6��PO!�LI�Oڞ�re�V�N�f@`��I�� =	_�SZ�Vmޘ��`�WA�Imߠ�STAT �k�% @��4�F��T�$#�x �2D�WP  ��P� G��=��������_JMP�ERR 1ޱ
�  �p2345678901��� 	�:�-�?�]�c����� ������������$�MLOW�ޘ�����g_TI/�˘'���MPHASE  �k�ԓ� ��SH�IFT%�1 Ǚ��<z��_� ���F/| Se������ �0///?/x/O/a/��/�/�/�/�/�����k�	VSFT1�\�	V��M+3 S�5�Ք p���ſA�  B8[0�[0�Πpg3a1Y2�_3Y�7ME��K�͗q	6e���&%���M���b��	���$��TDINEND3�4��4OH�+�G�1�OS2OIV I�{��]LRELEv�I��4.�@��1_AC�TIV�IT��B��A �m��/_��B�RDBГOZ�YBO�X �ǝf_\���b�2�TI�190.0.�P8�3p\�V254tp^�Ԓ	 �S��_�[b��r�obot84q_   p�9o\�pc�PZoMh�]�Hm�_Jk@1�o�ZA+BCd��k�,���P \�Xo}�o0); M�q����� ���>��aZ�b��_V