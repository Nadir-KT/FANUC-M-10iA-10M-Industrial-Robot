��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �� �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ڏ1�	 H PC�UREQ1 � $SOFT; �T_ID�TOT�AL_EQ� $� � NO�PS_�SPI_INDE���$�X�SC�REEN_NAM�E �SI�GN��� P�K_FIL	$�THKYMPAN�E�  	$D�UMMY12 �� u3|4|&��ARG_STR�1 � $T�ITP$I��1�{������5�6�7�8
�9�0��z�P����1�1��1 '1
'2"GS�BN_CFG1 � 8 $CN?V_JNT_* |�$DATA_C�MNT�!$FL�AGS�*CHE�CK�!�AT_C�ELLSETUP�  P $HOME_IO,�G�%�#MACR=O�"REPR�(-�DRUN� D|�3SM5H UTO�BACKU0� $ENAB���!EVIC�T]I � D� �DX!2ST� ?0B��#$INTERV�AL!2DISP_�UNIT!20_D�On6ERR�9FR�_F!2IN,G�RES�!0Q_<;3!4C_WA�471^�:OFF_ N�3wDELHLOGn285Aa2?i1@FN?�� -M���W+0�$Y $D�B� 6COMW!2MO� "0G_A.o	 \rVE�1�$F��A{$�O��D�B�CTMP�1_F�E2�G1_P�3�B�2�XD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYPuAHK�BD_S�B�1AG�N Gn $SLOT_NUM�JQPREV,DBU�� g1� ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�AETE�_OKRUS�P7_CRQ$;4�V�� 0LACIw�1�RAPk �1x@ME>@$D�V�Q��Pv�A{�BLv� OUzR ,mAЧ0�!� B� LM�_O�^eR�"CAsM_;1 xr~$ATTR4�NP� ANN�@5I�MG_HEIGH|Q�cWIDTH4�VT� �UU0F_�ASPECQ$�M�0EXP��@A�X�f�CFT ?X $GR� � �S�!�@B@NFL�I�`t� UIREx 3dTuGITCHCj�`N� S�d_L�`2�C�"�`EDlpE
� J�4S�0� �zsa�4 hq;G0 �� 
$WARNM��0f�!,P� �s�pN{ST� CORN�"�a1FLTR�uTRkAT� T�p H0ACCa1���{��ORI
`"S={R�T0_S�B�CHuG,I1 [ �Tp�"3I9�TYL12�pHK*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7j��8��9�CO�$ <� $6xK3� 1w`O_M�@�C/ t � E#63NGP�ABA� �c���ZQ���`���@nr��� ��P�0��`�,� �v�p�PzP�b26����"J�_)R��BC�J��3�JVP��tBS��}�Aw��"�@G CP_�*0OFSzR @�� RO_K8���aIyT�3��NOM_�0R�1ĥ3�PT� �� $���AxP��K}EX�� �0g0�I01��p�
$TF�a��C$MD3��T�O�3�0U� �� K�Hw2�C1|�	EΡg0wE{vF�vF�`�Pp@�a2 m
P$A`PU�3N)#�dR*��AX�!sDETAI�3BUFV��p@1� |�p۶�pPIZdT� PP[�MZ��Mg�Ͱj�F[�SIMQSI�"0��A.�r���kx Tp�|zM��P�B�FAkCTrbHPEW7�`P1Ӡ��v��MCd�� �$*1JB8�p<�*1DECHښ��H���-�c� � �+PNS_EMP���$GP���,P_���3�p�@Pܤ��TC��|r��0�s��b��0�� �B���!
���J�R� ��SEGFRR��Iv �aR�Tkp9N&S,�PVF4Ǳ>� &k�Bv �u�cu��aE�� !2��p+�MQ��E�SIZ�3����T��P�����>�aRSINF��� ��kq���������LX�����F�CRCMu�3CClpG��p� ��O}���b�1��������2�V�DxIC��C ���r����P��{� SEV �zF_�եF�pNB0�?�p�����A�! �r �Rx����V�lp�2ݠ�aR�t�,�g�_�R>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!��$SK��2GD  � �"�"�@�PR8� 
R��D���# l>�q1$��$��
+�L9$?(�V�)%@?R4C&_?R4gENE��'~?��AA�!RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@����C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!��DCS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�g ��QSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc �@Sp�i�a+ �j�fib��pOGIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�P6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6Cq~��DM�SWU. 8!�KgEYI��5�TM�10�s�qoA�vINޱE�Ca, / D��H7OST�P!4����<���<�°<��p<�E�M'���Z�D`SBL�� UL��0  ��	����DT��01 � $|��9USAMPL�@��/���決�$ I@|갯 $SUBӄ���w0QS�����#��SAV�����c�S< X9�`�fP$�0E!�� YN_B�#2 M0�`DI�d�pO|��m��#$F�R_I�C� �ENC2s_Sd3  ���< 3�9���� c����4�"��2�A9��ޖ5���`ǻ�@Q@K&D-!�a�AVER�q��λ�DSP
���PC�_�q��"�|�ܣ�V7ALU3�HE�(��M�IP)���OP5Pm �TH�*�D�S" T�/�Fb�;�d����d D��`��{ET6 H(rLL_DUǀ�a�@`��k���֠OT�"�U�/���q@@NO�AUTO70�!$}�x�~�@s��|��Cp���C� 2���z�L�� 8H *��L� ��� Բ@sv��`� �� ÿ� ��Xq��cq���q���q���7��8��9��0T���1�1 �1-�U1:�1G�1T�1aʕ1n�2|�2��2� �2-�2:�2G�2�T�2a�2n�3|�3R�3� �3-�3:�U3G�3T�3a�3nʅ4|�ͱ����9� <���z�ΓKI`����H硵��FEq@�{@: ,��&a?g P_P?��>�����E�@�ᶰ��QQ��;֐$�TP�$VARqI����,�UP2Q`3< W�߃TD��g����`������v����BAC�"= T2����$)�,+r³�p IFI��p�� �q M�P"�P�F�l@``>t ;h��6����ST� ���T��M ����0	��i���F����������kRt ����FOR�CEUP�b܂FL+US
pH(N��� ���6bD_CM�@E �7N� (�v�P��REM� Fa���@j���
K�	N���EFF/���@3IN�QOV���OVA�	TROV� DT)��DTMX:e �P:/���Pq�vXpCL�N _�p��@ ��	_�|��_T: �|�J&PA�QDI����1��0�Y0RQDm�_+qH���M���CL�d#�RIV�{�ϓN"EAR/�I�O�PCP��B�R��CM�@N 1b =3GCLF��!�DY�(��a�#5T��DG���� �%��&��SS� )�? �P(q1�1�`_(1"811�EC1�3D;5D6�GRA����@�����PW��ON2EBU�G�S�2�C`gϐ_?E A ��?����TERM:�5B�9ORIw�0C�9SM_-`���0�D�:A�9E�9UP>��F� -Qϒ�A�P�3�@B$S�EGGJ� EL�UU�SEPNFI���pBx��1@��4>DC$sUF�P��$����Q�@C���G�0T������SNSTj�P�ATۡg��APTH	J�A�E*�Z%qB\`@F�{E��F�q�pARxP<Y�aSHFT͢qA|�AX_SHOR$��>��6 @$GqPE���OVR���aZP�I@P@$U?r *aAGYLO���j�I�"���Aؠ��ؠERV ��Qi�[Y)��G�@R���i�e��i�R�!P�uASYM���uqA#WJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P���WkOR�@M��k0�SMT��G��GR��3�aPA�@���p|5�'�H � j��A�TOCjA7pP<]Pp$OPd�O�P�C�%�p�O!���RE.pR�C�AOX�?��Be5pR�E�ruIx'QG�e$PW�R) IMdu�RR_p$s��c�B Iz2�H8�=�_ADDR~H�H_LENG�BP�q�q:�x�R��So�mJ.�SS��SK������� ��-�SE�*��G2�HS�N�MN1K	�`j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ����Q8� ��OUPW3�bE_>�I��!q�a1�� ������|���������-���:���iIOX2S=�D�e��y^���L $��<p�!_OFF[r_�oPRM_�z�a�TTP_�H��M; (�pOBJ�"�p�G�$H�LE�C|��ٰN � 9�.*�AB_�T��
��S�`�S��LV��K�RW"duHITCOmU?BGi�LO�q����d� Fpk��GpSS� ���HW�h�wA��O.��`I�NCPUX2VISIO��!��¢.�á�<�á-� �IOL]N)�P 87�R'�^[p$SL�bd oPUT_��$dp��Pz �� F_�AS2Q/�$L D���D�aQT U�0]PA������PHY`G灱Z�̱5�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp����x��ٶ��UJ���S����NE�WJsOG�G �DIS��b&�KĠ��3T |���AV��`_�CTR<!S^�FLAGf2&�;LG�dU �n�:���3LG_SIZ���ň��=���FD��I����Z �ǳ� �0�Ʋ�@s��-ֈ�-ր=�-���-��0-�ISGCH_��Dq��N?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHrܘ�I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn��0I�BWUFF1XY��PT�$�� �v��Rf�x�`1�A�rYY���P �����pOS�1�2�3���_|�0Z �  ��aiE�*��IDX�dP�RhrO�+��AV&ST��R��Yz�~<! Y$EK&CK+���Z&m&�5�0[ L��o�0�� ]PL�6pwq�t^����t�L6�_ \ �����瀰�7��#�0C��] ��CLD�P��;eTRQLI��jd.�094FLG z�0r1R3�DM�R7Ɩ�LDR5<4R5ORG.���e2(`���V�8�.��T<�4�d^ ��q�<4��-4R5S�`T�00m��0DFRCLMC!D�?�?3I@���MIC��d_ d����RQm�q�DgSTB	�  �Flg�HAX;b �H>�LEXCESZr�RrBMup�a`�p�B�;d�rB`��`a��F_A�J��$[�O�H:0K�db \��ӂnS�$MB��LIБ~}SREQUIR�R�>q�\Á�XDEBUT��oAL� MP�c�b�a��P؃ӂ!BoAND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@qܮ�o� �SPS�T8� e�rLO�C�RI�p�EXfA�p��A�AOD�AQP�f X��ON��[rMF�����f )�"I��%�e��T���FX�@IGG� g �q��"E�0�h�#���$R�a%;#�7y��Gx��VvCPi�D'ATAw�pE:�y���RFЭ�NVh t_ $MD�qIёA)�v+�tń�tH�`��P�u�|��sANSAW}��t�?�uD��)�r�	@Ði �@CU��V�T0�A�oARR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2��RIN��v�<F?S�INTE����kE���,�V�����_Nl��ڂ��kDׄ�Rm�DIViFD�H�@ـn�$�V��'c!$���$Z�����~��[��oH �$�BELTb��!ACCEL+��ҡ���IRC�t����T</!��$PS�@#2L  �Ė83����x��� ��PATH���������3̒Vp�A_@�Q�.�4�B�C�_MGh�$D�DQ���G�$FW�h��p��m�����b�D}E��PPABNԗROTSPEED����00J�Я8��@���̐$USE_d��P��s�SY���c�A >qYNu@A�g��OFF�q�M�OUN�NGg�K�O9L�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I̒��4��\BݠVEO�w�Ͳ2�3_UPE�߳LOWL���00����D���BwP��� ��1RCʀƶMOSI�V�JRMO���@GP�ERCH  �OV��^��i�<!� ZD<!�c��d@�P��BV1�#P͑��L�0��EW��ĸUP��Ŝ���TRKr�"AYLOA'a�� Q-��̒<�1Ӣ`0 ��RT1I$Qx�0 MO���Ѐ�B R�0J��D��s��H����b�DUM2�(�S_BCKLSH_C̒��>�=�q� #�U��ԑ���2�t�]ACLALvŲ�1nМP�CHK00'%SD�RTY4�k��y�1�q_6#2�_UM�$Pj�Cw�_�SCL���ƠLMT_J1_LO��@���q��E�����๕�幘SPC��7������PCo���H� �PU�2m�C/@�"XT_�c�CN_��N��e���SFu���V�&#�� ��9�̒��=�C�u�SH6#��c����1�р��o�0�͑
��_�P�At�h�_Ps�W�_ 10��4�R�01D�VG��J� L�@J�OG|W���TORQU��ON*�Mٙ�sRH�L���_W��-�_=���C��I��I�IJ�II�F�`�JLAX.�1[�VC��0�D�BO1U�@i�B\�JRKU��	@D�BL_SMd�BM�%`_DLC�BGR�V��C��I��H�_� �*COS+\�(LN�7+X >$C�9)I�9)u*c,�)�Z2 HƺMY�@!�( "TH&-�)T�HET0�NK2a3I��"=�A CB6CB=�C�A�B(2061C�616SBC�T2N5GTS QơC� �aS$" �4c#�7r#$DUD�EX�1s� t��B�6���AQ|r�f'$NE�DpIB U�H\B5��$!��!A�%�E(G%(!LPH$U�2׵�2SXpCc% pCr%�2�&�C�J�&!�EVAHV6H3�YLVhJUVuKV�KV�KV�KV�KV�IHAHZF`RPXM��wXuKH�KH�KUH�KH�KH�IO2L�OAHO�YWNOhJO�uKO�KO�KO�KO
�KO�&F�2#1ic%��d4GSPBALA�NCE_�!�cLE6k0H_�%SP��T&��bc&�br&PFUL�C�hr�grr%Ċ1=ky�UTO_?�j�T1T2Cy��2N &�v�ϰctw�g�p�0(Ӓ~���T��O���>� INSEGv�!��REV�v!���DI�F��1l�w�1m�0OB�q
�����MIϰ1��LCHgWAR����AB&~u�$MECH,1�� :�@�U�AX:�P���Y�G$�8pn 
pZ��|���ROBR��CR̒��N��&��MSK_�`f�p� P Np_��R ����΄ݡ�1��Ұ�Т΀ϳ��΀"�IN��q�MTCOM�_C@j�q  �L��p��$NO�RE³5���$�7r 8� GR�E��SD�0ABF�$?XYZ_DA5A���DEBU�qI���Q�s �`$�COD�� ��k�F��f�$BUFIwNDXР  ���MOR��t $-�U��)��r�B������Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��E����͐OPWOܭŀv0��SY�SBU�@ʐ$SO!P����#�U"��p�PRUN�I�PA��DH�D����_O�U�=��qn�$^}�IMAG��ˀ��0P�qIM����I�N�q���RGOVCRDȡ:���|�P~���Р�0L_6p���Li��RB���0��M���EDѐF� J��N`M*��ཷ��˱SL�`ŀw x $OVSL�vwSDI��DEXm�@g�e�9w�����V� ~�N���w����Û���ȳ�M�o ���q<��� x �HˁE�F�ATUS
���C�0àǒ�çBTM����If�¿�4����(�ŀy �DˀEz�g���PE��r�����
���EXE��V��E�Y�$Ժ �ŀz @ˁ��UP�{�h�$�p��XN����9�H� ��PG"�{ h �$SUB��c�@_���01\�MPWAI2��P����LO��-��F�p�$RCV?FAIL_C�-��BWD"�F���DE�FSPup | Lˀ`�D�� U�UNI��S���RX`���_L�pP��M���P�ā}���� B�~���|��`ҲNN�`KET��y���P� $�~���0SIZE��ଠ{����S<�OR��FORMAT/p � F��ᖫrEMR��y�UqX���@�PLI7�~ā  $�P_SWI��Ş�_PL7�AL_ S�ސR�A��B��(0C��Df�$E�h����C_=�U�� � � ���~�J3�0�����TIA4��5��6��MOM������h �B�AD��*��* PU70NRW��W �U������ A$PI�6���	�� )�4l�}69��Q����c�SPEED�PG q�7�D�>D�� ��>tMt[��SAM�`痰>��MOV���$��p �5��5�D�1�$2�������{�Hip�IN?,{� F(b+=$�H*�(_$�+�+GAMM�f�1{�$GET��ĐH��D����
^pLIB�R�ѝI��$HIB��_��Ȑ*B6E��b*8A$>G086LW= e6\<G9�686��R���ٰV��$PGDCK�Q�H�_����;"��z�.%�7��4*�9� �$IM_SRO��D�s"���H�"�LE��O�0\H��6@��Q� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_�D�E��NO��C gA�Ҷ��@�$����I ��	�I� %Z[� �� RX" ��m���"�q �'"�8�Hӱ�t�W�UpS���Q�M��O㵐.'}q��C�g���@ʣ�ߑ���P�LM�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PLM���	� 0h�H�{�%X��O��z�Z�eT�M���� pS��C��O__0_B_�a:��_%�� |S��� �@	�v��v �@��ȯw�v��EM��% QmCbfr�B�ː��ftP��PM��Q]U� �U�Q���A-�QTH=�HO�L��QHYS�ES�,�UE��B��]O#��  ��P0��|�gAQ���ʠu�iZ���ŀ�ɂv�-�A;ӝROG��a2D�E�Âv�_�ĀZ�/INFO&��+�����b� �킍{ ((@SLEQ/ �#�����O�o���S`c0O�0�051EZ0NUe�_��AUT�Ab�COPAY��Ѓ�{��@M���N�����1�P�
� ���RGI�����X_�Pl�$�����`
�W��P��j@�G����EXT_CY�CtbCa�p�����h�_NA�!�$�\�<�RO�`]��� � m��P�OR�ㅣ���SReVt�)����DI �T_l���Ѥ{�ۧ�Шۧ �ۧ5٩6٩7�٩8��CaS�B쐒���$�F6���PL�A�A^�TAR���@E `�Z����9��d� ,(@FL�q`h��@YNL���Mz�C���PWR���쐔e�DELA�Ѱ�Y�pAD#q�ER.�QSKI�P�� ĕ�x�O��`NT!���P_x���ǚ@�b�p1� 1�1Ǹ�?� �?� �>��>�&�>�3�>�=9�J2R;쐷� 4��EX� TQ����ށ�Q���[�pKFд�8�RDCIf�� �U`�X}�R��#%M!*�0�)��$R�GEAR_0IO�TJBFLG�igpERa��TC݃����>��2TH2N���O 1�b��Gq �T�0 ����Mİ��`Ib���REuF�1�� l�h���ENAB��lcTPE?@���!(ᭀ ����Q�#�~�+2 VH� ��2�Қ��@�"�4�F�X�j�3���{��������j�4�Ҝ��
��.�@�R�j�5�ҝu�����P������j�6�Ҟ��@(:Lj�7���o�����j�8�Ҡ��"4�Fj�SMSK��R���a��E�At����MOTE�������@ "1��Q�I�O�5"%I��P��PsOWi@쐣  �D������h�쐤���Y"$DSB_SICGN4A�Qi�̰C�о�tRS232%��Sb�iDEVICE�US#�R�RPAR�IT�!OPBI�T�Q��OWCONTR��Qⱓ�R�CU� M�SUXTASK�3NB��0�$oTATU�P��IS@@쐦F�6�_�P�C}�$FREEFROMS]p�ai��GETN@S�UPD�l�ARB73P%0����� !m$U�SA���az9�L�EcRI�0f��pRY�5~"_�@f�P�1�!�6'WRK��D9�F�9ХFRIEND��Q4bUF��&�A@T�OOLHFMY5��$LENGTH_;VT��FIR�pqC��@�E� IUFI�N�R���RGI<�1�AITI:�xG�X��I�FG2�7G�1a����3�B�GPRR�DA��O_� o0e�I1RER�đ�3&����TC���AQJV�QG|�.2���F��1 �!d�9Z�8+5K�+5���E�y�L0�4�X ��0m�LN�T�3H@z��89��%�4�3G��IW�0�W�RdD� Z��Tܳ��K�a3d��{$cV 2��`H�1��I1H�02K2sk3K3Jci�a I�i�a�L��SL��RS$Vؠ�BV�EVk�(]V*R��� �,6Lc ���9V2F{/P:B��kPS_�Et�$rr8�C�ѳ$A0��wCPR���v�U�cSk�p� {��8��� 0��D�VX`�!�tX`�\`P�0P�Ё�
�5SK!/� �-qR��!�0���z�NJ AX�!h�A�@LlA��A�/THIC�1�������1TFE���q>��IF_CH�3A�I00�����G1�x�������9�Ɇ_J�F҇PR(���R�VAT�� �`-p��7@����DO�E���COU(��AX�Ig��OFFSE+�TRIG�SK��c@���Ѽ�e�[�K�Hk�<��8�IGMAo0�A�-��ҙ�ORG_�UNEV��� ��S�쐮d ��$������GROU��ݓTO2��!ݓwDSP��JOG'�L�#	�_P'�2OR�p��>P6KEPl�#IR�0�PM�RQ�AP�Q��E�0q�e����SYSG��"��PG��BRK*Rd�r�3�-�������ߒ<p�AD��ݓJ�BSO�C� N�DUM�MY14�p\@SV��PDE_OP3S�FSPD_OVR���ٰCO��"�OIR-��N�0.�Fr�l.��OV�SFc�2�f��F��!4�S���RA�"LCHDL>�RECOV��0��W�@M�յ�R�O3��_�0�s @�ҹ@VERE��$OFS�@CV� 0BWDG�ѴC��X�2j�
�TR�!���E_FDOj�MOB_CM��U�B ��BL=r0�w�=q�tV@fQ��x0sp��_�Gx���AM��k�J0������_M��2{�#�8$CA�{Й���8$HBK|1c�ыIO��.�:!aPPA"�N�3�^�F����:"�DVC_DB �C��d�w"����!�Ց1���ç�3����ATIO� �q0�qUC�&CAB� BS�PⳍP�Ȗ���_0c�SUBCP	Uq��S�Pa aáĀ}0�Sb��c��r"ơ$HW_C���:c��IcA�A-�l$U�NIT��l��AT�N�f����CYCL�ųNECA��[�F�LTR_2_FI`���(��}&��LP&������_SCT@SF�_��F����G���FqS|!�¹�CHAA�/����2��RSD��x"ѡb�r�: _T���PRO��O�� E%M�_��8u�q� u�q��DI��0e�RAILAC4��}RMƐLOԠdC��:anq��wq����+PR��SLQ\`f�C�ѷ 	��FUN9CŢ�rRINkP+a0�0 ��!RA� >R� 
Я�ԯW3AR�BLFQ���A�����DA`�����LDm0 �aB9��nqB�TIvrbؑ���PR�IAQ1�"AFS�P �!�����`%b����M�I1U�DFa_j@��y1°LME�{FA�@HRDY�4��Pn@RS@Q�0">�MULSEj@f�<b�q �X���ȑ���$.A$��1$c1Ó��߰� x~�EG0vpݓ�q!AR����09>B�%��A�XE��ROB��Wd�A4�_�-֣SY��h�!6��&S�'WR��r�-1���STR���5�9�E�� 	5B��=QB90�@6X������OT�0o ;	$�ARY8�w2h0���	%�FI��~;�$LINK��H��1�a_63�t5�q�2XYZ"� �;�q�3@��1�2�8%{0B�{D��� CFI��6G�0�
�{�_J��86��3aOP_O4Y;5�QTBmA"�B�C
�z�DU"�66CTURN3�vr�E`�1�9�ҍGFL�`@���~ �@�5<:7�^� 1�?0K�	Mc�68Cb�vrb�4�ORQ��X�>8 �#op������wq�Uf�8����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W���Tυ � ;����QH�!`�� ���U�Q�WkeK#kec�XER��	GE	0��S�dAWaǢ:D����7!�!AX �rB!{q��1u y-!y�pz�@z�@ z6Pz\Pz� z1 v�y�y�+y� ;y�Ky�[y�ky��{y��y�q�yDEBU��$����L�`!º2WG`  AB!��,��SV���� 
w���m���w����1 ���1���A���A��6Q ��\Q���!�m@��2.CLAB3B�U��x���S  Ð�ER���� � i$�@� Aؑ!p�PO��Z�q0w�^��_MRAȑ� d�  T�-�ER1R��TYz�B��I�V3@�cΑTO	Q�d:`L� �d2��]�X�C[! �� p�`T}0i��_�V1�r�a'�4�2B-�2<����@P�����F�$W��g��5V_!�l�$�P�����c��q"�	��SFZN_CFG_!� 4��?º�|��ų����@�ȲW �aV ��\$� � n���Ѵ��9c�Q��(��FA�He�,�XE�DM�(�����!s��Q�g�P{RV HEL}Lĥ� 56��B_BAS!�RSQR��ԣo �#S��T[��1r�%��2ݺU3ݺ4ݺ5ݺ6ݺ�7ݺ8ݷ��ROO0I䰝0�0NLK!�C�AB� ��ACK��IN��T:�1�@p�@ z�m�_PU!�CO� ��OU��P�� Ҧ) ��޶��T�PFWD_KAR�ӑ��RE~��P8��(�QUE������P
��CSTOPI_AL�����0&p���㰑�0SEMl�db�|�M��d�TY|�3SOK�}�DI����p�(���_TM\�MANRQ�ֿ0E�+�|�$KEYSWITCH&	����HE
�BEAT4��cE� LEҒ��
�U��FO�����_O_HOM�O�7REF�PPRz�(�!&0��C+�OA��ECO��B�rI�OCM�D8׵�p]���8�` � D�1$����U��&�MH��<�P�CFORC���� ���OM�  �� @V��|�U�,3P� 1-�`� 3�-�4��NPX_�ASǢ� 0ȰA�DD����$SI}Z��$VARݷ. TIP]�\�2�A򻡐���]�_�$ �"S꣩!Cΐ��OFRIF⢞�S�"�c���NF��V ��n` � x�`SI��TES�R6SSGL(T�2P&��AU�<� ) STMTQZ�Pm 6BW�P*S�HOWb��SV|�\$�� ���A00P�a�6�@@�J�T�5�	U6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	f0 u�	�0u�	�@u�[Pu%121?1�L1Y1f1s2��	2�	2�	2�	2��	2�	2�	22�2%222?2�L2Y2f2s3�P)3�	3�	3�	3��	3�	3�	33�3%323?3�L3Y3f3s4�P)4�	4�	4�	4��	4�	4�	44�4%424?4�L4Y4f4s5�P)5�	5�	5�	5��	5�	5�	55�5%525?5�L5Y5f5s6�P)6�	6�	6�	6��	6�	6�	66�6%626?6�L6Y6f6s7�P)7�	7�	7�	7��	7�	7�	77�7%727?7�,i7Y7Fi7s��&��VP�UPD>��  ��|�԰��YSLOǢ� � z��и����o�E��`>�^t��АAcLUץ����CU��z�wFOqID_L��ֿuHI�zI�$F�ILE_���t���$`�JvSA��� �h���E_BLC�K�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� ��LA��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ� ��TBCu�C� ��X -$�LENi��v�������I��G�LOW_A�XI�F1��t2�X�M����D�
 ��I�� ��}�TOR�����Dh��� L�=��⇒�s���#�_�MA`�ޕ��ޑT#CV����T��� &��ݡ����J�����IJ����Mo���J�Ǥ� �������2���� v�����F�JK���VKi�Ρv�Ρ3f��J0�ңJJڣ;JJ�AALң�(ڣ��4�5z�&��N1-�9���␅�L~�_Vj��+p����� ` �GRO�U�pD��B�NF�LIC��REQ�UIREa�EBU`A��p����2¯������c�� �\��APPR��C����
�EN�CsLOe��S_M �v�,ɣ�
���� ���MC�&���Ng�_MG�q�C� ��{�9���|�BRK�z�NOL��|ĉ R��_LI|��Ǫ�k�	J����P
���ڣ��@���&���/���6�ń6��8�����Ə� ��8�%�xW�2�e�PATHa׀z�p�z�=�vӥ�ϰ�6x�CN=�CA����l�p�IN�UC���bq��CO�UM��YZ������qE%���2�������PAYLO�A��J2L3pR_AN��<�L��F�B��6�R�{�R_F2LgSHR��|�LOG���р��ӎ���ACRL_u�������.���9H�p�$H{���FLEX
�s�J>�� :�/� ���6�2�����;�M�_�F16����n��� ������ȟ��Eҟ� ����,�>�P�b�� �d�{����������H��5�T��X�� v���EťmFѯ �������&�/��A�S�e�D�Jx�� � ������j�4pcAT����n�EL S �%øJ���ʰ;JE��CTR�Ѭ��TN��F&��HA_ND_VB[
�ܤpK�� $F2�{�6� �rSWi���r�U��� $$	Mt�h�R��08��@<b 35��^6A�p3�kƈ�q{9t�A�̈p��A���A�ˆ0��U���D*��D��P��G��ICST��$A��$AN��DYˀ�{�g4�5D� ��v�6�v��5缧�^�@��P������#�,�5�>�
�K�� &0�_�ER!V9�SQOASYM��] ��¤��x��ݑ���_SHl�������sT�(����(�:�JA���S�pcir��_VI�#�Oh9�``V_UN!I��td�~�J���b �E�b��d��d�f��n���������uN����2�H�������"CqEN� a�D	I��>�ObtC�Dpx��� ��2IxQA ����q��-��s �� ������ ��OMME��rr/�TVpPT�P ���qe�i����P�x ���yT�Pj� $�DUMMY9�o$PS_��RFq�s  ��:� �8��!~q� X�����K�STs�ʰSB}R��M21_Vt�8$SV_ERt�qO��z���CLRx�EA  O�r?p? Oր� � D $�GLOB���#LO ��Յ$�o��P�!wSYSADR�!�?p�pTCHM0 �� ,����W_NA��/�e�$%�SR��l (:]8:m�K6�^2 m�i7m�w9m��9���� ���ǳ���ŕߝ�9ŕ ���i�L���m���_�_�_�Tr�XSCSRE�ƀ�� ��3STF���}�pТR6�C�] _v AŁ�� T����TYP �r�K��u�!u����O�@IS�!���tC�UE{t� �����H�S���!R�SM_�XuUNE�XCEPWv��CpS_��{ᦵ�ӕ���÷���COU ���o 1�O�UET��փr���PROG�M� FLn!$CMU��PO*q�����I_�pH;� �s 8��N�_HE
p���Q��pRY �?���,�J�*���c�?�OUS�� �� @d���$B�UTT��R@���C�OLUM�íu�S�ERVc#=�PAN�Ev Ł� � N�PGEU�!�F��~9�)$HELP��^WRETER��)� ����Q�������@� P�P �IN��s�PNߠw v��1����� ����LN�� �䟀�_��k�$H��M TEX�#�����FLAn +REL�V��D4p�������M��?,��ӛ$�����P=�USR�VIEWŁ� <�d��pU�p0NFyIn i�FOCU��ni�PRILPm+��q��TRIP)��m�UNjp{t� �QP��XuWARN|Wud�SRTOLS��ݕ�����O|SO;RN��RAUư��9T��%��VI|�zu�� $�P�ATHg��CAC�HLOG6�O�LIMybM���'��"��HOST6�!��r1�R�OBOT,5���IMl� D�C� g!��E�L���i��VCPU_AVA�ILB�O�EX7�!BQNL�(���A�� Q���Q ��ƀ��  QpC���@_$TOOL6�$��_JMP� �<I�u$SS�!$}TPVSHIF��|s�P�p�6�s����R���OSURzW�pRADIz��2�_�q�h�g! ؎q)�LUza$�OUTPUT_BM��IML�oR6�(`)�@TIL<SCO�@Ce�;�� 9��F��T��a�� o�>�3�����w�I2u���V�zu���%�DJU��|#�/WAIT����ک�%ONE��Y�BOư ��� $@p%�C�SB�n)TPE��NEC���x"�$t$���*B_T��R��%�qR� $���sB�%�tM�+���t�.�F�R!݀��O�Pm�MAS�_DUOG�OaT	�D�����C3S�	�O2DELcAY���e2JO�� n8E��Ss4'#J�aP60%�����Y_��O2�$��2���5��`?� �=pZABC~S��  $�2��J�
���$$C�LAS������AB���'@@VI�RT��O.@ABS��$�1 <E�� < *AtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v�����M@�[�AXLրK�*B�ndC  ���IN��ā��PRE������LARMRECOV <Il䂥�NG�� \K	 =#�
J�|\�M@PPLIC��?<E�E��Handlin�gTool �� �
V7.50P�/28 *A��^���
�_SW UP*A� F��F0ڑ����A��~�� 20�К*A���	Ց��h�jFB �7DA5��  ~'@�^@�𞝓None������� ��T�y�*A4�]x��P_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ��i�n�����#B)B ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��e��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���oe�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� ��PB�Z?����5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`��S:��r������Up�_)o�S  K�3Ph���R�PX�_mo8j����a�Oko�o9i�(�+(�9!Rhg�o�o�l�Kof�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`(ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCPU�eB��CF��;.<C����C5`SXE@D��nyDQ��D���>��D�;D�����F��>F�$�G}RB�7Gzր��SY��)!�vqG���Em�U(�.��(�(�1�<�q�G�x2��eҢ �� a�D�j�怀ES\E@EX��EQ�EJP� F�E�F�� G�ǎ^F� E�� FB�� H,- Ge�߀H3Y��� � >�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE ��O@b 
�(�;��"�  <�6�z�Rb���?�j�C4�)�SZm� W��{�Jm�C��B-G�Cu��@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"�� , 
�^��P�o xvf`MT�I^��rl@�:sONTImM������Zv�i
õ�cMOTN�END���dREC�ORD 1(R�8a��ua�O��q� �sb�.�@�R��xZ� ������ɏۏ폄� ��#���G���k�}��� ��<�ş4��X��� 1�C���g�֟������ ��ӯ�T�	�x�-��� Q�c�u���������� >����)Ϙ�Mϼ� F�࿕ϧϹ���:��� ����%�s`Pn&�]�o� �ϓ�~ߌ���8�J��� ��5� ��k����� ���J�����X��|� ��C�U�����������0�����	��dbTOLERENCqdsBȺb`L�͐P�CS_CFG �)�k)wdMC�:\O L%04dO.CSV
�Pc��)sA �CH� z�P)~���hM�RC_OUT �*�[�`+P SG�N +�e�r���#�10-MAY�-20 10:4�7*V27-JAN�j21:48�k? P;����)~�`pa�m��PJPѬ�VERSION� SV2�.0.�6tEFLOGIC 1,�[/ 	DX�P7)��PF."PROG_�ENB�o�rj UL�Sew �T�"_WRSTJNEp�V�r�`dEMO_OPT?_SL ?	�es�
 	R575)s7)�/??*?<?|'�$TO  �-د�?&V_@pEX�Wd�u�3PAT�H ASA\p�?�?O/{ICT�a-Fo`-�gds�egM%&ASTBF_TTS�x@�Y^C��SqqF�P�MAU� t/XrMS%WR.�i6.|
S/�Z!D_N�O0_�_T_C_x_g_�_�tSBL_FAUL"y0�[3wTDIAU �16M6p�A�1234567G890gFP? BoTofoxo�o�o�o�o �o�o�o,>Phb�S�pP�_ ���_s�� 0`�� ���)�;�M�_�q� ��������ˏݏ��|�)UMP�!� �^�TR�B�#+�=��PMEfEI�Y_T�EMP9 È�3p@�3A v�UNI�.�(YN_BRK �2Y)EMGDI_STA�%W!b�ՐNC2_SCR 3��1o"�4� F�X�fv���������#��ޑ14���@�)�;�����ݤ5�����x�f	u� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/߭P�b� t�� ��xߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N���r��� ������������ &8J\n��� �����"`� FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/4?,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O?�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�O�O�o �o�o
.@Rd v������� ��*�<�N�`�r��� �o����̏ޏ���� &�8�J�\�n����������ȟڟ����H�E�TMODE 16v��� ���ƨ
R�d�v�נR�ROR_PROG7 %A�%�:߽��  ��TABLE  A�������#�L�RRSEV_?NUM  ��Q���K�S���_�AUTO_ENB�  ��I�Ϥ_N�Oh� 7A�{��R�  *����J��������^�+��pĿֿ迄�HISO��͡I�}�_ALM �18A� �;�����+�e�wωϐ�ϭϿ��_H���  A���|��4��TCP_VER �!A�!����$E�XTLOG_RE�Q��{�V�SI�Z_�Q�TOL  �͡Dz��=�#׍�XT_BW�D����r���n�_D�I�� 9���}�z�͡m���STE�P����4��OP_�DO���ѠFA�CTORY_TU�N�dG�EATU�RE :�����l�Hand�lingTool� ��  - C�English� Diction�ary��ORDE�AA Vis��� Master����96 H��n�alog I/O����H551��u�to Softw�are Upda�te  ��J��m�atic Bac�kup��Part�&�groun�d Edit�� � 8\apC_amera��F���t\j6R�ell����LOADR�o�mm��shq��T7I" ��co���
! o���pa�ne�� 
!���tyle se�lect��H59��nD���onit�or��48����t�r��Reliab����adinDiagnos"�����2�2 ual �Check Sa�fety UIF� lg\a��ha�nced Rob� Serv q �ct\��lUse�r FrU��DI�F��Ext. D�IO ��fiA �d��endr E�rr L@��IF��r��  �П�9�0��FCTN M�enuZ v'��7}4� TP In���fac  SU_ (G=�p��_k Excn g��3��High-S�per Ski+� � sO�H9 � mm�unic!�onsg�teur� �����V����coknn��2��EN���Incrstr�u���5.fd�KAREL C�md. L?ua�A� O�Run-;Ti� Env����K� ��+%�s#�S�/W��74��Li�censeT� � (Au* ogB�ook(Sy��m�)��"
M�ACROs,V/�Offse��ap���MH� ����pf�a5�MechStop Prot��� d�b i�S�hif���j54�5�!xr ��#��,��lb ode �Switch��mK\e�!o4.�&� pro�4��g���Multi-�T7G��net.�Pos Re�gi��z�P��t� Fun���3 9Rz1��Numx ������9m�1�  A�djuj��1 J�7�7�* ����6t�atuq1EIKoRDMtot��_scove�� ���@By- }ues�t1�$Go� � U5\�SNPX b�"���YA�"LibAr����#�� �$�~@h�pd]0�Jt�s in VCC!M�����0�  �u!Ξ�2 R�0�/I��08��TMIL{IB�M J92�@�P�Acc>�F�9=7�TPTX�+�B�RSQelZ0�M8� Rm��q%��69�2��Unexce{ptr motnT  CVV�P���KC����+-��~K�  II)�VSP� CSXC�&.c��� e�"�� t�@�Wew�AD �Q�8bvr nmeYn�@�iP� a0�y�0�pfGrid~Aplay !� �nh�@*�3R�1M-1�0iA(B2015 �`2V"  F����scii�loa�d��83 M��l�����Guar�d 'J85�0�mP'�L`����stuaPat�&]$Cyc���|0�ori_ x%Dat�a'Pqu���ch��1��g`� j� RLJam�5���I_MI De-B(\A^�cP" #^0C�  etkc^0a�sswo%q�)65�0�ApU�Xnt\��Pven�CTq�H�5�0YEL?LOW BO?Y���� Arc�0vis���Ch�Weld�Qcial4Izt��Op� ��gs�` �2@�a��poG yRjT1 NE�#3HT� xyWb��#! �p�`gd`����p\� =P��JPN� ARCP*PRx�A�� OL�pwSup̂fil�pp��J�� ��cro�6�70�1C~E�d��SuS�pe�tex�$Y �P� So7 t� /ssagN5 <Q�B�P:� �9 "0�Qr�tQC��P�l0dpn�笔�rpf�q�e��ppmasc�bin4psyn��' ptx]08�H�ELNCL V�IS PKGS �Z@MB &��B� J8@IPE �GET_VAR �FI?S (Uni�� LU�OOL: �ADD�@29.F�D�TCm���E�@D�Vp���`A�ТNO� WTWTEST� �� ��!��c�F�OR ��ECT ��a!� ALSE �ALA`�CPMO�-130��� b D�: HANG F�ROMg��2��R�709 DRAM� AVAILCH�ECKS 549���m�VPCS S�U֐LIMCHK���P�0x�FF P�OS� F�� q�8-12 CH�ARS�ER6�OG�RA ��Z@AVE�H�AME��.SV���Вאn$��9�m� "y�TRCv� �SHADP�UPD�AT k�0��ST�ATI��� MU�CH ���TIM�Q MOTN-0�03��@OBO�GUIDE DAUGH���b��@$Gtou� �@C� �0���PATH�_�M�OVET�� R6�4��VMXPAC�K MAY AS�SERTjS��CY�CL`�TA��BE COR 71�1�-�AN��RC O�PTIONS  ��`��APSH-1N�`fix��2�SO���B��XO򝡞�_TP��	�i��0j��du�{byz p wa���y�٠HI������U��pb XSPD T�B/�F� \hch�ΤB0���END�C�E�06\Q�p{ s>may n@�p�k��L ��traff#�	� ��~1�from sysvar scr�0qR� ��d�DJU����H�!A��/��S?ET ERR�D��P7����NDAN�T SCREEN� UNREA V�M �PD�D��PA����R�IO J�NN�0�FI��B���GROUNנD� Y�Т٠�h�S�VIP 53 QS���DIGIT V�ERS��ká�NE�W�� P06�@C�1IMAG�ͱ���8� DI`���p�SSUE�5��EP�LAN JON� gDEL���157QzאD��CALLI�ॡQ��m���IPN�D}�IMG N9� PZ�19��MN;T/��ES ���`wLocR Hol߀�=��2�Pn� PG:t��=�M��can������С: 3D �mE2view d3 X��ea1 �0�b�pof Ǡ"H�Cɰ�ANNOT� ACCESS �M cpie$Etn.Qs a� loMd�Flex)a:��w^$qmo G�sA9�a-'p~0��h0pa���eJ AUTO-�0��!ipu@Т<ᾡ�IABLE+� �7�a FPLN: �L�pl m� M�D<�VI�и�WI�T HOC�Jo�~1Qui��"��N���USB�@�Pt & remov����D�vAxis F�T_7�PGɰCP�:�OS-144� � h s 26�8QՐOST�p  �CRASH DU���$P��WORD�.$�LOGIN̈P��P:	�0�046 issueE��H�: Slow� st�c�`6Й���໰IF�IM�PR��SPOT:�Wh4���N1STY<��0VMGR�b�N�CAT��4oRR�E�� � 58t�1��:%�RTU!Pre -M a�SE:�@!pp���AGpL��9m@all��*0va�OCB WA����"3 CNT0 �T9DWroO0al�arm�ˀm0d �t�M�"0�2|� o�Z@OME<�� ���E%  #1-�SR�E��M�st}0g �    5KA�NJI5no M�NS@�INIS�ITALIZ'� E�f�we��6@� �dr�@ fp "~��SCII L�afails w�>�SYSTE[��i��  � Mq�1�QGro8�m n@�@vA����&��n᰼0q��RWRI O�F Lk��� \r�ef"�
�up� d�e-rela�Qd� 03.�0SSc}hőbetwe4�IND ex ɰTPa�DO� l�y �ɰGigE�s�operabil.`p l,��HcB�̚@]�le�Q0cf�lxz�Ð���OS� {����v4pfigi GLA�$�c2��7H� lap�0A[SB� If��g�2 l\c�0�/��E�� EXCE �㰁�P���i�� Do0��Gd`]Ц�fq��l lxt��EFal��#0�i�O�Y��n�CLOS��SR�Nq1NT^�F�U�FqKP�ANIO V7/ॠ1�{����DB �0��ᴥ�;ED��DET|�'�� �bF�NLINEb�BUG�T���C"RLIB��A���ABC JARK�Y@��� rkey��`IL���PR��N\��ITGAR� D$��R �Er *�T���a�U�0��h�[�Z�E V� TAS�K p.vr�P�2" .�XfJ�srn8�S谥dIBP	c�v��B/��BUS��UNN� j0-�{�d�cR'���LOE�wDIVS�CULs0$cb����BW!���R~�W`P�����ITd(঱tʠ�OF���UNEXڠ+���p��FtE��SVEM�G3`NML 50�5� D*�CC_SAFE�P*� �ꐺ� PET��'P�`�gF  !���IR����c i S>� K���K�H GUN�CHG��S�MEKCH��M��T*��%p6u��tPORY_ LEAK�J����SPEgD��2Vw 74\GRI�x�Q�g��CTLN��TRe @�_�p ���EN'�IN�����0�$���r��T3)�iԗSTO�A�s�L���͐X	���q��Y� ��TO2�J m���0F<�K����DU��S��O��3 �9�J F�&���SSVGN-1#I���'RSRwQDAU�Cޱ � �T6�g��� 3�]�~��BRKCTR/"� �q\j5��_�QܺS�qINVJ0D ZO�Pݲ���s��г��Ui ɰ̒�a�DU{AL� J50e��x�RVO117 AW�TH!Hr%�N�7247%�52��|�&aol ���R���at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���Md��Rǰt� \fosB�A�0Np�c�����{�U��ROP 2��b�pB��ITP4aM��b !AUt �c0< � plete��N@� z1^qR�635 (Acc_uCal2kA���I) "�ǰ�1a\�Ps��ǐ� bЧ0�P򶲊���ig\�cbacul "A3p_ �1��ն���_etaca��AT����PC�`�����_p�.pc!Ɗ��:�circB���5��tl��Bɵ�:�fm+�Ί�V�b�ɦ�r�?upfrm.����ⴊ�xed��Ί�~�'pedA�D �}b�ptlibB�� ߆_�rt��	Ċ�_0\׊ۊ�6�fm�݊��oޢ�e��̆Ϙ���c��Ӳ�5�j>�����tcȐ��	�r����emm 1��T�sl^0���T�mѡ�#�rm�3��ub Y�q�st�d}��pl;�&�c1kv�=�r�vf�䊰���9�vi����u�l�`�0fp�q �.yf��� daq; �i Data Ac_quisi��n��
��T`��1�8�9��22 DMCM RRS2Z��75��9 3 Rg710�o59pq5\?��T "���1 (D�T� n k@��������E Ƒȵx��Ӹ�etdmm F��ER����gE<��1�q\mo?۳ �=(G���[(

�2�` ! �@J�MACRO��Sk�ip/OffseP:�a��V�4o9� &qR662���Rs�H�
 6Bq8�����9Z�43 J�77� 6�J783�o ��n�"v��R5IKCBq2� PTLC�Zg� R�3 (�s,� �������03��	зJԷ\sfm�nmc "MNM�C����ҹ�%mnf�FMC"Ѻ0ª etmcr� �8����� ,��lD�l �  874\prdq>,jF0����axisHPro�cess Axe�s e�rol^P�RA
�Dp� 56 �J81j�59� 5�6o6� ���0w�6�90 98� [!IDV�1��2(x2��2ont�0�
�����m2���?C��etis "ISD��x9�� FpraxRA�M�P� D��de�fB�,�G�isb/asicHB�@޲�{6�� 708�6
��(�Acw:�����@�D
�/,��AMOX��  ��DvE��?;T��>Pi� RAFM';�]�!PAM�V�W�Ee�U0�Q'
bU�75�.��ceNe� nterface^�1' �5&!54�K��b(Devam±�/�#��Э/<�Tane`"D�NEWE���btpd/nui �AI�_s~2�d_rsono����bAsfjN��bdv_arFvf�xhp�z�}w��hkH9xs�tc��gAponlGzv{�ff��r ���z�3{q'Td~>pchampr;re�p� ^5977� �	܀�4}0��mɁ�/������lf�!�pcc7hmp]aMP&B<�� �mpev������pcs��YeS~�� Macro�O	D��16Q!)*�:$��2U"_,��Y�(PC ��$_;������o|��J�gegemQ@�GEMSW�~ZG�g�esndy��OD�n�dda��S��syT�Kɓ�su^Ҋ����n�m���L��  �	��9:p'ѳ޲���spotplus�p���`-�W�l�J�s⽱t[�׷p�key �ɰ�$��s�-Ѩ�m�~��\featu 0�FEAWD�oolo�srn'!2 �p���a�As3��tT�.� (N. A.)��!e!�J# (j�,��oBIB�o�D -�.�n��k9�"K��u[-�_���}p� "PSEq�W����wop "sEЅ�&�:�J����� �y�|��O8��5��R ɺ���ɰ[��X�� �����%�(
ҭ�q HL�0k�
�z�a !�B�Q�"(g�Q �����]�'�.����ɀ&���<�!ҝ_�#��tpJ�H�~Z��j����� y������2��e��� ���Z����V��!%���=�]�͂��^2�@i[RV� on�QYq͋JF0� 8ހ�`�	�(^�dQueue���X\1�ʖ`�+F1�tpvtsn��N�&��ftpJ0v �R�DV�	f��J1 Q4���v�en��k/vstk��mp��~btkclrq���get�����r��`kack8�XZ�strŬ�%��stl��~Z�np:!�`���q/��ڡ6!l�/Yr�mc�N+v3�_� ���l�.v�/\jF��� �`Q�΋ܒ��N50 (FRA���+��͢frap�arm��Ҁ�} 6��J643p:V�E�LSE
#�VA�R $SGSYS�CFG.$�`_U?NITS 2�DG0~°@�4Jgfr��4A�@FRL-��0ͅ�3 ې���L�0NE�:� =�?@�8�v�9~Qx3�04��;�BPRS�M~QA�5TX.$VNUM_OL��85��DJ507��l�? Functʂ"q�wAP��琉�3 HH�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6 N�kAP����S��"TPPR���Q.A�prnaSV�ZSx��AS8Dj510U�-�`cr�`8 ��ʇ��DJR`jYȑH � �Q �PJ�6�a21��48AAVM 5�Q�b0 lB�`TUP� xbJ5459 `b�`616���0VCAM 9��CLIO b1��5 ���`M�SC8�
rP R`\�sSTYL �MNIN�`J62�8Q  �`NRExd�;@�`SCH ���9pDCSU Me�te�`ORSR �Ԃ�a04 kR_EIOC �a5�`542�b9vpP<� nP�a�`�R�`7�`��MASK H�o�.r7 �2�`O'CO :��r3��p�b�p���r0X��a�`�13\mn�a39 HRM"�q�q�ҿLCHK�uO�PLG B��a03� �q.�pHCR �Ob�pCpPosi��`fP6 is[rJ�554�òpDSWĤbM�D�pqR�a37� }Rjr0 �1�s4i �R6�7��52�rs5 �2�r7 1� �P6���Regi��@T�uFRDM��uSaq%�4�`93�0�uSNBA�uSwHLB̀\sf"p�M�NPI�SP{VC�J520���TC�`"MNрT�MIL�IFV�P�AC W�pTPT�Xp6.%�TEL�N N Me�0�9m3UECK��b�`UFR�`��V�COR��VIPL:pq89qSXC�S�`�VVF�J�TP ��q��R626l�u� S�`Gސ�2�IGUI�C��PG�St�\ŀH863`�S�q�����q34sŁ684���a��@b>�3 :B��1 \T��96 .�+E�g51 y�q53�3f�b1 ���b1 n��jr9 ���`VAT9 ߲�q75 s�F�<�`�sAWSM��`�TOP u�ŀR582p���a80 
�ށgXY q���0 ,b��`885�QXрO�Lp}�"pE࠱tp��`LCMD��ET3SS���6 �V��CPE oZ1�V�RCd3
�NLH�h���001m2Ep��3� f��p��4 /1�65C��6l���7zPR��008 tB~��9 -200�`�U0�pF�1޲1 ��޲2L"���p��޲y4��5 \hmp~޲6 RBCF�`0ళ�fs�8 �Ҋ���~�J�7 rbc	fA�L�8\PC�����"�32m0u�n�K�R�ٰn�5 5EW�
n�9 z��40Y kB��3 ��6ݲ��`00iB/��6$�u��7�u��8 µ������sU0�`�t �1 05\rb��2 E���K���j�2��5˰��60��a�HУ`:�63�jAF�_����F�7 ڱ݀H�80�eHЋ��cU0��I7�p��1u��8u��9 73�������D7� ��5t�9+7 ��8U�1��2J��1�1:���h���1np�"��8(�U1��\pyl��,࿱�v ��B�854��1hV���D�4��im�с1�<���>br�3�pr�4@pGPr�6 !B���цp��1�����1�`͵155ض1g57 �2��62�S����1b��2����1Π"�2���B�6`�1<c�4 L7B�5 DR��8_�{B/��187 u�J�8 06�90� rBn�1 (��202 0EW,ѱ�2^��2��90�U2��p�2��2 b��4:��2�a"RB����9\�U2�`w�l���O4 60Mp��7��`����b�s
5 ���3����pB"9 3a ����`ڰR,:�7 �2��V�2��5@���2^��a^9��B�qr����n�5����5᥁"�8a�Ɂ}Չ5B���5����`U�A���� ��86 �6 S�0��5�p�2�#�529 �2^�Tb1P�5~�2`P���&P5��8��5��u�!�5��ٵ5+44��5��R�ąPa nB^z�c (�a4�����U5J�
V�5��1�1^��%������5 b21���gA��58W8-2� rb��5N�E�G5890r� 1�95 �"������c 8"a��|�L ���!J"E5|6��^!�6���B�"8�`#��+�8�%�6B�AME�"1w iC��622�B�u�6V��d� 4��8�4�`ANRSP�e?/S� C�5� �6� ��� \� �6� ��V� 3t��� TG20CA�R��8� pHf� 1DH�� AOE�� �� ,�|�� �0\�� �!64K��ԓrA� �1� (M-7�!/50T�[PM��P�Th:1�C�#Pe� �3��0� 5`M75T1"� �D8p� �0Gc�� u�4��i1-710i�1� Skd�7j�z�?6�:-HS,�  �RN�@�UB�f�X�=m75sA*A6a�n���!/CB�B2.6A �0;A�CIB�A�2P�QF1�UB2�21� �/70�S� �4��� �Aj1�3p���r�#0 B2\m*A@C@��;bi"i1K�u"A~A�AU� imm7c7@��ZA@I�@�Df�Ab�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A��EA�5B�4>\77
B7=Q�D�2�Q$B�E)7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E"l7�@7�A
1�E�V~`��W2%Q�R9ї@0L_�#����"A����b��H3s=rA/2 �R5nR4�74rNUQ1�ZU�A�s\m9
1M�92L2�!F!^Y�ps�� 2ci��-?�qhimQ�t  w043�C�p�2�mQ�r�H_ �H20��Evr�QHsXBSt62�q`s����� ��P�xq350_*A3I)�2�d�u0�@� '4kTX�0�pa3i1�A3sQ25�c��s�t�r�VR1%e�q0 
��j1��O2 �A �UEiy�.�‐ �0C2h20$CXB79#A�����M Q1]�~�� 9 �Q��?PQ��qA!Pvs � 5	15aU���?P�Ņ���ဝQ9A6�zS*�7�qb5�1��8��Q��00P(��V7]u�aitE1���ïp�?7� !?�z��rbUQRB1PM=�Qa9p��H��QQ�25L��@�����Q��@L���8ܰ��y00\r�y�"R2BL�tN�  ��� �1D�l�2�qeR�5���_b�3�X]1/m1lcqP1�a�ED�Q� 5F����!5���@M-16Q�� f� ��r��Q�e� ��� PN�LT_�1��i1��9453��@�e�|�b1l>F1u*AY2�
��R8�Q���RJ�J3�D}T� 85
Qg�/0��*A!P� *A�Ð𫿽�2ǿپ6t�6=Q���P�X���� AQ� g� *ASt]1^u�ajrI�B ����~�|I�b��yI�\m�Qb�I�uz�A��c3Apa9q� B6S���S��m���}�85�`N�N�   �(M���f1���6��P��161��5�s`҃SC��U��A����5\set06c��f��10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C����5�B��B��h`�F��� X0���A:���C�M��!AZ��@��4�6i����� e�O�-	���f 1��F �ᱦ�1F�8Y	���T6HL3��BU66~`���U�dU�9D20Lf0��Qv�  ��fjq��N������ 0v
� ��i	�	��72lqQ2�������� \chngmOove.V��d��|��@2l_arf 	�f~��6���� ��9C�Z���~���kr41 S���0��V���t�����U�p7nuqQ%�A]��V�1\�Qn�BJ�2W�EM!5���)�#:�64��F�e50S�\��0�=� PV���e�������E�����m7shqQSH"U��)��9�!A��(���� ,�l�����TR1!��,�6�0e=�4F�����2��	 R-������ �����Ж��4���LSR�)"�!lO�A��Q�) %!� 16�
U/��2�"2�E��9p���2X� SA/Ai��'�
7F�H�@ !B�0��D���5V� �@2cVE��p��T��pt갖�1L~E�#�Fd�Q��9E�#De/��RT��59���	�A�E�iR������9\m20�20��+�-u�19r4�`�E1�=` O9`�1"ae��O��2��_$W}am41��4�3�/d1c_std��1)�!�`�_T��r�_ 4\jdg�a�q�PJ%!~` -�r�+bgB��#c'300�Y�5j�QpQb1�bq��vB��v�25�U�����qm43� �Q<W�"Ps� �A��e����t� i�P�W.��c�F�X.�e�kE14�4y4�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf��`coWo!\�2a��K2A;_2��QW2�`bF�(�V11�23�`���X5�Ra21�J�*9�a:88J9X�l5�m1a첚��*���(85�&��������P6���R,52&A����,fA9IfI'50\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP 1��vB)e�m�����ު1p� �1D��l�27�F�KAR�EL Use S���FCTN��� �J97�FA+�� �(�Q޵�p%�)?�Vj�9F?(�j�Rtk208 "Km�6Q�yB�j��iæPr�9�sx#��v�krcfp��RCFt3���Q��k�cctme�!ME�g����6�mainj�dV�� ��ru��kDº�c���o����&J�dt�F �»��.vrT�f�����E�%�!��5�FRj73�B�K���UER�HJn�O  J�� (ڳF���F�q�Y�&T��`p�F�z��19�tkvBr���V�h�9p�E�y�<�k������;�v���"CT��f���� )�
І��)�V	�6� ���!��qFF��1q� ��=�����O�?�$"����$��je���TC�P Aut�r�<5�20 H5�J5�3E193��9��96�!8��9��	 �B�574��52�J:e�(�� Se%!Y������u��ma�Pqtool�ԕ�����~�conrel�F�trol Rel�iable�RmvCU!��H51�����8 a551e"�CNRE¹I��c�&��it�l\s�futst "UaTա��"X�\u�� g@�i�6Q]V0�B,Eѝ6A� �Q�)C ���X��Yf�I�1|�6s@6i��T6I U��vR�d�
$e%1���2�C58�E6��8`�Pv�iV4OFH58SOteJ� mvBM6E~O58�I�0�E�#+@� &�F�0���F�P6a����)/++�</N)0\�tr1�����P ,�lɶ�rmask�i�msk�aA���k�y'd�h	A	�P�sD�isplayIm��`v����J887# ("A��+Heůצprds��Iϩǅ�Uh�0pl�2�R2���:�Gt�@��PRD �TɈ�r�C�@Fm��D��Q�AscaҦ� �V<Q&��bVvbrl �eې@��^S��&5U�f�j8710�yl 	��Uq���7�&�p��p��P^@�P�firmQ����Pp�2�=b�k�6�r�3��6��t7ppl��PL���O�p<b�ac�q	��g1�J�U�d�J��gait_9e��Y�&��Q����	�Shap��e?ration�0��R67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G����qF�205p�5pS���Ձ�retsap��BP�O�\s� O"GCR�ö? �q/ngda�G���V��st2axU��Aa]��bad�_�btputl/�&�e�>��tplibB_���=�2.����5���c3ird�v�slp���x�hex��v�re8?�Ɵx�key�v�cpm��x�us$�6�gcr��F�����8�[�q27j92�v��ollismqSk��9O�ݝ� (pl�.���t��p!o��2 9$Fo8��cg7no@ƿtptcls` C�LS�o�b�\�km�ai_
�s>�v�o	��t�b���ӿ�E�H��6�1enu5�01�[m��uti|a|$calmaUR���CalMateNT;R51%�i=1]@ -��/V� ��Z�� �tfq1�9 "K9E��L����2m�CLcMTq�S#��et ��LM3!} �F�c��nspQ�c���c�_moq��� ��c1_e�����su��ޏ� �_ �@�5�G�join�i�j��oX��ł&cWv	 ���N�v9e��C�clm�&A�o# �|$finde��0STD �ter FiOLANG���R���
��n3��z0Cen���r,������ J����� ���K�〪Ú�=���_Ӛ��r~� "FNDR��� 3��f��tguid�䙃N�."��J�tq�� ��������� ����J����_������c��	m�Z��?\fndr.��n#�>
B2p��Z�CP� Ma�����38PA��� c��6� (�� �N�B�������H 2�$�81��m_���"ex�z5� .Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$�r*$ ��*$r*$%/s#C�d/�.,P�/0*ʲD�PN��$���$*�G}r�$k Exc�'{IF�$MASK�%�93 H5�%H5�58�$548 H��$4-1�$��#1(�$�0 E�$��$-b��$���!UPDT ��B�4�b�4�2�49�0`�4a�3�9j0"M�4<9�4  ��4��4tpsh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4���3adq\�5K�979":E�ajO l "DQ^E^�3�i�Dq ��4ҲO ?R�? ��q�5��T���3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F��t�4��.�5y N� >�2il(in�4��31 JH1�2Q4�2�51ݠ�4rmal� �3)�REo�Z_�� �Ox����4��^F�?onorTf��7_ja�UpZҒ4l�5rmsAU��Kkg���4�$HCd\��fͲ�eڱ�4�REM����4yݱ"u@�RERG5932fO��47Z�>�5lity,�U��8e"Dil\�5�r�o ��7987�?8�25 �3hk910�3 ��FE�0=0P_�Hl\mhm�5� �qe�=$�^�
E��u<�IAymptm�U��BU��vste�y\� 3��me�b�DvI�[�Qu �:F�Ub�*_�
E&,�su��_ E�r��ox���4hu#se�E-�?�sn��������FE��,�box�����c݌,"��� ����z��M��g��pdspw)�	�� 9���b���(��1���c��Y�R��  �>�P���W��������'�0ɵ�[���͂���  �w ,�@� �zA�bumpšuf��B*�Box%��7Aǰ60�BBw���MC� (6�,f�t{ I�s� ST���*��}B�����w��"BBF
�>�`����)��\bbk968 "�4��։�bb�9va69�����etbŠ��X�����ed	�F��1u�f� �sea"������'�\��,���b�ѽ�o6�H�
�	x�$�f���!y����Q[�! tpermr�fd� TPl0~o� Recov,���3D��R642� � 0��C@}s� tN@��(U�rro����yu2r��  ?�
  �����$$CLe� O�������������$z�_DIGsIT��������.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$j����+c:PRODU�CTM�0\PGSTKD��V&ohozf�99��D����$FEAT_I�NDEX��xd���  
��`ILECOMPW ;���#��`��cSETUP2� <�e�b��  N �a�c_�AP2BCK 1�=�i  �)�wh0?{%&c�� ��Q�xe%�I� m���8��\�n� ���!���ȏW��{� �"���F�Տj���w� ��/�ğS������� ��B�T��x������ =�үa������,��� P�߯t������9�ο �o�ϓ�(�:�ɿ^� ��Ϗϸ�G���k�  �ߡ�6���Z�l��� ��ߴ���U���y�� ���D���h��ߌ�� -���Q��������� @�R���v����)��� ��_�����*��N ��r��7�� m�&�3\�i�
pP 2#p�*.VRc�*��� /���PC/1/FR6:/].��/+T�`�/�/F%�/�,�`xr/?�*.F�D8?	H#&?e<�/<�?;STM �2�?н.K �?�=i�Pendant �Panel�?;H �?@O�7.O�?y?�O:GIF�O�O�5�OoO8�O_:JPG _J_��56_�O_�_�	P�ANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEINS.XML���0\���qC�ustom To�olbar	���PASSWORD�yFRS:\�L�� %Pas�sword Config���֏e� Ϗ�B0���T�f��� �������O��s�� ����>�͟b��[��� '���K��򯁯��� :�L�ۯp�����#�5� ʿY��}��$ϳ�H� ׿l�~�Ϣ�1����� g��ϋ� ߯���V��� z�	�s߰�?���c��� 
��.��R�d��߈� ��;�M���q���� ��<���`������%� ��I��������8 ����n���!�� W�{"�F� j|�/�Se ��/�/T/�x/ /�/�/=/�/a/�/? �/,?�/P?�/�/�?? �?9?�?�?o?O�?(O :O�?^O�?�O�O#O�O GO�OkO}O_�O6_�O /_l_�O�__�_�_U_ �_y_o o�_Do�_ho �_	o�o-o�oQo�o�o �o�o@R�ov ��;�_��� *��N��G������ 7�̏ޏm����&�8� Ǐ\�돀��!���E� ڟi�ӟ���4�ßX� j��������įS���w������B�#��$�FILE_DGB�CK 1=���/���� ( �)
SU�MMARY.DG<L���MD:������Diag Summary���Ϊ
CONSLO�G�������D�ӱ�Console �logE�ͫ��MEMCHECK:��!ϯ���X�Mem�ory Data|��ѧ�{)��HADOW�ϣϵ��J���Shado�w Change�sM�'�-��)	FTP7Ϥ�3ߨ����Z�mment� TBD��ѧ0=�4)ETHERNET�������T��ӱEthern�et \�figu?rationU�ؠ~��DCSVRF��p�߽�����%��� verify �all��'�1PY=���DIFF�����[���%��d�iff]������1pR�9�K��� ����X��CHGAD������c��r����2ZAS�� ��GD ���k��z��FY3bI[�� �/"GD ���s/����/�*&UPDATE�S.� �/��FR�S:\�/�-ԱU�pdates L�ist�/��PSRBWLD.CM(?����"<?�/Y�PS�_ROBOWEL ��̯�?�?��?&�O -O�?QO�?uOOnO�O :O�O^O�O_�O)_�O M___�O�__�_�_H_ �_l_o�_�_7o�_[o �_lo�o o�oDo�o�o zo�o3E�oi�o ���R�v� ��A��e�w���� *���я`�������� �O�ޏs������8� ͟\�����'���K� ]�쟁����4���ۯ j������5�įY�� }������B�׿�x� Ϝ�1���*�g����� Ϝ���P���t�	�� ��?���c�u�ߙ�(� ��L߶��߂���(� M���q� ���6��� Z������%���I��� B�����2�����h�����$FILE�_� PR� ���������MDONLY� 1=.�� 
 ���q����� �����~%� I�m�2� �h��!/�./W/ �{/
/�/�/@/�/d/ �/?�//?�/S?e?�/ �??�?<?�?�?r?O �?+O=O�?aO�?�O�O &O�OJO�O�O�O_�O�9_�OF_o_
VIS�BCKL6[*�.VDv_�_.PF�R:\�_�^.P�Vision V?D file�_�O 4oFo\_joT_�oo�o �oSo�owo�oB �of�o�+�� �����+�P�� t������9�Ώ]�� ����(���L�^���� ���5���ܟk� ��� $�6�şZ��~������
MR_GRPw 1>.L���C4  B���	� W������*u���R�HB ��2 ���� ��� ���B�����Z�l��� C���D�������Ŀ���I�?�L���]J�h�F�5�UT	zQ�񌲿�ֿ Gk�W�E��ED��+-���:���@<W^�@��A��_f��?m�A����r��E�� F�@ �������J���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6�\b��B��<%���A�o=�@�0eߋ�NҞ�A��߲� v���r������
�C� .�@�y�d������ ��������?�Z�l�v��BH�� ��R�@(h�E��������
0�PJ��P��V"��ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�OPгߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������>[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U��0
//./A�#��� �~/����/�/�/ �/� ?2?D?V?h?�/ ?�?�?�?�?�?�?� ��@O?dO�/�O�O �O�O�?�O�O__*_ MON_�Or_�_�_�_�_ 	OO-O�_A_&ouOJo \ono�o�o=o�o�o�o �oo�o4FXj |�_�_�_o�7o ��0�B�T�#x��� �������e����� ,�>�����ŏ�� �Ο������:� L�^�p�����'���ʯ ܯ� �O�a�s����� l���������ƿؿ�� ��� �2�D�g��z� �Ϟϰ����#�5�G� I��}�R�d�v߈ߚ� iϾ��������)߫��<�N�`�r��XST_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������O�C�R.RDzVT=#��K@9�BOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ�{
�Å��ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A���   @�<�P�R�
h�BD�b�A��j�����������Dz۩���������j��(� �� -���C���'�7�������Y����� �??�ff ��g|y ������q:a��
>+�  PƱj�(�����7	���|�?˙���xZ�p<
�6b<߈;����<�ê<�? <�&Jσ��AI�ɳ+���?offf?I�?&��k�@�.��J<?�`�q�.� �˴fɺ�/��5/� ���j/U/�/y/�/�/ �/�/�/?�/0?q��F�?l??�?/�?+)�?�?�E��� E�I�G+� F��?)O�?9O_O`JO�OnO�Of�BL޳B�?_h�.��O�O�� %_�OL_�?m_�?�__�_�_�_�_�
�h�yÎg>��_�Co�_goRodo�o�GA�ds�q�C�o�o�o|����$]�Hq���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?��$�?�K�0���
=ç>�����3�W
=�s#�W��e�צ��@����{�����<���(�B�u���=B0�������	L��H��F�G���G���H�U`E����C�+���I�#�I��H�D�F��E��RC�j=���
I��@H��!H�( E?<YD0q� $��H�3�l�W���{� �������՟���2� �V�A�z���w����� ԯ��������R� =�v�a���������� ��߿��<�'�`�K� ��oρϺϥ������ ��&��J�\�G߀�k� �ߏ��߳�������"� �F�1�j�U��y�� ����������0���T�?�Q����(�1�3�3/E�����5�������M3ǭ8�����M4M�gs&IB+�2D�a���{�^^	����(��uP2P7Q4_A��M0bt��R�����,�/   �/� b/P/�/t/�/ *a)_ 3/�/�/�%1a?��/?;?M?_?q?  �?�/�?�?�?�?O~ 2 F�$�v'Gb�/�A��@�a,�`�qC��C@�o�O�2���OF� D�zH@�� F�P D���O�O�ys<O!_3_E_W_i_s�?���@@pZJ.t22!2~
 p_�_�_ �_	oo-o?oQocouo��o�o�o�o��Q ���+��1��$�MSKCFMAP�  �5� �6�Q�Q"~�c�ONREL  �
q3�bEX_CFENB?w
s�1uXqFNC_QtJOGOVLIM?w�dIpMrd�bKEY�?w�u�bRUN�|�u�bSFSPDTY�avJu3s�SIGN?QtT1�MOT�Nq�b_�CE_GRP 1-p�5s\r��� j�����T��⏙�� ����<��`��U��� M���̟��🧟�&� ݟJ��C���7����� ��گ�������4�V��`TCOM_CF/G 1q}�Vp�􂿔�
P�_ARC�_\r
jyUAP�_CPL��ntNO�CHECK ?{ 	r� �1�C�U�g�yϋϝ� ����������	��({�NO_WAIT_�L�	uM�NTX��r{�[m�_ER�RY�2sy3� A&�������r�cx� ��T_MO��}t��,  �I$�|k�3�PARAM��u{��V[���!�u?�� =9@345678901� �&���E�W�3�c������{������� �����=�UM_?RSPACE �V�v��$ODRD�SP���jxOFF�SET_CART�ܿ�DIS��PEN_FILE� �q��c֮�OPTI�ON_IO��PWORK v_�ms �P(�R��@�6$j.j	 ��Hj(6$�p=��_DSBL  Ċ5Js�\��RI_ENTTO>p9!sC��Pq=#��UT_SIM_D�
r�b� V� LCT ww�bc���U)+$_PEXE�d&RATp �vju��p��2X�j)TU�X)TX�##X d-�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O?O�H2�/oO�O�O�O��O�O�O�O�O_]�< ^O;_M___q_�_�_�_ �_�_�_�_o���X��OU[�o(�꘯(���$o��, ��IpB` �@D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	l�mb�`�xJ�`�����a�< ��`��m�a, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�b���� �N U�B[�'!o�:q�pC\�C�@@sBq�|���= m�
�A\��h@ߐ�n����Z��B\��A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�����(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��� ��3 ���Ӱ��ɆDT� Qy-����D � ��ӱ4�P :� L :�GP:�D :�@ :�U8�8�	8�
8�U8�8�8�8�Q8�X@:�8�8�8�8�8��:�E8�8�x�:�8�PP�:�d :�8�8�P��:�
�:�!8�"8�Q#8���:�%8�&8�U'8�(8�)8�*8�T��:�,8�-8�.8�/8�08�18�,��� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�X�(�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_d��_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п�_��� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p�������� //$)�$�PGTRACEL�EN  #!  ��" ��8&_UP z/���g!o S!�h 8!_CFG7 {g%Q#"!�x!�$J �#|"DEFSPD |�,�!!J �8 IN~ TRL }�-�" 8�%�!PE__CONFI� ~g%��g!�$\�%�$LID�#�-�74GRP 1��7Q!�#!A ����&ff"!A�+33D�� D�]� CÀ A)@+6�!�" d�$�9��9*1*0� 	 �+9�(�&�"�? ��	C�?�;B@3AO��?OIO3OmO"!>�?T?�
5�O�O��N�O =��=#�
�O_�O_J_ 5_n_Y_�O}_�_y_�_<�_�_  Dzco" 
oBo�_Roxoco �o�o�o�o�o�o�o�>)bM��;�
V7.10be�ta1�$  �A�E�rӻ�A " �p?!G���q>���r�܁0�q�ͻqBQ��qA\�p�q�4T�q�p�"�BȔ 2�D�V�h�w��p�?�?)2{ȏw�׏ ���4��1�j�U��� y�����֟������ 0��T�?�x�c����� ��ү����!o�,�ۯ P�;�M���q�����ο ���ݿ�(��L�7��p�+9��sF@  �ɣͷϥ�g%����� �+�!6I�[߆����� �ߵߠ���������!� �E�0�B�{�f��� ����������A� ,�e�P���t������� �����=(a L^������ �'9$]�Ϛ� �ϖ�������/ <�5/`�r߄ߖߏ/> �/�/�/�/�/?�/1? ?U?@?R?�?v?�?�? �?�?�?�?O-OOQO <OuO`O�O�O�O�O�� �O_�O)__M_8_q_ \_n_�_�_�_�_�_�_ o�_7oIot���o �o���o�o�o(/! L/^/p/�/{*o�� �������A� ,�e�P�b��������� �Ώ��+�=�(�a� L���p������Oߟ� ��� �9�$�]�H��� l�~�����ۯƯ��� #�No`oro�on��o�o �o�oԿ���8J \ng����vϯϚ� ������	���-��Q� <�u�`�r߫ߖ��ߺ� ������;�M�8�q� \��������z���� ��%��I�4�m�X��� |�����������:� L�^���Z������� ����$�6�H� Swb���� ���//=/(/a/ L/�/p/�/�/�/�/�/ ?�/'??K?]?H?�? ��?�?f?�?�?�?O �?5O OYODO}OhO�O �O�O�O�O�O&8J 4_F_����_�_� �_�_"4-o�O*o coNo�oro�o�o�o�o �o�o)M8q \������� ��7�"�[�m��?�� ��R�Ǐ���֏�!� �E�0�i�T���x��� �����_$_V_ �2��l_~_�_�����R�$�PLID_KNO�W_M  �T������SoV ��U͠�U��
�� .�ǟR�=�O�����m�ӣM_GRP 1���!`0u��T@Rٰo�ҵ�
�� �Pзj��`���!� J�_�W�i�{ύϟϱ����������߱�MR������T��s�w� s��ߠ޴߯߅��� �߻�����A���'� ���������� ����=���#����������}������S��S�T��1 1��U�# ���0�_ A .��,>Pb� �������3 (iL^p��P���2*N���<-/3/)/;/M/4f/x/�/�/5�/�/�/�/A6??(?:?7S?e?w?�?8�?�?�?��?MAD  �d#`PAR�NUM  �w�%OSCH?J �ME
�G`A�Iͣ�EUPD`OrE
a�OT_CMP_��B@�P�@'˥TER_wCHK'U��˪?R$_6[RSl�¯��G_MOA@�_�U_�_~RE_RES_G ��>�oo8o+o \oOo�oso�o�o�o�o��o�o�o�W �\ �_%�Ue Baf�S � ����S0�� ��SR0��#��S�0 >�]�b��S�0}������RV 1�����rB�@c]��t�(�@c\����D�@c[�$���RT?HR_INRl�DA���˥d,�MASS69� ZM�MN8�k��MON_QUEUE ���˦��x�� RDNPUbQN8{�P[��END���_�ڙEXE�ڕ�@B�E�ʟ��OPTI�OǗ�[��PROG�RAM %��%���ۏ�O��TAS�K_IAD0�OCFG ���tO��Š�DATA���Ϋ@��27�>�P�b� t���,�����ɿۿ������#�5�G���IN+FOUӌ������ �ϭϿ��������� +�=�O�a�s߅ߗߩ߀���������^�jč�� yġ?PDI�T �ίc���W�ERFL
��
RGADJ �n�A����?����@�~��IORITY{��QV���MPDSP(H�����Uz����oOTOEy�1�R� (!AF4��E�P]���!t�cph���!u�d��!icm���ݏ6�XY_ȡ�R��ۡ)� a*+/ ۠� W:F�j��� ���%7[�B�*��POR�T#�BC۠�����_CARTRE�P
�R� SKSTyAz��ZSSAV����n�	2500H863���r�$�!�R�����q�n�}/�/�'� UR�GE�B��rYWFF� DO{�rUVWV���$�A�WRUP_�DELAY �|R��$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?�3AQSKIP!�vn�l#x 	1/ +O+ OROdOvO9Hn� �O�G�O�O�O�O�O_ �O_D_V_h_._�_z_ �_�_�_�_�_
o�_.o @oRoovodo�o�o�o �o�o�o�o*<�Lr`���n��?$RCVTM������pDCR!��LЈqC`N��C�d�C��o�?��>��L�<|�{4M�g��&��/����%�t����|��}'�4Oi��O� <
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E0�kATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960�iW+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�M)�$bR  ��ϰ�P{_�P_INTVAL�@�����JR_OPT�ION�V �E�BpVAT_GRPw 2����G(y_Ho �e_ vo�o�oYo�o�o�o�o �o*<�bOoND pw������ 	���?�Q�c�u��� ��/���ϏᏣ���� )�;���_�q������� ��O�ɟ���՟7� I�[�m�/�������ǯ ٯ믁��!�3���C� i�{���O���ÿտ� ��ϡ�/�A�S�e�'� �ϛϭ�oρ������ �+�=���a�s߅�G� �߻����ߡ���'� 9�K�]��߁���� y����������5�G��Y��E�$SCAN�_TIM�AYue�w�R �(�#�((�<0.aWaPaP
T�q>��Q��o������OO"2/���d;2"BaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>HE�̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:L!`O�UT",REC 1�Z� d �  	  	������

 �Z�{0 H6lZ�~�� ���� //D/2/ h/z/\/�/�/�/�/�/ �/�/?�/,?R?@?v? d?�?�?�?�?�?�?�? OO(ONO<OrOTOfO �O�O�O�O�O�O_&_ _J_8_Z_\_n_�_�_ �_�_�_�_�_"ooFo 4oVo|o^o�o�o�o�o �o�o�o0TB xf����(� ��,��P�>�`��� h���������Ώ�� (�:��^�L���p��� ����ܟ���� �6� $�Z�H�~���r����� دƯ����2��&� h�V���z�����Կ� ȿ
�����.�d�R� �Ϛ�|ϾϬ������ ���<��`�N�pߖ� �ߺߨ���������8�&�\�J�l��jV� 1�w Pl��	>� � ��&��
TYPE�VFZN_CF�G �x��d7�GRP� 1�A�c ,�B� A� D;�� B���  B�4RB21^HELL:�(
 X����%RSR���� E0iT�x�� ����/S�ew�����%@w�����#�1����A��2#�d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he�s_ (_:_L_^_��_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}4xcopy �fr:\*.* �virt:\tm�pback�Q=>�192.168.�4�P46:216�4 �R�_�_�_�K}5�Ua�_�_�V�_go�yo�o}9�Ts:o�rderfil.dat.l@oVo�o�o�}0�Rmdb: +o�oRb�ocu�b �_2o?U��
�o ��Sod�v����o�o 6Q���+Ə O`�r����*�<�� ޟ���'���K�\��n����
xyzrate 61 +�@=�O�������>��1356 ��ү c�u�������5�6�ٿ ����"���5�ѿb��tφ��6����em}p:�6088 W�����ύ�.��*.d�������`�r߄ߗ�1 +�=�O������� )�������c�u� ��5����������"� ������b�t������� ��:�V����������8 ��gy��� ��9�T���	�� @��cu���-? ����/��N _/q/�/�ߨ�:/L/�/��/?( �ǖ792 �/�/b?t?�?#8��*?<0�?�?�?-/ �?39�?aOsO��O�Ϫ?��̑534 Ӑ�O�O�O� ߺO�H �O`_r_�_�/��;_M_ �_�_o�'?�T�_�_ couo�o��?5O�G�o �o�o"O�o�H�ob t���/�/QcU� �
�/��T`�g� y����o�o9T��� 	���@ҏc�u�������$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1����?���% ֟��&�	��\�?� f���u��������ϯ ��"��F�)�;�|�_� ������ֿ��˿�� �B�%�f�I�[Ϝ�� ���ϵ�������,�� 6�b�E߆�i�{߼ߟ� ����������L�/� V��e������� �����6��+�l�O� v��������������� 2V9K�o ������� &R5vYk�� ���/��<// F/r/U/�/y/�/�/�/ �/?�/&?	??\??? f?�?u?�?�?�?�?�? �?"OOFO)O;O|O_O �O�O�O�O�O�O_�O _B_%_f_I_[_�__ �_�_�_�_�_�_,oo 6oboEo�oio{o�o�o �o�o�o�oL/ V�e����� ���6��+�l�O��v�������PARAoM �����_ �	��P�����OFT_�KB_CFG  �ヱ���PIN_�SIM  ����C�U�g�����RV�QSTP_DSB�,�򂣟����SR� �/�� & �MULTIROBOTTASK������TOP_�ON_ERR  ����PTN� /�@��A	�RING_�PRM� ��V�DT_GRP 1y�ˉ�  	�� ����������Я��� ��*�Q�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߣߠ߲��� ��������0�B�i� f�x���������� ���/�,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZ�~��� ����/ /G/D/ V/h/z/�/�/�/�/�/ �/?
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8___\_��VPRG_COUNT���@���RENB�U��UM�S��__U�PD 1�/�8  
s_�oo*o SoNo`oro�o�o�o�o �o�o�o+&8J sn������ ���"�K�F�X�j� ��������ۏ֏��� #��0�B�k�f�x��� ������ҟ������ C�>�P�b����������ӯί�����UY?SDEBUG�P�P��)�d�YH�SP_�PASS�UB?~Z�LOG ��U+�S)�#�0��  ��Q)�
M�C:\��6���_M�PC���U���Q�ñ8� �Q�SAV �����ǲ&��ηSV;�TE�M_TIME 1���[ (  �w�"����$T1?SVGUNS�P�U�'�U���ASK_OPTION�P��U�Q�Q��BCC�FG ��[u� qn�A�a�`a� gZo��߃ߕ��߹��� ����:�%�^�p�[� ��������� ��� ��6�!�Z�E�~�i���������&������� &8��nY�} �?��ԫ �� (L:p^�� �����/ /6/ $/F/l/Z/�/~/�/�/ �/�/�/�/�/2?8  F?X?v?�?�??�?�? �?�?�?O*O<O
O`O NO�OrO�O�O�O�O�O _�O&__J_8_n_\_ ~_�_�_�_�_�_�_o �_ o"o4ojoXo�oD? �o�o�o�o�oxo .TBx��j� �������,� b�P���t�����Ώ�� ޏ��(��L�:�p� ^�������ʟ��o ��6�H�Z�؟~�l� ������د���ʯ � �D�2�h�V�x�z��� ¿���Կ
���.�� >�d�Rψ�vϬϚ��� ��������*��N�� f�xߖߨߺ�8����� ����8�J�\�*�� n������������ "��F�4�j�X���|� ������������0 @BT�x�d� ����>, Ntb����� �/�(//8/:/L/ �/p/�/�/�/�/�/�/ �/$??H?6?l?Z?�? ~?�?�?�?�?�?O� &O8OVOhOzO�?�O�O �O�O�O�O
__�O@_ ._d_R_�_v_�_�_�_ �_�_o�_*ooNo<o ^o�oro�o�o�o�o�o �o J8n$O �����X����4�"�X�B�v��$�TBCSG_GR�P 2�B���  �v� 
 ?�  �� ����׏�������1���U�g�z���ƈ�_d, ���?v��	 HC��d�>�����e�CL � B���Пܘ������\)��Y�  A�ܟ$�B��g�B�Bl�i�X�������X��  D	 J���r�����C���H��үܬ���D�@v� =�W�j�}�H�Z���ſ@��������v��	V3.00~��	m61c�	*X�P�u�g�pœ>���v�(:�� q��p͟�  O�����p�����z�J�CFG �B�e�� �����������=�� =�c�q�K�qߗ߂߻� ���������'��$� ]�H��l������ ������#��G�2�k� V���z����������� ���p*<N�� �l������ �#5GY}h ����v�b��>� // /V/D/z/h/�/ �/�/�/�/�/�/?
? @?.?d?R?t?v?�?�? �?�?�?O�?*OO:O `ONO�OrO�O�O��O �O�O_&__J_8_n_ \_�_�_�_�_�_�_�_ �_�_oFo4ojo|o�o �oZo�o�o�o�o�o�o B0fT�x� ������,�� P�>�`�b�t�����Ώ �������&�L��O d�v���2�����ȟʟ ܟ� �6�$�Z�l�~� ��N�����دƯ��  �2��B�h�V���z� ����Կ¿����.� �R�@�v�dϚψϪ� �Ͼ�������<�*� L�N�`ߖ߄ߺߨ��� �ߚ�������\�J� ��n��������� �"���2�X�F�|�j� �������������� .TBxf�� �����> ,bP�t��� ��/�(//8/:/ L/�/�ߚ/�/�/h/�/ �/�/$??H?6?l?Z? �?�?�?�?�?�?�?O �?ODOVOhO"O4O�O �O�O�O�O�O
_�O_ @_._d_R_�_v_�_�_ �_�_�_o�_*ooNo <oro`o�o�o�o�o�o �o�o&�/>P�/ ������� ��4�F�X��(��� |�����֏����Ə 0��@�B�T���x��� ��ҟ������,�� P�>�t�b��������� ������:�(�^� L�n�������2d� ����̿�$�Z�H�~� lϢϐ��������Ϻ�  ��0�2�D�zߌߞ� ��j����������
� ,�.�@�v�d���� ����������<�*� `�N���r��������� ����&J\� t��B���� ��F4j|� �^����/��  2 6# �6&J/6"�$TBJ�OP_GRP 2���� � ?�X,i#��p,� �_xJ� �6$��  �< ��� �6$ @�2 �"	 �C��} �&b  Cق'<�!�!>���
55�9>�0+1�33�=�CL� f�ff?+0?�ff�B� J1�%Y?d7�.���/>��2\�)?0�5���;���hCY� � � @� �!B�  �A�P?�?�3EC�  D�!�,�0*B�Oߦ?�3JB��
:���Bl�0���0�$�1�?O6!A�ə�AДC�1D9�G6�=q�E6O�0�p��B�Q�;�A�� �o��@L3D	�@��@__�O�O>B��\JU�OHH�1ts>�A@33@?1� C�� �@�_�_&_8_�>��D�UV_0�xLP�Q30<{�zR� @�0�V�P!o3o�_ <oRifoPo^o�o�o�o Ro�o�o�o�oM( �ol�p~��p4�6&�q5	V�3.00�#m61c�$*(��$1!�6�A� Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,IR�CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;S@�;Q��|8�`�rz@/&�8�6&�<��1�w�^$ESTPARS  *(�{ _#HR��ABL/E 1�p+Z�6#�|�Q� � 1�|�B|�|�5'=!|�	|�E
|�|�˕6!|��|�|���RD	I��z!ʟܟ� ��$���O������¯�ԯ�����S��x#  V���˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������U-���� ĜP�9�K�]�o��-��?�Q�c�u���6�NUoM  �z!� >  Ȑ����_CFG ������!@b IMEBF_TT����x#���a�VER��b�w��a�R 1�p+
 �(3�6"1 ��   6!���������� � 9�$�:�H�Z�l�~��� ������������^$R��_��@x�
b MI_CHANm�� x� kDBGL�V;0o�x�a!n E�THERAD ?U�� �y�$�"�\&n ROUT6��!p*!*~�SNMASK�|x#�255.h��fx^$OOLO_FS_DI��[���	ORQCTRL �p+;/��� /+/=/O/a/s/�/�/ �/�/�/��/�/�/!?���PE_DETA�I��PON_S�VOFF�33P_?MON �H�v��2-9STRTCH/K ���42�VTCOMPAT�a8�24:0FPRO�G %�%M�ULTIROBO�TTO!O06�PL�AY��L:_INSWT_MP GL7�YDUS���?�2LC�K�LPKQUICK�MEt �O�2SCR�E�@�
tps��2�A�@�I���@_Y���9�	SR_GRP 1��_ ���\� l_zZg_�_�_�_�_�_�^�^�oj�Q'ODo /ohoSe��oo�o�o �o�o�o�o!W E{i�������	12345C67��!���X�E�1�V[
 �}�ipnl/a�gen.htmno����𤏶�ȏ~�Pa�nel setup̌}�?��0�B�T�f� ��񏞟�� ԟ���o����@� R�d�v������#�Я �����*���ϯů r���������̿C�� g��&�8�J�\�n�� ���϶���������u� �ϙ�F�X�j�|ߎߠ� ���;�������0��B��*NUALRM�b@G ?��  [������������  ��%�C�I�z�m��������v�SEV  �����t�ECFG Ձ=]/B�aA$   B�/D
 ��/C�W i{�������� PRց;� �To\o�I�6?K0(%����0� ����//;/&/ L/q/\/�/�/�/l�Dc �Q�/I_�@HIST 1ׁ9�  (  ���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1 Ec0p?�?8�?�?/C�� >?P=962n?�?
OO.O�?�?�136c?|O�O �O�OAOSO�?�O__ 0_�O�O_Lu_�_�_�_ :_�/�_�_oo)o;o �__oqo�o�o�o�oHo��o�o%7I~� �a81�ou���� ��o���)�;�M� �q���������ˏZ� l���%�7�I�[�� �������ǟٟh��� �!�3�E�W������ ����ïկ�v��� /�A�S�e�Pb���� ��ѿ������+�=� O�a�s�ϗϩϻ��� ����ߒ�'�9�K�]� o߁�ߥ߷������� �ߎ�#�5�G�Y�k�}� ������������� ��1�C�U�g�y���v� ����������	� ?Qcu��(� ���)�M _q���6�� �//%/�I/[/m/ /�/�/�/D/�/�/�/ ?!?3?�/W?i?{?�? �?�?�����?�?OO /OAOD?eOwO�O�O�O �ONO`O�O__+_=_ O_�Os_�_�_�_�_�_ \_�_oo'o9oKo�_ �_�o�o�o�o�o�ojo �o#5GY�o}�������?���$UI_PANE�DATA 1������?  	�}�0�`B�T�f�x��� )�� ��mt�ۏ����#� 5���Y�@�}���v��� ��ן�������1���U�g�N������ �1��Ïȯگ��� �"�u�F���X�|��� ����Ŀֿ=����� �0�T�;�x�_ϜϮ� ���Ϲ������,ߟ�M��j�o߁ߓߥ� �������`��#�5� G�Y�k��ߏ����� ����������C�*� g�y�`���������F� X�	-?Qc�� ��߫���� ~;"_F�� |�����/� 7/I/0/m/�����/�/ �/�/�/�/P/!?3?� W?i?{?�?�?�??�? �?�?O�?/OOSOeO LO�OpO�O�O�O�O�O _z/�/J?O_a_s_�_ �_�_�O�_@?�_oo 'o9oKo�_oo�oho�o �o�o�o�o�o�o#
 GY@}d��&_ 8_����1�C�� g��_��������ӏ� ��^���?�&�c�u� \�������ϟ���ڟ �)��M������� ����˯ݯ0����� 7�I�[�m�������� ��ٿ�ҿ���3�E� ,�i�Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#� ������ ��$�6�� Z�A�~�e�w����� �������2��V�h��O�����v�p��$U�I_PANELI�NK 1�v��  � � ��}1234567890�� ��	-?G ��� o�����a���#5G�	��h��p&���  R �����Z�� $/6/H/Z/l/~//�/ �/�/�/�/�/�/
?2? D?V?h?z??$?�?�? �?�?�?
O�?.O@ORO dOvO�O O�O�O�O�O �O_�O�O<_N_`_r_�_�_�0,���_�X �_�_�_ o2ooVoho Ko�ooo�o�o�o�o�o �o��,>r}�� �������� ��/�A�S�e�w�� ������я���tv� z����=�O�a�s� ������0S��ӟ��� 	��-���Q�c�u��� ����:�ϯ���� )���M�_�q������� ��H�ݿ���%�7� ƿ[�m�ϑϣϵ�D� �������!�3�Eߴ_ i�{�
�߂����߸� �����/��S�e�H� ���~��R~'�'�a ��:�L�^�p����� ���������� �� 6HZl~��� #�5��� 2D ��hz����� c�
//./@/R/� v/�/�/�/�/�/_/�/ ??*?<?N?`?�/�? �?�?�?�?�?m?OO &O8OJO\O�?�O�O�O �O�O�O�O[�_��4_ F_)_j_|___�_�_�_ �_�_�_o�_0ooTo fo��o��o��o�o �o,>1bt ����K��� �(�:����{O�� ����ʏ܏�uO�$� 6�H�Z�l��������� Ɵ؟����� �2�D� V�h�z�	�����¯ԯ ������.�@�R�d� v��������п��� ϕ�*�<�N�`�rτ� �O�Ϻ�Io������� ��8�J�-�n߀�cߤ� �����߽����o1� �oX��o|������ �������0�B�T� f�������������� S�e�w�,>Pbt ��'���� �:L^p�� #���� //$/ �H/Z/l/~/�/�/1/ �/�/�/�/? ?�/D? V?h?z?�?�?�???�? �?�?
OO.O��ROdO �߈OkO�O�O�O�O�O �O_�O<_N_1_r_�_�g_�_7OM�m��$UI_QUICKMEN  ��_Aob�RESTORE �1�  �|��Rto�o�im�o�o�o�o �o:L^p�% ������o�� ��Z�l�~�����E� Ə؏���� �ÏD� V�h�z���7������� /���
��.�@��d� v�������O�Я��� ��ßͯ7�I���m� ������̿޿���� &�8�J��nπϒϤ� ��a�������Y�"�4� F�X�j�ߎߠ߲��� ���ߋ���0�B�T��gSCRE`?�#mu1sc�o`u2��3��4���5��6��7��8<��bUSERq�v�2��Tp���ks����U4��5��6��7���8��`NDO_C�FG �#k  �n` `PDAT�E ����NonebSEU�FRAME  �TA�n�RTOL_ABRTy�l���ENB����GRP� 1�ci/aCz  A�����Q��  $6HRd���`U�����MS�K  �����N&v�%�U�%����bVISCAND�_MAX�I����FAIL_ISMG� �PݗP#���IMREGNU�M�
,[SIZl�n`�A�,V?ONTMOU���@���2��a��a����FR:\ �� MC:�\�\LOG�B@F� !�'/!�+/O/�Uz �MCV�8#UDM1r&EX{+�S�P>PO64_��0�'fn6PO���LIb�*�#V����,f@�'�/�w =	�(SZV�.w����'WAI�/�STAT ߄���P@/�?�?�:$�?�?��2DWP�  ��P G<@+b=��� H��O_JMPER�R 1�#k
  ��2345678901dF�ψO{O�O �O�O�O�O_�O*__�N_A_S_�_
� ML�OWc>
 �_T�I�=�'MPHASE  ���F��PSHIF�T�1 9�]@<�\�Do�U#oIo�o Yoko�o�o�o�o�o�o �o6lCU� y����� ���	�V�-�e2����	�VSFT1�2	�VM�� �5ԑ1G� ���%Aȯ  B8̀̀�"@ pكӁ˂�у��Fz�ME@�?�{�\�!c>&%�aM1�i�k�0�{ �$`0TDINEND��\�O� �z�����S��w��P���ϜRELE�Q��Y����\�_ACTI�V��:�R�A ���e���e�:�RD�� ���YBOX c�9�د�6��0�2���19o0.0.�83�;�254��QF�	 �X�j���1�rob�ot���   �p�૿�5pc��̿�����7�𼻲�-�f�ZABC
�����,]@U��2ʿ �eϢωϛϭϿ��� �� ���V�=�z�a�Hs߰�E�Z��1�Ѧ