��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �� �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ڏ1�	 H PC�UREQ1 � $SOFT; �T_ID�TOT�AL_EQ� $� � NO�PS_�SPI_INDE���$�X�SC�REEN_NAM�E �SI�GN��� P�K_FIL	$�THKYMPAN�E�  	$D�UMMY12 �� u3|4|&��ARG_STR�1 � $T�ITP$I��1�{������5�6�7�8
�9�0��z�P����1�1��1 '1
'2"GS�BN_CFG1 � 8 $CN?V_JNT_* |�$DATA_C�MNT�!$FL�AGS�*CHE�CK�!�AT_C�ELLSETUP�  P $HOME_IO,�G�%�#MACR=O�"REPR�(-�DRUN� D|�3SM5H UTO�BACKU0� $ENAB���!EVIC�T]I � D� �DX!2ST� ?0B��#$INTERV�AL!2DISP_�UNIT!20_D�On6ERR�9FR�_F!2IN,G�RES�!0Q_<;3!4C_WA�471^�:OFF_ N�3wDELHLOGn285Aa2?i1@FN?�� -M���W+0�$Y $D�B� 6COMW!2MO� "0G_A.o	 \rVE�1�$F��A{$�O��D�B�CTMP�1_F�E2�G1_��3�B�2�XD��#
 d $�CARD_EXI�ST4$FSS�B_TYPuAH�KBD_S�B�1A�GN Gn $�SLOT_NUM�JQPREV,DB�U� g1� ;1_ED�IT1 � *1G=� S�0�%$EP�$�OP�AEToE_OKRUS�oP_CRQ$;4x�V� 0LACIw�1�RAPk �1x@M}E@$D�V��Q�Pv�A{�B�L� OUzR ,�mA�0�!� B� L�M_O�^eR�"C�AM_;1 x�r$ATTR84NP� ANN�@5�IMG_HEIG�HQ�cWIDTH�4VT� �UU0F�_ASPECQ;$M�0EXP��@�AX�f�CFT X $GR� �� S�!�@B@NF�LI�`t� UIR�E 3dTuGITCH�C�`N� S�d_Ld�`�C�"�`EDlpE� J�4S�0� �z�sa4 hq;G0 �� 
$WARNM�0f�!,P� �s�p�NST� CORN��"a1FLTR�uT�RAT� T�p H0ACCa1���{�ORI
`"S={�RT0_S�B�C�HG,I1 �[ Tp�"3I9�T�Y12�pHK*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6���7��8��94�ACO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0���`�� �v�p��PzPb26����"J��_R��BC�J��3�JVP��tB�S��}Aw��"�@G C�P_*0OFSzR; @� RO_K8����aIT�3��NOM	_�0�1ĥ3W ��T �� $���AxP��K}EX�� �0�g0I01��p�
$TyFa��C$MD3���TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF0�vF�40CPp@�a�2 
P$A`PU8�3N)#�dR�*�AX�!sDETAI�3BUFV�p@�1 |�p۶�pP�IdT� PP[�M�Z�Mg�Ͱj�F[�SIMQSI�"0��A�.����_�Pkx 	Tp|zM��P�B��FACTrbHPE�W7�P1Ӡ��v��M]Cd� �$*1�JB�p<�*1DEC�Hښ�H��a� �� +PNS_EMP��$GP���,P!_��3�p�@Pܤ��TC��|r��0�s�� b�0�� �B���!
����JR� ��SEGF�R��Iv �aR�TrkpN&S,�PVF4|��� &k� Bv�u�cu��aE�� !2���+�MQ��E�SIZ�3����T��P���|��aRSINF� ����kq���������LX�����F�CRCMu�3CClpG�� p���O}���b�1����P���2�V�DxIC��C���r����P��{�� EV �zF_J��F�pNB0�?�������A�! � r�Rx����V�lp�2���aR�t�,�g�R>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!��$SK��2&nQDB�"�"@�;PR8� 
� ����# >�q1M$��$��+�L9�$?�A
�V�%�@?�AR�PC&�_?(ӫPE��'�~?(�� RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@����C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!��DCS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�g �QSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc��@Sp�i�a+ �j�f�_�ΰAPIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�� 6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6Cq�"MSW�U. 8��KEYI��5�TM�1�s�qLoA�vINޱ�D, �/ D��HOST�P!4���<���`<�°<��p<�EM'����Z�� SBL� U}L��0  �	8����DT�0?1 � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0�QS�����#��SAV �����c�S< 9�`��fP$�0E!� YwN_B�#2 0��DI�d�pO|�m��#�$F�R_IC�� �ENC2_Sd3  ��< 3�9���� cgp����B4�"��2�A��ޖ5���`ǻ��@Q@K&D-!�a�A�VER�q����D3SP
���PC_�q���"�|�ܣ�VALMU3�HE�(�M�sIP)���OPPm �TH�*���S" T�/�Fb�;�d����d ������1�6 H(rLL_DUǀ�a�@��k���֠OT�"U�/����"@@NOAUTO70�$}�x�~�R@s��|�C͠��IC� 2p�z�L�� 8H *��L� ���Բ@sv��` � �� ÿ���Xq��cq����q���q��7��8J��9��0���1�U1 �1-�1:�1G�U1T�1a�1n�2|ʩ2��2 �2-�2�:�2G�2T�2a�2*n�3|�3�3� �U3-�3:�3G�3T�U3a�3n�4|�w�8����9 <���z�ΓKI����H硵ƣ�FEq@{@: y,��&a? PF_P?��>�����E�@��̱QQ��;�fp$TP�$�VARI����,�U�P2Q`< W�߃TD��g���`������wZ���BAC�"G= T2����$)�,p+r³�p IFI�� �p�� q M�P"B`�s�l@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� Fa@��j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(�q�#5T�DG���� �%��pFSS� )�?C P(q1�1�`Q_1"811�EC�13D;5D6�GR)A���@�����P�W�ON2EBUG�S�2�&�gϐ_E A ��z?�P�TERM�5�B�9ORIw�0C��9SM_-`���0Dj�:A�9E�9UP���F� -Qϒ�A�P�3�@B$SE�GGJ� EL�UUS]EPNFI��pB�x��1@��4>DC$U9F�P��$���QD�@C���G�0T��ܘ��SNSTj�PA�Tۡg��APTHJ�A�E*�Z%qB\`F� {E��F�q�pARxPY�aSHFT͢qA�A>X_SHOR$�>�J�6 @$GqPE���OVR���aZPI�@P@$U?r *aAY#LO���j�I�"�p�Aؠ��ؠERV� �Qi�[Y)��G�@R��Pi�e�i�R�!P�u�ASYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U���C�%UP���P���WO�R�@M��k0SkMT��G��GR��3�aPA�@��&�5��'�H � j�NA�TOCjA7pP]Pp$OPd�O��(C�%�p�O!��KRE.pR�C�AO�,?��Be5pR�Eru�Ix'QG�e$PWRf) IMdu�RR_$s� �5��B I�z2H8�=�_ADD�RH�H_LENG��B�q�q:�x�R��S�o�J.�SS��SK������ ��-�SqE*�����HSN�[MN1K	�j�05�@r�֣OL��\��WpW�Q�>pACRO �p���@H ����Q�� ��OUPW3�b_">�I��!q�a1���� ����|���������-���:���iIO
X2S=�D�e���p<`���L $��p��!_OFF[r_�P�RM_�rr�H�TTP_�H��M; (�pOBJ�"�p�G�$H�LE�C|��ٰN � 9�.*�AB_�T��
��S�`�S��LV��K�RW"duHITCOmU?BGi�LO�q����d� Fpk��GpSS� ���HW�h�wA��O.��`I�NCPUX2VISIO��!��¢.�á�<�á-� �IOL]N)�P 87�R'�^[p$SL�bd oPUT_��$dp��Pz �� F_�AS2Q/�$L D���D�aQT U�0]PA������PHY`G灱Z�[p4�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp࿷�x��ٶ����UJ��S����N�E�WJOG�G �D{IS�� �KĠL��3T |��AV���`_�CTR!S^�FgLAGf2&�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_H��Dq��N?���V��EE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�B�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S S�n��0I�BUFF�1XY��PT�A$�� �v��f�p��*1�A�rYY��P ������pOS1�2��3���_�0Z �  ��aiE�\*��IDX�dP�R�hrO�+��A&STʠ�R��Yz�<! /Y$EK&CK+����Z&m&�5�0[ L��o�0��]PL� 6pwq�t^����w��7�?_ \ �`�Р瀰�7��#�0C��]{ ��CLDP��>;eTRQLI�jd8.�094FLGz�0�r1R3�DM�R7��LqDR5<4R5ORG.� ��e2(`���V�8.��T8<�4�d^ �q�<4(��-4R5S�`T00m���0DFRCLM�C!D�?�?3I@�� M9IC��d_ d����RQm�q�DSTB	�  �Fg�H�AX;b �H�LE�XCESZr�rBMup�a`��B;d�ѨrB`��`a��F_�A�J��$[�O�H0K��db \��ӂS�$�MB��LIБ}SREQUIR�R>q�\<Á�XDEBU��oAL� MP�c�ba��Ph؃ӂ!BoAND�ф�`�`d�҆�c�cDC1��IN�����`@�(h?Nz�@q��o��4�TPST8� �e�rLOC�RYI�p�EX�fA�px��A�AODAQP�7f X��ON��[rMF�����f)�"I���%�e��T� �FX�@IGG� g �q��"E�0��#���$R�a%;#7y���Gx��VvCPi�DAT	Aw�pE:�y��RF����NVh t W$MD�qIё)�v+�tń�tH�`�P�ux�|��sANSW}�P�t�?�uD�)�r��	@Ði �@C�U��V�T0�AoAR;R2�j Dɐ�Q�ނ�Bd$CALI��@F�G�s�2�R�IN��v�<� INTE���kE���,�XV�����_Nl���ڂ��kDׄRm�DIViFDH�@ـn�$V��'c!;$��$Z������~�[��o�H �$BELT|b��!ACCEL+q��ҡ��IRC��t����T/!��$SPS�@#2LPqЀƔ83������� ��P�ATH��������3̒Vp�A_�Q�.�4��B�Cᐈ�_MGh�$DDQ���G�$FW���p��m�؝���b�DE��PP�ABNԗROTS�PEED����00J��Я8��@��P$OUSE_��P��Fs�SY��c�A >q�YNu@Ag��OF�F�q�MOUN�N�Gg�K�OL�H�INC*��a��q��Bj�<L@�BENCS��q`�Bđ���D��IN#"�I̒��4�\BݠVE�O�w�Ͳ23_UP�E�߳LOWL ���00����D���B wP��� �1RCʀƶ�MOSIV�JRMO����@GPERCH  �OV��^� �i�<!�ZD<!�c�� d@�P��V1�#P͑��L���EW��ĸ�UP������TR�Kr�"AYLOA 'a�� Q-�̒<�1Ӣ`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H����b��DUM2(�S_BCKLSH_C̒ ��>�=�q�#�U��ԑ����2�t�]ACLAL�vŲ�1n�P�CH�K00'%SD�RTY@4�k��y�1�q_6#N2�_UM$Pj�Cw��_�SCL��ƠLM?T_J1_LO��@���q��E�����p�๕�幘SPC��07������PCo���!H� �PU�m�C/@�"sXT_�c�CN_��1N��e���SFu���V�&#����9�̒��2=�C�u�SH6#�� c����1�Ѩ�o�0�͑�
��_�PAt�h�_	Ps�W�_10��4�R�P01D�VG�J� L�@�J�OGW���TO7RQU��ON*�M����sRHљ��_W��-�_=��C��I���I�I�II�F��`�JLA.�1[�VEC��0�D�BO1Up�@i�B\JRKU���	@DBL_S�Md�BM%`_DLC�BGRV��C��I��H_� ��*COS+\�(LN�7+X>$C�9)I�@9)u*c,)�Z2 �HƺMY@!�( "T�H&-�)THET0�NK23I��"=��A CB6CB=�C �A�B(261C�616�SBC�T25GTS QơC��aS$" ��4c#�7r#$DU D�EX�1s�t��B�6��r.�Q|r�f$NE�D�pIB U�\B5��$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2�&P�C�J�&!�VAHV6HT3�YLVhJVuKV�KUV�KV�KV�KV�IHAHZF`RXM��wXuKUH�KH�KH�KH�KUH�IO2LOAHO�Y�WNOhJOuKO�KO��KO�KO�KO�&F��2#1ic%�d4GSP�BALANCE_l�!�cLEk0H_�%SP��T&�bc&�br&PFULC�hr�g�rr%Ċ1ky�UT�O_?�jT1T2Cy��2N&�v�ϰct�w�g�p�0Ӓ~���T���O���� INSsEGv�!�REV�v�!���DIF��1�l�w�1m�0OB0�q
����MIϰ1�~�LCHWAR��波AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|���7ROBR�CR���N��&�MSK�_�`f�p P 
Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�M?TCOM_C@j�q  L��p��?$NORE³5�y��$�r 8� �GR�E�SD�0A�BF�$XYZ_�DA5A���DEBaU�qI��Q�s �`�$�COD�� ���k�F�f�$BUFINDXРw  ��MOR��/t $-�U��)��r�B��������G�ؒu � $SIMULT ��~��< ���OBJE�` ��ADJUS>�1�A'Y_Ik��D_�����C�_FIF�=�T� ��Ұ��{��p@� �����p�@��D��FRI��ӥT��RIO� ��E�{�͐�OPWO�ŀv}0��SYSBU�@ʐ$SOP�����#�U"��pPRUN,�I�PA�DH�D�\���_OU�=���qn�$}�IMA�G��ˀ�0P�qIM����IN�q���?RGOVRDȡ:����|�P~���Р�0L�_6p���i��RB����0��M���E�DѐF� ��N`Md*���ŷ�˱SL�`�ŀw x $OwVSL�vSDI��DEXm�g�e�9w�$����V� ~�N���@w����Ûǖȳ�M�h ��q<��� x HˁE�F�ATUS���Cp�0àǒ��BTM��*��If���4����\(�ŀy DˀEz�g���PE�r�����
���EXE��V���E�Y�$Ժ ŀz @�ˁ��UP{�h�$�p��XN���9ԼH� �PG"�{� h $SUB���c�@_��01\�M/PWAI��P���ՓLO��-�F�p��$RCVFAILs_C�-�BWD"�|F���DEFSPup | Lˀ`�D�p� U�UNI���S���R`���_UL�pP���P�ā}��� B�~���|�t�`ҲN�`KET��Jy���P� $�~��=�0SIZE��h��{���S<�OR��?FORMAT/p 㰷 F���rEMR���y�UX�����P�LI7�ā  �$�P_SWIp�����_PL7�?AL_ �ސR�A��B�(0C��Dnf�$Eh�����C_=�U� �� � ���~�J�3�0����TIA4���5��6��MOM������� �B�AD��*��* PU70NRW���W ��V����� A$PI�6���	 ��)�4l�}6�9��Q���c�SPEED�PGq�7�D� >D����>tMpt[��SAM�`�痰>��MOV ���$��p�5��5�D�1�$2��������{�Hip�IN?,{�F(b+=$��H*�(_$�+�+GAM�M�f�1{�$GE�T��ĐH�D����
�^pLIBR�ѝI.��$HI��_��Ȑ$*B6E��*8A$>G086LW=e6\<G9�6�86��R��ٰV��$PDCK�DQ�H�_����;" ��z�.%�7�4*�9�� �$IM_SRO�D�s"���LH�"�LE�O�0\H��6@�@�U� �ŀ��P�qUR_S�CR�ӚAZ��S_?SAVE_D�E��NO��CgA�Ҷ� �@�$����I��	�I � %Z[� ��RX"  ��m���"�q�'" �8�Hӱt�W�UPpS��хDM��O� ��.'}q��Cg���@�ʣ�ߑ�R�M�AÂ� � $PY���$WH`'�NG p���H`��Fb��Fb��Fb��PLM���	� 0(h�H�{�X��O��z��Z�eT�M���� pS��C��O__�0_B_�a��_%�� |S����@	�v��v@ �@���w�v��EM���% fR�fr�B��ː��ftP��P�M��QU� ��U�Q��A-�QTH�=�HOL��QHY�S�ES�,�UE���B��O#��  ��P0�|�gAQ���ʠJu���O��ŀ�ɂ�v�-�A;ӝROG��a2D�E�Âv�x_�ĀZ�INFO&���+����b�R�O�I킍 ((@SLEQ/�#�����H�o���S`c0O�0��01EZ0NU�e�_�AUT�Ab�COPY��Ѓ�{��@M��N�����1�P��
� ��RGI���f��X_�Pl�$��(���`�W��P��j@��G���EXT_CYCtb��pr����h�_NA�c!$�\�<�RO�`~]�� � m��POR�ㅣ����SRVt�)����DI �T_l���Ѥ{��ۧ��ۧ �ۧ5٩6J٩7٩8��R�S�BZ쐒��$�F6����PL�A�A^�TAR��@E `�Z��p���<��d� ,(@cFLq`h��@YNL�ꟼM�C���PW�RЍ�쐔e�DE�LAѰ�Y�pAD�#q�QSKIPN�� ĕ�x�O�`�NT!���P_ x���ǚ@�b�p1� 1�1Ǹ�?� �?���>��>�&�>�3�>�9��J2R;쐖� 4��EX� TQ ����ށ�Q���[�K�Fд�8�RDCIf�S �U`�X}�R��#%M!*�0�)��$RGoEAR_0IO�T�JBFLG�igpE	Ra��TC݃�����ӟ2TH2N��� �1�b��Gq TN�0 ����M����`Ib���REF:�1�� l�h���ENAB��lcTPE?@���!(ᭀ�� ��Q�#�~�+2 H�W���2�Қ���"�P4�F�X�j�3�қ{�@��������j�4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:Lj�7�ҟo@�����j�8�����"4Fj�SMSK������a��E�A��MOT-E������@ "�1��Q�IO�5"%Ip��Pb���POWi@쐣  �����X��gpi�쐤��Y"$DSB_SIGN4AȩQi�̰C���tRS�232%�Sb�iDEVICEUS#|�R�RPARIT򱾈!OPBIT�Q���OWCONTR`��Qⱓ�RCU� �M�SUXTASK��3NB��0�$TATU�P��� @@쐩�F�6�_�PC}��$FREEFRO�MS]p�ai�GET\N@S�UPDl�ARB���SP%0����� !m$USAࢰ�az9�L�ERI��0f��pRY�5~"_ľ@f�P�1�!�6WR	K��D9�F9Х?FRIEND�Q4b�UF��&�A@TOO�LHFMY5�$L�ENGTH_VT��FIR�pqC�@�yE� IUFIN�R:���RGI�1�OAITI:�xGX�l�I�FG2�7G1a�0���3�B�GPRR�DA���O_� o0e�I1R�ER�đ�3&���TCp���AQJV�G|�.2���F��1�!d� 9Z�8+5K�+5��E�y�|L0�4�X �0*m�LN�T�3Hz��8P9��%�4�3G��W�0�W�RdD�Z��T�ܳ��K�a3d��$cV 2���1��RI1H�02K2sk3K3Jci�aI�i��a�L��SL��R$V�ؠ�BV�EVk��A (bQ*R��� �,6Lc ���9V2F{/P:B��kPS_�E��$rr8�C�ѳ$A0��wCPR���v�U�cSk��� {�d�"�1���# 0���VX`�!�t�X`��0P�Ё�
z�5SK!� �-q�R��!0���z�N�J AX�!h�A�@LxlA��A�THIC�1��������1TFE����q>�IF_CH��3A�I0�����G�1�x������9�nɆ_JF҇PR(����RVAT�� �-p��7@����sDO�E��COU(���AXIg��OF�FSE+�TRIG �SK��c���Ѽ�e�[��K�Hk���8�IGM�Ao0�A-��ҙ�ORG_UNEV�Ξ� �S�쐮Od �$�������GROU��ݓTO�2��!ݓDSP��JcOG'��#	�_P'��2OR���>P6KEPl�IR�0�P�M�RQ�AP�Q��Ep�0q�e���SYSG���"��PG��BRK *Rd�r�3�-�������ߒ<pAD��ݓJ�OBSOC� N�DUMMY14�p�\@SV�PDE_O�P3SFSPD_WOVR��ٰCO�L�"�OR-��N�0b.�Fr�.��OV�CSFc�2�f��F���!4�S��RA�"LC�HDL�RECOQV��0�W�@M��յ�RO3��_��0� @�ҹ@V�ERE�$OFSf�@CV� 0BWDG��ѴC��2j�
�TR��!��E_FD}Oj�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��2_�Gxǋ�AM��k�0J0������_M��2x{�#�8$CA��{Й���8$HBKX|1c��IO��.�:!aPPA"�N�3��^�F���:"�DVC_DB�C��d�w"�Ј��!��1���ç�3�����ATIO� ��q0�UC�&CAB�BS�PⳍPȲȖ��_0c�SUOBCPUq��S�P a aá�}0�Sb��c���r"ơ$HW_C ���:c��IcA�A-��l$UNIT��l���ATN�f����C�YCLųNECA���[�FLTR_2_FI���(��}&���LP&�����_SC-T@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb�r�v: _T��PRO��,O�� EM�_��98u�q u�q���DI�0e�RAI�LAC��}RMƐL!OԠdC��:anq��Xwq����PR��SLQIkfC�ѷ 	���FUNCŢ�rRI�NkP+a�0 ��!RA� >R 
Я��ԯWAR�BLFQ��A�����DA�����LDm0�aB9��nqBTIvrbؑ����PRIAQ1�"AFS�P�!����P�`%b���M�I1U�DF_j@��y1°�LME�FA�@HR�DY�4��Pn@RS�@Q�0"�MULS�Ej@f�b�q ��X��ȑ���$�.A$�1$c1�Ó���� x�~�EG70ݓ�q!A1R����09>B�%���AXE��RO%B��W�A4�_�-֣CSY���!6��&S�'�WR���-1���SCTR��5�9�E�� 	5B��=QB�90�@6������OT��0o 	$�ARAY8�w20���	%��FI��;�$LI�NK�H��1�a_�63�5�q�2XYZ"��;�q�3@��1)�2�8{0B�{�D��� CFI���6G��
�{�_�J��6��3aOP�_O4Y;5�QTB�mA"�BC
�z�DU�"�66CTURN 3�vr�E�1�9�ҍGFL�`���~ �@�5�<:7�� 1�J?0K�Mc�68Cpb�vrb�4�ORQ�� X�>8�#op�������wq�Uf�����TOV	E�Q��M;�E#�UK#�UQ"�VW�ZQ�W ���Tυ� ;����Q H�!`�ҽ��U�Q�Wke0K#kecXER���	GE	0��S�dA WaǢ:D���7!�!AX�rB!{q�� �1uy-!y�pz �@z�@z6Pz\Pz � z1v�y�y �+y�;y�Ky�[y �ky�{y��y�q�yoDEBU��$� ���L�!º2WG`  CAB!�,��SV���� 
w���m��� w����1���1���A�� �A��6Q��\Q���!�pm@��2CLAB3B��U�����S � ÐER��
0 O� $�@� Aؑ!p�PO��Z�xq0w�^�_MRAȑ_� d  T��-�ERR��T)Yz�B�I�V3@�cNΑTOQ�d:`L� H�d2�]�X�C[!_ � p�`T}0i��_V1�r�a'�4�2-�2<�����@P�����F�$W���g��V_!�l�$�P����c��q"��	�SFZN_wCFG_!� 4�� ?º�|�ų����@�ȲW [V ��\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(����$�!s�Q�g�P{RV �HELLĥ�� 56�B_BAS�!�RSR��ԣo ��#S��[��1r�%���2ݺ3ݺ4ݺ5*ݺ6ݺ7ݺ8ݷ���ROOI䰝0�0NLK!�CAB� ���ACK��IN��T�:�1�@�@ z�m�_�PU!�CO� ��OU��P� Ҧ) ��޶���TPFWD_�KARӑ��RE�~��P��(�QU�E�����P
��CSTOPI_AL������0&���㰑�0S#EMl�b�|�M��dЛTY|�SOK�}�D�I�����(���_�TM\�MANRQ�ֿ0E+�|�$K�EYSWITCH�&	���HE
�B�EAT��cE� LQEҒ���U��FO������O_HOM��O�REF�PPARz��!&0��C+�9OA�ECO��B<�rIOCM�D8׆��]���8�` �# D�1����U��&��MH�»P�CFOR�C��� p ��O}M�  � @V�T�|�U,3P� 1-��`� 3-�4��N�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��C@�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fim7s�&��VP��UPD��  ���|�԰��YSL}OǢ� � z� �и���o�E��`>�^t��АALUץ�����CU���wFOqID�_L�ӿuHI�zI~�$FILE_����t��$`�JvSAΒ�� h���E_BLCK�#�C,�D_CPU<�{�<��o����tJr��Rw ��
PW �O� ��LA��Sp��������RUNF� Ɂ��Ɂ����F�ꁡ�|ꁬ� �TBCu��C� �X -$�LENi��v�������I��G�LO�W_AXI�F1��t2X�M����D�4
 ��I�� ��}�GTOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑTCV����T���&��ݡ����HJ�����J����Mo�"��J�Ǜ �������2��� v�����6F�JK��VKi�Ρ4v�Ρ3��J0�ң�JJڣJJ�AAALң�ڣ��4�5z�&�N1-�9����␅�L~�_Vj��x+p���� ` ��GROU�pD��B>�NFLIC��REQUIREa�EBUA��p����2¯�����c��� \��APP�R��C���
�E�N�CLOe��SC_M v�,ɣ�
�ޣ�� ���MCp�&���g�_MG�q�C� �{�9���|�wBRKz�NOL��t|ĉ R��_LI|�H�Ǫ�k�J����P
� ��ڣ�����&���/�"��6��6��8��Y�|���� ���8�%�W�2�e�PATHa�z�p�z�=�vӴ��ϰ�x�CN=�CaA�����p�IN��UC��bq��CO�U�M��YZ������qE�%���2������PA�YLOA��J2L�3pR_AN��<�L���F�B�6�R�{�R_?F2LSHR��|�LOG��р��ӎ���ACRL_u��������.���H�p�$yH{���FLEX
��s�J�� :�/����6�2���0��;�M�_�F16�� ��n���������ȟ��Eҟ�����,�>� P�b���d�{�����@�������5�T��X��v���Eť mFѯ��������&�/�A�S�e�D�J>x�� � ������j�4pAT����n��EL  �%øJڪ��ʰJE��CTYR�Ѭ�TN��F&���HAND_VB�[
�pK�� $�F2{�6� �rS�Wi��r�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�
�K�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������uN���2�H̟�����"CqENL� �pDI��>�Obtq D�Dpx�� �
�2IxQA����q���-��s �� �����{ ��OMME���rr/�TVpP�T�P ���qe�i� ���P�x ��yT�Pj�� $DUMM�Y9�$PS_f��RFq�sp$:�� ���!~q�c X����K�STs��ʰSBR��M2�1_Vt�8$SV_ERt�O��z���WCLRx�A  O�r�?p? Oր � �D $GLOB���#LO��Յ$�po��P�!SYS�ADR�!?p�pTC}HM0 � ,�����W_NA���/�e�$%SR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T�RF�TXSCR�E�ƀ�� ��STF���}�pТ6�SQP] _v AŁ�� T����TYP �r�K��u�!u����O�@IS�!���uD�UE{t� �����H�S���!R�SM_�XuUNE�XCEPWv��CpS_��{ᦵ�ӕ���÷���COU ���o 1�O�UET��փr���PROG�M� FLn!$CMU��PO*q��d��I_�pH;� �s 8��N�_HE
p���Q��pRY �?���,�J�*���c�?�OUS�� �� @d���$B�UTT��R@���C�OLUM�íu�S�ERVc#=�PAN�Ev Ł� � N�PGEU�!�F��~9�)$HELP��^WRETER��)� ����Q�������@� P�P �IN��s�PNߠw v��1����� ����LN�� �䟀�_��k�$H��M TEX�#�����FLAn +REL�V��D4p�������M��?,��ӛ$�����P=�USR�VIEWŁ� <�d��pU�p0NFyIn i�FOCU��ni�PRILPm+��q��TRIP)��m�UNjp{t� �QP��XuWARN|Wud�SRTOLS��ݕ�����O|SO;RN��RAUư��9T��%��VI|�zu�� $�P�ATHg��CAC�HLOG6�O�LIMybM���'��"��HOST6�!��r1�R�OBOT,5���IMl� D�C� g!��E�L���i��VCPU_AVA�ILB�O�EX7�!BQNL�(���A�� Q���Q ��ƀ��  QpC���@_$TOOL6�$��_JMP� �<I�u$SS�!$>��VSHIF��|s�P�p�6�s���yR���OSUR=W�pRADIz��2�_�q�h�g! �q�)�LUza$O�UTPUT_BM��IML�oR6(`�)�@TIL<SC	O�@Ce�;��9 ��F��T��a��o��>�3�����w�2Ju�( V�zu���%�DJU��|#�/WAIT����ک�%ONE��Y�BOư ��� $@p%�C�SB�n)TPE��NEC���x"�$t$���*B_T��R��%�qR� $���sB�%�tM�+���t�.�F�R!݀��O�Pm�MAS�_DUOG�OaT	�D�����C3S�	�O2DELcAY���e2JO�� n8E��Ss4'#J�aP60%�����Y_��O2�$��2���5��`?� �=pZABC~S��  $�2��J�
sp�$$C�LAS������Asp�'@@VI�RT��O.@ABS��$�1 <E�� < *AtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v�����M@�[�AXLր`�&A�ndC  ���IN��ā��PRE������LARMRECOV <Il䂥�NG�� \K	 =#�
J�|\�M@PPLIC��?<E�E��Handlin�gTool �� �
V7.50P�/28 *A��^���
�_SW UP*A� F��F0ڑ����A�~�� 20�К*A���	Ց��h�j(B �7DA5��  ~'@�^@�𞝓None������� ��T�y�*A4�]x��P_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ��i�n�����#B)B ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��&��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���o&�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� ��PB�Z?����5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`��S:��r������Up�_)o�S  K�3Ph���R�PX�_mo8j����a�Oko�o9i�(�+(�9!Rhg�o�o�l�Kof�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`(ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCPU�eB��CF��;.<C����C5`SXE@D��nyDQ��D���>��D�;D�����F��>F�$�G}RB�7Gzր��SY��)!�vqG���Em�U(�.��(�(�1�<�q�G�x2��eҢ �� a�D�j�怀ES\E@EX��EQ�EJP� F�E�F�� G�ǎ^F� E�� FB�� H,- Ge�߀H3Y��� � >�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE ��O@b 
�(�;��"�  <�6�z�Rb���?�j�C4�)�SZm� W��{�Jm�C��B-G�Cu��@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"�� , 
�^��P�o xvf`MT�I^��rl@�:sONTImM������Zv�i
õ�cMOTN�END���dREC�ORD 1(R�8a��ua�O��q� �sb�.�@�R��xZ� ������ɏۏ폄� ��#���G���k�}��� ��<�ş4��X��� 1�C���g�֟������ ��ӯ�T�	�x�-��� Q�c�u���������� >����)Ϙ�Mϼ� F�࿕ϧϹ���:��� ����%�s`Pn&�]�o� �ϓ�~ߌ���8�J��� ��5� ��k����� ���J�����X��|� ��C�U�����������0�����	��dbTOLERENCqdsBȺb`L�͐P�CS_CFG �)�k)wdMC�:\O L%04dO.CSV
�Pc��)sA �CH� z�P)~���hM�RC_OUT �*�[�`+P SG�N +�e�r���#�10-MAY�-20 10:4�7*V27-JAN�j21:48�k? P;����)~�`pa�m��PJPѬ�VERSION� SV2�.0.�6tEFLOGIC 1,�[/ 	DX�P7)��PF."PROG_�ENB�o�rj UL�Sew �T�"_WRSTJNEp�V�r�`dEMO_OPT?_SL ?	�es�
 	R575)s7)�/??*?<?|'�$TO  �-د�?&V_@pEX�Wd�u�3PAT�H ASA\p�?�?O/{ICT�a-Fo`-�gds�egM%&ASTBF_TTS�x@�Y^C��SqqF�P�MAU� t/XrMS%WR.�i6.|
S/�Z!D_N�O0_�_T_C_x_g_�_�tSBL_FAUL"y0�[3wTDIAU �16M6p�A�1234567G890gFP? BoTofoxo�o�o�o�o �o�o�o,>Phb�S�pP�_ ���_s�� 0`�� ���)�;�M�_�q� ��������ˏݏ��|�)UMP�!� �^�TR�B�#+�=��PMEfEI�Y_T�EMP9 È�3p@�3A v�UNI�.�(YN_BRK �2Y)EMGDI_STA�%W!b�ՐNC2_SCR 3��1o"�4� F�X�fv���������#��ޑ14���@�)�;�����ݤ5�����x�f	u� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/߭P�b� t�� ��xߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N���r��� ������������ &8J\n��� �����"`� FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/4?,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O?�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�O�O�o �o�o
.@Rd v������� ��*�<�N�`�r��� �o����̏ޏ���� &�8�J�\�n����������ȟڟ����H�E�TMODE 16v��� ���ƨ
R�d�v�נR�ROR_PROG7 %A�%�:߽��  ��TABLE  A�������#�L�RRSEV_?NUM  ��Q���K�S���_�AUTO_ENB�  ��I�Ϥ_N�Oh� 7A�{��R�  *����J��������^�+��pĿֿ迄�HISO��͡I�}�_ALM �18A� �;�����+�e�wωϐ�ϭϿ��_H���  A���|��4��TCP_VER �!A�!����$E�XTLOG_RE�Q��{�V�SI�Z_�Q�TOL  �͡Dz��=�#׍�XT_BW�D����r���n�_D�I�� 9���}�z�͡m���STE�P����4��OP_�DO���ѠFA�CTORY_TU�N�dG�EATU�RE :�����l�Hand�lingTool� ��  - C�English� Diction�ary��ORDE�AA Vis��� Master����96 H��n�alog I/O����H551��u�to Softw�are Upda�te  ��J��m�atic Bac�kup��Part�&�groun�d Edit�� � 8\apC_amera��F���t\j6R�ell����LOADR�o�mm��shq��T7I" ��co���
! o���pa�ne�� 
!���tyle se�lect��H59��nD���onit�or��48����t�r��Reliab����adinDiagnos"�����2�2 ual �Check Sa�fety UIF� lg\a��ha�nced Rob� Serv q �ct\��lUse�r FrU��DI�F��Ext. D�IO ��fiA �d��endr E�rr L@��IF��r��  �П�9�0��FCTN M�enuZ v'��7}4� TP In���fac  SU_ (G=�p��_k Excn g��3��High-S�per Ski+� � sO�H9 � mm�unic!�onsg�teur� �����V����coknn��2��EN���Incrstr�u���5.fd�KAREL C�md. L?ua�A� O�Run-;Ti� Env����K� ��+%�s#�S�/W��74��Li�censeT� � (Au* ogB�ook(Sy��m�)��"
M�ACROs,V/�Offse��ap���MH� ����pf�a5�MechStop Prot��� d�b i�S�hif���j54�5�!xr ��#��,��lb ode �Switch��mK\e�!o4.�&� pro�4��g���Multi-�T7G��net.�Pos Re�gi��z�P��t� Fun���3 9Rz1��Numx ������9m�1�  A�djuj��1 J�7�7�* ����6t�atuq1EIKoRDMtot��_scove�� ���@By- }ues�t1�$Go� � U5\�SNPX b�"���YA�"LibAr����#�� �$�~@h�pd]0�Jt�s in VCC!M�����0�  �u!Ξ�2 R�0�/I��08��TMIL{IB�M J92�@�P�Acc>�F�9=7�TPTX�+�B�RSQelZ0�M8� Rm��q%��69�2��Unexce{ptr motnT  CVV�P���KC����+-��~K�  II)�VSP� CSXC�&.c��� e�"�� t�@�Wew�AD �Q�8bvr nmeYn�@�iP� a0�y�0�pfGrid~Aplay !� �nh�@*�3R�1M-1�0iA(B2015 �`2V"  F����scii�loa�d��83 M��l�����Guar�d 'J85�0�mP'�L`����stuaPat�&]$Cyc���|0�ori_ x%Dat�a'Pqu���ch��1��g`� j� RLJam�5���I_MI De-B(\A^�cP" #^0C�  etkc^0a�sswo%q�)65�0�ApU�Xnt\��Pven�CTq�H�5�0YEL?LOW BO?Y���� Arc�0vis���Ch�Weld�Qcial4Izt��Op� ��gs�` �2@�a��poG yRjT1 NE�#3HT� xyWb��#! �p�`gd`����p\� =P��JPN� ARCP*PRx�A�� OL�pwSup̂fil�pp��J�� ��cro�6�70�1C~E�d��SuS�pe�tex�$Y �P� So7 t� /ssagN5 <Q�B�P:� �9 "0�Qr�tQC��P�l0dpn�笔�rpf�q�e��ppmasc�bin4psyn��' ptx]08�H�ELNCL V�IS PKGS �Z@MB &��B� J8@IPE �GET_VAR �FI?S (Uni�� LU�OOL: �ADD�@29.F�D�TCm���E�@D�Vp���`A�ТNO� WTWTEST� �� ��!��c�F�OR ��ECT ��a!� ALSE �ALA`�CPMO�-130��� b D�: HANG F�ROMg��2��R�709 DRAM� AVAILCH�ECKS 549���m�VPCS S�U֐LIMCHK���P�0x�FF P�OS� F�� q�8-12 CH�ARS�ER6�OG�RA ��Z@AVE�H�AME��.SV���Вאn$��9�m� "y�TRCv� �SHADP�UPD�AT k�0��ST�ATI��� MU�CH ���TIM�Q MOTN-0�03��@OBO�GUIDE DAUGH���b��@$Gtou� �@C� �0���PATH�_�M�OVET�� R6�4��VMXPAC�K MAY AS�SERTjS��CY�CL`�TA��BE COR 71�1�-�AN��RC O�PTIONS  ��`��APSH-1N�`fix��2�SO���B��XO򝡞�_TP��	�i��0j��du�{byz p wa���y�٠HI������U��pb XSPD T�B/�F� \hch�ΤB0���END�C�E�06\Q�p{ s>may n@�p�k��L ��traff#�	� ��~1�from sysvar scr�0qR� ��d�DJU����H�!A��/��S?ET ERR�D��P7����NDAN�T SCREEN� UNREA V�M �PD�D��PA����R�IO J�NN�0�FI��B���GROUNנD� Y�Т٠�h�S�VIP 53 QS���DIGIT V�ERS��ká�NE�W�� P06�@C�1IMAG�ͱ���8� DI`���p�SSUE�5��EP�LAN JON� gDEL���157QzאD��CALLI�ॡQ��m���IPN�D}�IMG N9� PZ�19��MN;T/��ES ���`wLocR Hol߀�=��2�Pn� PG:t��=�M��can������С: 3D �mE2view d3 X��ea1 �0�b�pof Ǡ"H�Cɰ�ANNOT� ACCESS �M cpie$Etn.Qs a� loMd�Flex)a:��w^$qmo G�sA9�a-'p~0��h0pa���eJ AUTO-�0��!ipu@Т<ᾡ�IABLE+� �7�a FPLN: �L�pl m� M�D<�VI�и�WI�T HOC�Jo�~1Qui��"��N���USB�@�Pt & remov����D�vAxis F�T_7�PGɰCP�:�OS-144� � h s 26�8QՐOST�p  �CRASH DU���$P��WORD�.$�LOGIN̈P��P:	�0�046 issueE��H�: Slow� st�c�`6Й���໰IF�IM�PR��SPOT:�Wh4���N1STY<��0VMGR�b�N�CAT��4oRR�E�� � 58t�1��:%�RTU!Pre -M a�SE:�@!pp���AGpL��9m@all��*0va�OCB WA����"3 CNT0 �T9DWroO0al�arm�ˀm0d �t�M�"0�2|� o�Z@OME<�� ���E%  #1-�SR�E��M�st}0g �    5KA�NJI5no M�NS@�INIS�ITALIZ'� E�f�we��6@� �dr�@ fp "~��SCII L�afails w�>�SYSTE[��i��  � Mq�1�QGro8�m n@�@vA����&��n᰼0q��RWRI O�F Lk��� \r�ef"�
�up� d�e-rela�Qd� 03.�0SSc}hőbetwe4�IND ex ɰTPa�DO� l�y �ɰGigE�s�operabil.`p l,��HcB�̚@]�le�Q0cf�lxz�Ð���OS� {����v4pfigi GLA�$�c2��7H� lap�0A[SB� If��g�2 l\c�0�/��E�� EXCE �㰁�P���i�� Do0��Gd`]Ц�fq��l lxt��EFal��#0�i�O�Y��n�CLOS��SR�Nq1NT^�F�U�FqKP�ANIO V7/ॠ1�{����DB �0��ᴥ�;ED��DET|�'�� �bF�NLINEb�BUG�T���C"RLIB��A���ABC JARK�Y@��� rkey��`IL���PR��N\��ITGAR� D$��R �Er *�T���a�U�0��h�[�Z�E V� TAS�K p.vr�P�2" .�XfJ�srn8�S谥dIBP	c�v��B/��BUS��UNN� j0-�{�d�cR'���LOE�wDIVS�CULs0$cb����BW!���R~�W`P�����ITd(঱tʠ�OF���UNEXڠ+���p��FtE��SVEM�G3`NML 50�5� D*�CC_SAFE�P*� �ꐺ� PET��'P�`�gF  !���IR����c i S>� K���K�H GUN�CHG��S�MEKCH��M��T*��%p6u��tPORY_ LEAK�J����SPEgD��2Vw 74\GRI�x�Q�g��CTLN��TRe @�_�p ���EN'�IN�����0�$���r��T3)�iԗSTO�A�s�L���͐X	���q��Y� ��TO2�J m���0F<�K����DU��S��O��3 �9�J F�&���SSVGN-1#I���'RSRwQDAU�Cޱ � �T6�g��� 3�]�~��BRKCTR/"� �q\j5��_�QܺS�qINVJ0D ZO�Pݲ���s��г��Ui ɰ̒�a�DU{AL� J50e��x�RVO117 AW�TH!Hr%�N�7247%�52��|�&aol ���R���at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���Md��Rǰt� \fosB�A�0Np�c�����{�U��ROP 2��b�pB��ITP4aM��b !AUt �c0< � plete��N@� z1^qR�635 (Acc_uCal2kA���I) "�ǰ�1a\�Ps��ǐ� bЧ0�P򶲊���ig\�cbacul "A3p_ �1��ն���_etaca��AT����PC�`�����_p�.pc!Ɗ��:�circB���5��tl��Bɵ�:�fm+�Ί�V�b�ɦ�r�?upfrm.����ⴊ�xed��Ί�~�'pedA�D �}b�ptlibB�� ߆_�rt��	Ċ�_0\׊ۊ�6�fm�݊��oޢ�e��̆Ϙ���c��Ӳ�5�j>�����tcȐ��	�r����emm 1��T�sl^0���T�mѡ�#�rm�3��ub Y�q�st�d}��pl;�&�c1kv�=�r�vf�䊰���9�vi����u�l�`�0fp�q �.yf��� daq; �i Data Ac_quisi��n��
��T`��1�8�9��22 DMCM RRS2Z��75��9 3 Rg710�o59pq5\?��T "���1 (D�T� n k@��������E Ƒȵx��Ӹ�etdmm F��ER����gE<��1�q\mo?۳ �=(G���[(

�2�` ! �@J�MACRO��Sk�ip/OffseP:�a��V�4o9� &qR662���Rs�H�
 6Bq8�����9Z�43 J�77� 6�J783�o ��n�"v��R5IKCBq2� PTLC�Zg� R�3 (�s,� �������03��	зJԷ\sfm�nmc "MNM�C����ҹ�%mnf�FMC"Ѻ0ª etmcr� �8����� ,��lD�l �  874\prdq>,jF0����axisHPro�cess Axe�s e�rol^P�RA
�Dp� 56 �J81j�59� 5�6o6� ���0w�6�90 98� [!IDV�1��2(x2��2ont�0�
�����m2���?C��etis "ISD��x9�� FpraxRA�M�P� D��de�fB�,�G�isb/asicHB�@޲�{6�� 708�6
��(�Acw:�����@�D
�/,��AMOX��  ��DvE��?;T��>Pi� RAFM';�]�!PAM�V�W�Ee�U0�Q'
bU�75�.��ceNe� nterface^�1' �5&!54�K��b(Devam±�/�#��Э/<�Tane`"D�NEWE���btpd/nui �AI�_s~2�d_rsono����bAsfjN��bdv_arFvf�xhp�z�}w��hkH9xs�tc��gAponlGzv{�ff��r ���z�3{q'Td~>pchampr;re�p� ^5977� �	܀�4}0��mɁ�/������lf�!�pcc7hmp]aMP&B<�� �mpev������pcs��YeS~�� Macro�O	D��16Q!)*�:$��2U"_,��Y�(PC ��$_;������o|��J�gegemQ@�GEMSW�~ZG�g�esndy��OD�n�dda��S��syT�Kɓ�su^Ҋ����n�m���L��  �	��9:p'ѳ޲���spotplus�p���`-�W�l�J�s⽱t[�׷p�key �ɰ�$��s�-Ѩ�m�~��\featu 0�FEAWD�oolo�srn'!2 �p���a�As3��tT�.� (N. A.)��!e!�J# (j�,��oBIB�o�D -�.�n��k9�"K��u[-�_���}p� "PSEq�W����wop "sEЅ�&�:�J����� �y�|��O8��5��R ɺ���ɰ[��X�� �����%�(
ҭ�q HL�0k�
�z�a !�B�Q�"(g�Q �����]�'�.����ɀ&���<�!ҝ_�#��tpJ�H�~Z��j����� y������2��e��� ���Z����V��!%���=�]�͂��^2�@i[RV� on�QYq͋JF0� 8ހ�`�	�(^�dQueue���X\1�ʖ`�+F1�tpvtsn��N�&��ftpJ0v �R�DV�	f��J1 Q4���v�en��k/vstk��mp��~btkclrq���get�����r��`kack8�XZ�strŬ�%��stl��~Z�np:!�`���q/��ڡ6!l�/Yr�mc�N+v3�_� ���l�.v�/\jF��� �`Q�΋ܒ��N50 (FRA���+��͢frap�arm��Ҁ�} 6��J643p:V�E�LSE
#�VA�R $SGSYS�CFG.$�`_U?NITS 2�DG0~°@�4Jgfr��4A�@FRL-��0ͅ�3 ې���L�0NE�:� =�?@�8�v�9~Qx3�04��;�BPRS�M~QA�5TX.$VNUM_OL��85��DJ507��l�? Functʂ"q�wAP��琉�3 HH�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6 N�kAP����S��"TPPR���Q.A�prnaSV�ZSx��AS8Dj510U�-�`cr�`8 ��ʇ��DJR`jYȑH � �Q �PJ�6�a21��48AAVM 5�Q�b0 lB�`TUP� xbJ5459 `b�`616���0VCAM 9��CLIO b1��5 ���`M�SC8�
rP R`\�sSTYL �MNIN�`J62�8Q  �`NRExd�;@�`SCH ���9pDCSU Me�te�`ORSR �Ԃ�a04 kR_EIOC �a5�`542�b9vpP<� nP�a�`�R�`7�`��MASK H�o�.r7 �2�`O'CO :��r3��p�b�p���r0X��a�`�13\mn�a39 HRM"�q�q�ҿLCHK�uO�PLG B��a03� �q.�pHCR �Ob�pCpPosi��`fP6 is[rJ�554�òpDSWĤbM�D�pqR�a37� }Rjr0 �1�s4i �R6�7��52�rs5 �2�r7 1� �P6���Regi��@T�uFRDM��uSaq%�4�`93�0�uSNBA�uSwHLB̀\sf"p�M�NPI�SP{VC�J520���TC�`"MNрT�MIL�IFV�P�AC W�pTPT�Xp6.%�TEL�N N Me�0�9m3UECK��b�`UFR�`��V�COR��VIPL:pq89qSXC�S�`�VVF�J�TP ��q��R626l�u� S�`Gސ�2�IGUI�C��PG�St�\ŀH863`�S�q�����q34sŁ684���a��@b>�3 :B��1 \T��96 .�+E�g51 y�q53�3f�b1 ���b1 n��jr9 ���`VAT9 ߲�q75 s�F�<�`�sAWSM��`�TOP u�ŀR582p���a80 
�ށgXY q���0 ,b��`885�QXрO�Lp}�"pE࠱tp��`LCMD��ET3SS���6 �V��CPE oZ1�V�RCd3
�NLH�h���001m2Ep��3� f��p��4 /1�65C��6l���7zPR��008 tB~��9 -200�`�U0�pF�1޲1 ��޲2L"���p��޲y4��5 \hmp~޲6 RBCF�`0ళ�fs�8 �Ҋ���~�J�7 rbc	fA�L�8\PC�����"�32m0u�n�K�R�ٰn�5 5EW�
n�9 z��40Y kB��3 ��6ݲ��`00iB/��6$�u��7�u��8 µ������sU0�`�t �1 05\rb��2 E���K���j�2��5˰��60��a�HУ`:�63�jAF�_����F�7 ڱ݀H�80�eHЋ��cU0��I7�p��1u��8u��9 73�������D7� ��5t�9+7 ��8U�1��2J��1�1:���h���1np�"��8(�U1��\pyl��,࿱�v ��B�854��1hV���D�4��im�с1�<���>br�3�pr�4@pGPr�6 !B���цp��1�����1�`͵155ض1g57 �2��62�S����1b��2����1Π"�2���B�6`�1<c�4 L7B�5 DR��8_�{B/��187 u�J�8 06�90� rBn�1 (��202 0EW,ѱ�2^��2��90�U2��p�2��2 b��4:��2�a"RB����9\�U2�`w�l���O4 60Mp��7��`����b�s
5 ���3����pB"9 3a ����`ڰR,:�7 �2��V�2��5@���2^��a^9��B�qr����n�5����5᥁"�8a�Ɂ}Չ5B���5����`U�A���� ��86 �6 S�0��5�p�2�#�529 �2^�Tb1P�5~�2`P���&P5��8��5��u�!�5��ٵ5+44��5��R�ąPa nB^z�c (�a4�����U5J�
V�5��1�1^��%������5 b21���gA��58W8-2� rb��5N�E�G5890r� 1�95 �"������c 8"a��|�L ���!J"E5|6��^!�6���B�"8�`#��+�8�%�6B�AME�"1w iC��622�B�u�6V��d� 4��8�4�`ANRSP�e?/S� C�5� �6� ��� \� �6� ��V� 3t��� TG20CA�R��8� pHf� 1DH�� AOE�� �� ,�|�� �0\�� �!64K��ԓrA� �1� (M-7�!/50T�[PM��P�Th:1�C�#Pe� �3��0� 5`M75T1"� �D8p� �0Gc�� u�4��i1-710i�1� Skd�7j�z�?6�:-HS,�  �RN�@�UB�f�X�=m75sA*A6a�n���!/CB�B2.6A �0;A�CIB�A�2P�QF1�UB2�21� �/70�S� �4��� �Aj1�3p���r�#0 B2\m*A@C@��;bi"i1K�u"A~A�AU� imm7c7@��ZA@I�@�Df�Ab�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A��EA�5B�4>\77
B7=Q�D�2�Q$B�E)7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E"l7�@7�A
1�E�V~`��W2%Q�R9ї@0L_�#����"A����b��H3s=rA/2 �R5nR4�74rNUQ1�ZU�A�s\m9
1M�92L2�!F!^Y�ps�� 2ci��-?�qhimQ�t  w043�C�p�2�mQ�r�H_ �H20��Evr�QHsXBSt62�q`s����� ��P�xq350_*A3I)�2�d�u0�@� '4kTX�0�pa3i1�A3sQ25�c��s�t�r�VR1%e�q0 
��j1��O2 �A �UEiy�.�‐ �0C2h20$CXB79#A�����M Q1]�~�� 9 �Q��?PQ��qA!Pvs � 5	15aU���?P�Ņ���ဝQ9A6�zS*�7�qb5�1��8��Q��00P(��V7]u�aitE1���ïp�?7� !?�z��rbUQRB1PM=�Qa9p��H��QQ�25L��@�����Q��@L���8ܰ��y00\r�y�"R2BL�tN�  ��� �1D�l�2�qeR�5���_b�3�X]1/m1lcqP1�a�ED�Q� 5F����!5���@M-16Q�� f� ��r��Q�e� ��� PN�LT_�1��i1��9453��@�e�|�b1l>F1u*AY2�
��R8�Q���RJ�J3�D}T� 85
Qg�/0��*A!P� *A�Ð𫿽�2ǿپ6t�6=Q���P�X���� AQ� g� *ASt]1^u�ajrI�B ����~�|I�b��yI�\m�Qb�I�uz�A��c3Apa9q� B6S���S��m���}�85�`N�N�   �(M���f1���6��P��161��5�s`҃SC��U��A����5\set06c��f��10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C����5�B��B��h`�F��� X0���A:���C�M��!AZ��@��4�6i����� e�O�-	���f 1��F �ᱦ�1F�8Y	���T6HL3��BU66~`���U�dU�9D20Lf0��Qv�  ��fjq��N������ 0v
� ��i	�	��72lqQ2�������� \chngmOove.V��d��|��@2l_arf 	�f~��6���� ��9C�Z���~���kr41 S���0��V���t�����U�p7nuqQ%�A]��V�1\�Qn�BJ�2W�EM!5���)�#:�64��F�e50S�\��0�=� PV���e�������E�����m7shqQSH"U��)��9�!A��(���� ,�l�����TR1!��,�6�0e=�4F�����2��	 R-������ �����Ж��4���LSR�)"�!lO�A��Q�) %!� 16�
U/��2�"2�E��9p���2X� SA/Ai��'�
7F�H�@ !B�0��D���5V� �@2cVE��p��T��pt갖�1L~E�#�Fd�Q��9E�#De/��RT��59���	�A�E�iR������9\m20�20��+�-u�19r4�`�E1�=` O9`�1"ae��O��2��_$W}am41��4�3�/d1c_std��1)�!�`�_T��r�_ 4\jdg�a�q�PJ%!~` -�r�+bgB��#c'300�Y�5j�QpQb1�bq��vB��v�25�U�����qm43� �Q<W�"Ps� �A��e����t� i�P�W.��c�F�X.�e�kE14�4y4�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf��`coWo!\�2a��K2A;_2��QW2�`bF�(�V11�23�`���X5�Ra21�J�*9�a:88J9X�l5�m1a첚��*���(85�&��������P6���R,52&A����,fA9IfI'50\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP 1��vB)e�m�����ު1p� �1D��l�27�F�KAR�EL Use S���FCTN��� �J97�FA+�� �(�Q޵�p%�)?�Vj�9F?(�j�Rtk208 "Km�6Q�yB�j��iæPr�9�sx#��v�krcfp��RCFt3���Q��k�cctme�!ME�g����6�mainj�dV�� ��ru��kDº�c���o����&J�dt�F �»��.vrT�f�����E�%�!��5�FRj73�B�K���UER�HJn�O  J�� (ڳF���F�q�Y�&T��`p�F�z��19�tkvBr���V�h�9p�E�y�<�k������;�v���"CT��f���� )�
І��)�V	�6� ���!��qFF��1q� ��=�����O�?�$"����$��je���TC�P Aut�r�<5�20 H5�J5�3E193��9��96�!8��9��	 �B�574��52�J:e�(�� Se%!Y������u��ma�Pqtool�ԕ�����~�conrel�F�trol Rel�iable�RmvCU!��H51�����8 a551e"�CNRE¹I��c�&��it�l\s�futst "UaTա��"X�\u�� g@�i�6Q]V0�B,Eѝ6A� �Q�)C ���X��Yf�I�1|�6s@6i��T6I U��vR�d�
$e%1���2�C58�E6��8`�Pv�iV4OFH58SOteJ� mvBM6E~O58�I�0�E�#+@� &�F�0���F�P6a����)/++�</N)0\�tr1�����P ,�lɶ�rmask�i�msk�aA���k�y'd�h	A	�P�sD�isplayIm��`v����J887# ("A��+Heůצprds��Iϩǅ�Uh�0pl�2�R2���:�Gt�@��PRD �TɈ�r�C�@Fm��D��Q�AscaҦ� �V<Q&��bVvbrl �eې@��^S��&5U�f�j8710�yl 	��Uq���7�&�p��p��P^@�P�firmQ����Pp�2�=b�k�6�r�3��6��t7ppl��PL���O�p<b�ac�q	��g1�J�U�d�J��gait_9e��Y�&��Q����	�Shap��e?ration�0��R67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G����qF�205p�5pS���Ձ�retsap��BP�O�\s� O"GCR�ö? �q/ngda�G���V��st2axU��Aa]��bad�_�btputl/�&�e�>��tplibB_���=�2.����5���c3ird�v�slp���x�hex��v�re8?�Ɵx�key�v�cpm��x�us$�6�gcr��F�����8�[�q27j92�v��ollismqSk��9O�ݝ� (pl�.���t��p!o��2 9$Fo8��cg7no@ƿtptcls` C�LS�o�b�\�km�ai_
�s>�v�o	��t�b���ӿ�E�H��6�1enu5�01�[m��uti|a|$calmaUR���CalMateNT;R51%�i=1]@ -��/V� ��Z�� �tfq1�9 "K9E��L����2m�CLcMTq�S#��et ��LM3!} �F�c��nspQ�c���c�_moq��� ��c1_e�����su��ޏ� �_ �@�5�G�join�i�j��oX��ł&cWv	 ���N�v9e��C�clm�&A�o# �|$finde��0STD �ter FiOLANG���R���
��n3��z0Cen���r,������ J����� ���K�〪Ú�=���_Ӛ��r~� "FNDR��� 3��f��tguid�䙃N�."��J�tq�� ��������� ����J����_������c��	m�Z��?\fndr.��n#�>
B2p��Z�CP� Ma�����38PA��� c��6� (�� �N�B�������H 2�$�81��m_���"ex�z5� .Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$�r*$ ��*$r*$%/s#C�d/�.,P�/0*ʲD�PN��$���$*�G}r�$k Exc�'{IF�$MASK�%�93 H5�%H5�58�$548 H��$4-1�$��#1(�$�0 E�$��$-b��$���!UPDT ��B�4�b�4�2�49�0`�4a�3�9j0"M�4<9�4  ��4��4tpsh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4���3adq\�5K�979":E�ajO l "DQ^E^�3�i�Dq ��4ҲO ?R�? ��q�5��T���3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F��t�4��.�5y N� >�2il(in�4��31 JH1�2Q4�2�51ݠ�4rmal� �3)�REo�Z_�� �Ox����4��^F�?onorTf��7_ja�UpZҒ4l�5rmsAU��Kkg���4�$HCd\��fͲ�eڱ�4�REM����4yݱ"u@�RERG5932fO��47Z�>�5lity,�U��8e"Dil\�5�r�o ��7987�?8�25 �3hk910�3 ��FE�0=0P_�Hl\mhm�5� �qe�=$�^�
E��u<�IAymptm�U��BU��vste�y\� 3��me�b�DvI�[�Qu �:F�Ub�*_�
E&,�su��_ E�r��ox���4hu#se�E-�?�sn��������FE��,�box�����c݌,"��� ����z��M��g��pdspw)�	�� 9���b���(��1���c��Y�R��  �>�P���W��������'�0ɵ�[���͂���  �w ,�@� �zA�bumpšuf��B*�Box%��7Aǰ60�BBw���MC� (6�,f�t{ I�s� ST���*��}B�����w��"BBF
�>�`����)��\bbk968 "�4��։�bb�9va69�����etbŠ��X�����ed	�F��1u�f� �sea"������'�\��,���b�ѽ�o6�H�
�	x�$�f���!y����Q[�! tpermr�fd� TPl0~o� Recov,���3D��R642� � 0��C@}s� tN@��(U�rro����yu2r��  ?�
  �����$$CLe� O�������������$z�_DIGsIT��������.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$j����+c:PRODU�CTM�0\PGSTKD��V&ohozf�99��D����$FEAT_I�NDEX��xd���  
��`ILECOMPW ;���#��`��cSETUP2� <�e�b��  N �a�c_�AP2BCK 1�=�i  �)�wh0?{%&c�� ��Q�xe%�I� m���8��\�n� ���!���ȏW��{� �"���F�Տj���w� ��/�ğS������� ��B�T��x������ =�үa������,��� P�߯t������9�ο �o�ϓ�(�:�ɿ^� ��Ϗϸ�G���k�  �ߡ�6���Z�l��� ��ߴ���U���y�� ���D���h��ߌ�� -���Q��������� @�R���v����)��� ��_�����*��N ��r��7�� m�&�3\�i�
pP 2#p�*.VRc�*��� /���PC/1/FR6:/].��/+T�`�/�/F%�/�,�`xr/?�*.F�D8?	H#&?e<�/<�?;STM �2�?н.K �?�=i�Pendant �Panel�?;H �?@O�7.O�?y?�O:GIF�O�O�5�OoO8�O_:JPG _J_��56_�O_�_�	P�ANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEINS.XML���0\���qC�ustom To�olbar	���PASSWORD�yFRS:\�L�� %Pas�sword Config���֏e� Ϗ�B0���T�f��� �������O��s�� ����>�͟b��[��� '���K��򯁯��� :�L�ۯp�����#�5� ʿY��}��$ϳ�H� ׿l�~�Ϣ�1����� g��ϋ� ߯���V��� z�	�s߰�?���c��� 
��.��R�d��߈� ��;�M���q���� ��<���`������%� ��I��������8 ����n���!�� W�{"�F� j|�/�Se ��/�/T/�x/ /�/�/=/�/a/�/? �/,?�/P?�/�/�?? �?9?�?�?o?O�?(O :O�?^O�?�O�O#O�O GO�OkO}O_�O6_�O /_l_�O�__�_�_U_ �_y_o o�_Do�_ho �_	o�o-o�oQo�o�o �o�o@R�ov ��;�_��� *��N��G������ 7�̏ޏm����&�8� Ǐ\�돀��!���E� ڟi�ӟ���4�ßX� j��������įS���w������B�#��$�FILE_DGB�CK 1=���/���� ( �)
SU�MMARY.DG<L���MD:������Diag Summary���Ϊ
CONSLO�G�������D�ӱ�Console �logE�ͫ��MEMCHECK:��!ϯ���X�Mem�ory Data|��ѧ�{)��HADOW�ϣϵ��J���Shado�w Change�sM�'�-��)	FTP7Ϥ�3ߨ����Z�mment� TBD��ѧ0=�4)ETHERNET�������T��ӱEthern�et \�figu?rationU�ؠ~��DCSVRF��p�߽�����%��� verify �all��'�1PY=���DIFF�����[���%��d�iff]������1pR�9�K��� ����X��CHGAD������c��r����2ZAS�� ��GD ���k��z��FY3bI[�� �/"GD ���s/����/�*&UPDATE�S.� �/��FR�S:\�/�-ԱU�pdates L�ist�/��PSRBWLD.CM(?����"<?�/Y�PS�_ROBOWEL ��̯�?�?��?&�O -O�?QO�?uOOnO�O :O�O^O�O_�O)_�O M___�O�__�_�_H_ �_l_o�_�_7o�_[o �_lo�o o�oDo�o�o zo�o3E�oi�o ���R�v� ��A��e�w���� *���я`�������� �O�ޏs������8� ͟\�����'���K� ]�쟁����4���ۯ j������5�įY�� }������B�׿�x� Ϝ�1���*�g����� Ϝ���P���t�	�� ��?���c�u�ߙ�(� ��L߶��߂���(� M���q� ���6��� Z������%���I��� B�����2�����h�����$FILE�_� PR� ���������MDONLY� 1=.�� 
 ���q����� �����~%� I�m�2� �h��!/�./W/ �{/
/�/�/@/�/d/ �/?�//?�/S?e?�/ �??�?<?�?�?r?O �?+O=O�?aO�?�O�O &O�OJO�O�O�O_�O�9_�OF_o_
VIS�BCKL6[*�.VDv_�_.PF�R:\�_�^.P�Vision V?D file�_�O 4oFo\_joT_�oo�o �oSo�owo�oB �of�o�+�� �����+�P�� t������9�Ώ]�� ����(���L�^���� ���5���ܟk� ��� $�6�şZ��~������
MR_GRPw 1>.L���C4  B���	� W������*u���R�HB ��2 ���� ��� ���B�����Z�l��� C���D�������Ŀ���I��9L����J�w�F�5�UT�Q��Ҳ��ֿ Gk�W�E��ED��+-���:���@<W^�@�mA��?f��?n�%A����r��E�� F�@ �������J���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6�\b��B��<%���A�o=�@�0eߋ�NҞ�A��߲� v���r������
�C� .�@�y�d������ ��������?�Z�l�v��BH�� ��R�@(h�E��������
0�PJ��P��V(��ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�OPгߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������>[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U��0
//./A�#��� �~/����/�/�/ �/� ?2?D?V?h?�/ ?�?�?�?�?�?�?� ��@O?dO�/�O�O �O�O�?�O�O__*_ MON_�Or_�_�_�_�_ 	OO-O�_A_&ouOJo \ono�o�o=o�o�o�o �oo�o4FXj |�_�_�_o�7o ��0�B�T�#x��� �������e����� ,�>�����ŏ�� �Ο������:� L�^�p�����'���ʯ ܯ� �O�a�s����� l���������ƿؿ�� ��� �2�D�g��z� �Ϟϰ����#�5�G� I��}�R�d�v߈ߚ� iϾ��������)߫��<�N�`�r��XST_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������O�C�R.RDzVT=#��K@9�BOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ�{
�Å��ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A���   @�<�P�R�
h�BD�b�A��j�����������Dz۩���������j��(� �� -���C���'�7�������Y����� �??�ff ��g|y ������q:a��
>+�  PƱj�(�����7	���|�?˙���xZ�p<
�6b<߈;����<�ê<�? <�&Jσ��AI�ɳ+���?offf?I�?&��k�@�.��J<?�`�q�.� �˴fɺ�/��5/� ���j/U/�/y/�/�/ �/�/�/?�/0?q��F�?l??�?/�?+)�?�?�E��� E�I�G+� F��?)O�?9O_O`JO�OnO�Of�BL޳B�?_h�.��O�O�� %_�OL_�?m_�?�__�_�_�_�_�
�h�yÎg>��_�Co�_goRodo�o�GA�ds�q�C�o�o�o|����$]�Hq���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?��$�?�K�0���
=ç>�����3�W
=�s#�W��e�צ��@����{�����<���(�B�u���=B0�������	L��H��F�G���G���H�U`E����C�+���I�#�I��H�D�F��E��RC�j=���
I��@H��!H�( E?<YD0q� $��H�3�l�W���{� �������՟���2� �V�A�z���w����� ԯ��������R� =�v�a���������� ��߿��<�'�`�K� ��oρϺϥ������ ��&��J�\�G߀�k� �ߏ��߳�������"� �F�1�j�U��y�� ����������0���T�?�Q����(�1�3�3/E�����5�������M3ǭ8�����M4M�gs&IB+�2D�a���{�^^	����(��uP2P7Q4_A��M0bt��R�����,�/   �/� b/P/�/t/�/ *a)_ 3/�/�/�%1a?��/?;?M?_?q?  �?�/�?�?�?�?O~ 2 F�$�v'Gb�/�A��@�a,�`�qC��C@�o�O�2���OF� D�zH@�� F�P D���O�O�ys<O!_3_E_W_i_s�?���@@pZJ.t22!2~
 p_�_�_ �_	oo-o?oQocouo��o�o�o�o��Q ���+��1��$�MSKCFMAP�  �5� �6�Q�Q"~�c�ONREL  �
q3�bEX_CFENB?w
s�1uXqFNC_QtJOGOVLIM?w�dIpMrd�bKEY�?w�u�bRUN�|�u�bSFSPDTY�avJu3s�SIGN?QtT1�MOT�Nq�b_�CE_GRP 1-p�5s\r��� j�����T��⏙�� ����<��`��U��� M���̟��🧟�&� ݟJ��C���7����� ��گ�������4�V��`TCOM_CF/G 1q}�Vp�􂿔�
P�_ARC�_\r
jyUAP�_CPL��ntNO�CHECK ?{ 	r� �1�C�U�g�yϋϝ� ����������	��({�NO_WAIT_�L�	uM�NTX��r{�[m�_ER�RY�2sy3� A&�������r�cx� ��T_MO��}t��, (�$�|k�3�PARAM��u{��V[���!�u?�� =9@345678901� �&���E�W�3�c������{������� �����=�UM_?RSPACE �V�v��$ODRD�SP���jxOFF�SET_CART�ܿ�DIS��PEN_FILE� �q��c֮�OPTI�ON_IO��PWORK v_�ms �P(�R��@�6$j.j	 ��Hj(6$�p=��_DSBL  Ċ5Js�\��RI_ENTTO>p9!sC��Pq=#��UT_SIM_D�
r�b� V� LCT ww�bc���U)+$_PEXE�d&RATp �vju��p��2X�j)TU�X)TX�##X d-�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O?O�H2�/oO�O�O�O��O�O�O�O�O_]�< ^O;_M___q_�_�_�_ �_�_�_�_o���X��OU[�o(�꘯(���$o��, ��IpB` �@D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	l�mb�`�xJ�`�����a�< ��`��m�a, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�b���� �N U�B[�'!o�:q�pC\�C�@@sBq�|���= m�
�A\��h@ߐ�n����Z��B\��A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�����(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��� ��3 ���Ӱ��ɆDT� Qy-����D � ��ӱ4�P :� L :�GP:�D :�@ :�U8�8�	8�
8�U8�8�8�8�Q8�X@:�8�8�8�8�8��:�E8�8�x�:�8�PP�:�d :�8�8�P��:�
�:�!8�"8�Q#8���:�%8�&8�U'8�(8�)8�*8�T��:�,8�-8�.8�/8�08�18�,��� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ��������� � �2�D�V�h�zߌ� �߰���������
�� .�@�R�d�v���� ����������*�<� N�X�(�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_d��_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п�_��� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p�������� //$)�$�PGTRACEL�EN  #!  ��" ��8&_UP z/���g!o S!�h 8!_CFG7 {g%Q#"!�x!�$J �#|"DEFSPD |�,�!!J �8 IN~ TRL }�-�" 8�%�!PE__CONFI� ~g%��g!�$\�%�$LID�#�-�74GRP 1��7Q!�#!A ����&ff"!A�+33D�� D�]� CÀ A)@+6�!�" d�$�9��9*1*0� 	 �+9�(�&�"�? ��	C�?�;B@3AO��?OIO3OmO"!>�?T?�
5�O�O��N�O =��=#�
�O_�O_J_ 5_n_Y_�O}_�_y_�_<�_�_  Dzco" 
oBo�_Roxoco �o�o�o�o�o�o�o�>)bM��;�
V7.10be�ta1�$  �A�E�rӻ�A " �p?!G���q>���r�܁0�q�ͻqBQ��qA\�p�q�4T�q�p�"�BȔ 2�D�V�h�w��p�?�?)2{ȏw�׏ ���4��1�j�U��� y�����֟������ 0��T�?�x�c����� ��ү����!o�,�ۯ P�;�M���q�����ο ���ݿ�(��L�7��p�+9��sF@  �ɣͷϥ�g%����� �+�!6I�[߆����� �ߵߠ���������!� �E�0�B�{�f��� ����������A� ,�e�P���t������� �����=(a L^������ �'9$]�Ϛ� �ϖ�������/ <�5/`�r߄ߖߏ/> �/�/�/�/�/?�/1? ?U?@?R?�?v?�?�? �?�?�?�?O-OOQO <OuO`O�O�O�O�O�� �O_�O)__M_8_q_ \_n_�_�_�_�_�_�_ o�_7oIot���o �o���o�o�o(/! L/^/p/�/{*o�� �������A� ,�e�P�b��������� �Ώ��+�=�(�a� L���p������Oߟ� ��� �9�$�]�H��� l�~�����ۯƯ��� #�No`oro�on��o�o �o�oԿ���8J \ng����vϯϚ� ������	���-��Q� <�u�`�r߫ߖ��ߺ� ������;�M�8�q� \��������z���� ��%��I�4�m�X��� |�����������:� L�^���Z������� ����$�6�H� Swb���� ���//=/(/a/ L/�/p/�/�/�/�/�/ ?�/'??K?]?H?�? ��?�?f?�?�?�?O �?5O OYODO}OhO�O �O�O�O�O�O&8J 4_F_����_�_� �_�_"4-o�O*o coNo�oro�o�o�o�o �o�o)M8q \������� ��7�"�[�m��?�� ��R�Ǐ���֏�!� �E�0�i�T���x��� �����_$_V_ �2��l_~_�_�����R�$�PLID_KNO�W_M  �T������SoV ��U͠�U��
�� .�ǟR�=�O�����m�ӣM_GRP 1���!`0u��T@Rٰo�ҵ�
�� �Pзj��`���!� J�_�W�i�{ύϟϱ����������߱�MR������T��s�w� s��ߠ޴߯߅��� �߻�����A���'� ���������� ����=���#����������}������S��S�T��1 1��U�# ���0�_ A .��,>Pb� �������3 (iL^p��P���2*N���<-/3/)/;/M/4f/x/�/�/5�/�/�/�/A6??(?:?7S?e?w?�?8�?�?�?��?MAD  �d#`PAR�NUM  �w�%OSCH?J �ME
�G`A�Iͣ�EUPD`OrE
a�OT_CMP_��B@�P�@'˥TER_wCHK'U��˪?R$_6[RSl�¯��G_MOA@�_�U_�_~RE_RES_G ��>�oo8o+o \oOo�oso�o�o�o�o��o�o�o�W �\ �_%�Ue Baf�S � ����S0�� ��SR0��#��S�0 >�]�b��S�0}������RV 1�����rB�@c]��t�(�@c\����D�@c[�$���RT?HR_INRl�DA���˥d,�MASS69� ZM�MN8�k��MON_QUEUE ���˦��x�� RDNPUbQN8{�P[��END���_�ڙEXE�ڕ�@B�E�ʟ��OPTI�OǗ�[��PROG�RAM %��%���ۏ�O��TAS�K_IAD0�OCFG ���tO��Š�DATA���Ϋ@��27�>�P�b� t���,�����ɿۿ������#�5�G���IN+FOUӌ������ �ϭϿ��������� +�=�O�a�s߅ߗߩ߀���������^�jč�� yġ?PDI�T �ίc���W�ERFL
��
RGADJ �n�A����?����@�~��IORITY{��QV���MPDSP(H�����Uz����oOTOEy�1�R� (!AF4��E�P]���!t�cph���!u�d��!icm���ݏ6�XY_ȡ�R��ۡ)� a*+/ ۠� W:F�j��� ���%7[�B�*��POR�T#�BC۠�����_CARTRE�P
�R� SKSTyAz��ZSSAV����n�	2500H863���r�$�!�R�����q�n�}/�/�'� UR�GE�B��rYWFF� DO{�rUVWV���$�A�WRUP_�DELAY �|R��$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?�3AQSKIP!�vn�l#x 	1/ +O+ OROdOvO9Hn� �O�G�O�O�O�O�O_ �O_D_V_h_._�_z_ �_�_�_�_�_
o�_.o @oRoovodo�o�o�o �o�o�o�o*<�Lr`���n��?$RCVTM������pDCR!��LЈqC`N��C�d�C��o�?��>��L�<|�{4M�g��&��/����%�t����|��}'�4Oi��O� <
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E0�kATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960�iW+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�M)�$bR  ��ϰ�P{_�P_INTVAL�@�����JR_OPT�ION�V �E�BpVAT_GRPw 2����G(y_Ho �e_ vo�o�oYo�o�o�o�o �o*<�bOoND pw������ 	���?�Q�c�u��� ��/���ϏᏣ���� )�;���_�q������� ��O�ɟ���՟7� I�[�m�/�������ǯ ٯ믁��!�3���C� i�{���O���ÿտ� ��ϡ�/�A�S�e�'� �ϛϭ�oρ������ �+�=���a�s߅�G� �߻����ߡ���'� 9�K�]��߁���� y����������5�G��Y��E�$SCAN�_TIM�AYue�w�R �(�#�((�<0.aWaPaP
T�q>��Q��o������OO"2/���d;2"BaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>HE�̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:L!`O�UT",REC 1�Z� d �  	  	������

 �Z�{0 H6lZ�~�� ���� //D/2/ h/z/\/�/�/�/�/�/ �/�/?�/,?R?@?v? d?�?�?�?�?�?�?�? OO(ONO<OrOTOfO �O�O�O�O�O�O_&_ _J_8_Z_\_n_�_�_ �_�_�_�_�_"ooFo 4oVo|o^o�o�o�o�o �o�o�o0TB xf����(� ��,��P�>�`��� h���������Ώ�� (�:��^�L���p��� ����ܟ���� �6� $�Z�H�~���r����� دƯ����2��&� h�V���z�����Կ� ȿ
�����.�d�R� �Ϛ�|ϾϬ������ ���<��`�N�pߖ� �ߺߨ���������8�&�\�J�l��jV� 1�w Pl��	>� � ��&��
TYPE�VFZN_CF�G �x��d7�GRP� 1�A�c ,�B� A� D;�� B���  B�4RB21^HELL:�(
 X����%RSR���� E0iT�x�� ����/S�ew�����%@w�����#�1����A��2#�d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he�s_ (_:_L_^_��_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}4xcopy �fr:\*.* �virt:\tm�pback�Q=>�192.168.�4�P46:216�4 �R�_�_�_�K}5�Ua�_�_�V�_go�yo�o}9�Ts:o�rderfil.dat.l@oVo�o�o�}0�Rmdb: +o�oRb�ocu�b �_2o?U��
�o���Sod�v����
�xyzrate 61 +�=�O�����������1356 ��ҏc�u����o �o56�ٟ���"���5�џb�t����6ܠ���emp:�60�88 W������.��*.d��Ʈϯ`�r�����1 +�=�O� ����)�Ҳ��ҿ c�uχϚ���5�ͧ�� �����"���̨��b� t߆ߙ����:�V���`��������8 �� g�y��ϰ�9�T��� ��	�߷�@���c�u� ����-�?������� ����N�_q������:L��< ��v792 ��bt�8���* <���/ �� 3�a/s/�/������q534�p�/�/�/ � ��/�(�/`?r?�? ���;?M?�?�?O� '�4�?�?cOuO�O�� �5/�'�O�O�O�"/ �O�(�Ob_t_�_��� �QCU_�_�_
o�_ �_T@�_goyo�o�O�O 9_T_�o�o	_�o@_ �ocu��_-o?o�_ ���o��No_� q����o�o1�oݏ� �&��J[�m������$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1����?���% ֟��&�	��\�?� f���u��������ϯ ��"��F�)�;�|�_� ������ֿ��˿�� �B�%�f�I�[Ϝ�� ���ϵ�������,�� 6�b�E߆�i�{߼ߟ� ����������L�/� V��e������� �����6��+�l�O� v��������������� 2V9K�o ������� &R5vYk�� ���/��<// F/r/U/�/y/�/�/�/ �/?�/&?	??\??? f?�?u?�?�?�?�?�? �?"OOFO)O;O|O_O �O�O�O�O�O�O_�O _B_%_f_I_[_�__ �_�_�_�_�_�_,oo 6oboEo�oio{o�o�o �o�o�o�oL/ V�e����� ���6��+�l�O��v�������PARAoM �����_ �	��P�����OFT_�KB_CFG  �ヱ���PIN_�SIM  ����C�U�g�����RV�QSTP_DSB�,�򂣟����SR� �/�� & �MULTIROBOTTASK������TOP_�ON_ERR  ����PTN� /�@��A	�RING_�PRM� ��V�DT_GRP 1y�ˉ�  	�� ����������Я��� ��*�Q�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߣߠ߲��� ��������0�B�i� f�x���������� ���/�,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZ�~��� ����/ /G/D/ V/h/z/�/�/�/�/�/ �/?
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8___\_��VPRG_COUNT���@���RENB�U��UM�S��__U�PD 1�/�8  
s_�oo*o SoNo`oro�o�o�o�o �o�o�o+&8J sn������ ���"�K�F�X�j� ��������ۏ֏��� #��0�B�k�f�x��� ������ҟ������ C�>�P�b����������ӯί�����UY?SDEBUG�P�P��)�d�YH�SP_�PASS�UB?~Z�LOG ��U+�S)�#�0��  ��Q)�
M�C:\��6���_M�PC���U���Q�ñ8� �Q�SAV �����ǲ&��ηSV;�TE�M_TIME 1���[ (  �w�"����$T1?SVGUNS�P�U�'�U���ASK_OPTION�P��U�Q�Q��BCC�FG ��[u� qn�A�a�`a� gZo��߃ߕ��߹��� ����:�%�^�p�[� ��������� ��� ��6�!�Z�E�~�i���������&������� &8��nY�} �?��ԫ �� (L:p^�� �����/ /6/ $/F/l/Z/�/~/�/�/ �/�/�/�/�/2?8  F?X?v?�?�??�?�? �?�?�?O*O<O
O`O NO�OrO�O�O�O�O�O _�O&__J_8_n_\_ ~_�_�_�_�_�_�_o �_ o"o4ojoXo�oD? �o�o�o�o�oxo .TBx��j� �������,� b�P���t�����Ώ�� ޏ��(��L�:�p� ^�������ʟ��o ��6�H�Z�؟~�l� ������د���ʯ � �D�2�h�V�x�z��� ¿���Կ
���.�� >�d�Rψ�vϬϚ��� ��������*��N�� f�xߖߨߺ�8����� ����8�J�\�*�� n������������ "��F�4�j�X���|� ������������0 @BT�x�d� ����>, Ntb����� �/�(//8/:/L/ �/p/�/�/�/�/�/�/ �/$??H?6?l?Z?�? ~?�?�?�?�?�?O� &O8OVOhOzO�?�O�O �O�O�O�O
__�O@_ ._d_R_�_v_�_�_�_ �_�_o�_*ooNo<o ^o�oro�o�o�o�o�o �o J8n$O �����X����4�"�X�B�v��$�TBCSG_GR�P 2�B���  �v� 
 ?�  �� ����׏�������1���U�g�z���ƈ�_d, ���?v��	 HC��d�>�����e�CL � B���Пܘ������\)��Y�  A�ܟ$�B��g�B�Bl�i�X�������X��  D	 J���r�����C���H��үܬ���D�@v� =�W�j�}�H�Z���ſ@��������v��	V3.00~��	m61c�	*X�P�u�g�pœ>���v�(:�� q��p͟�  O�����p�����z�J�CFG �B�e�� �����������=�� =�c�q�K�qߗ߂߻� ���������'��$� ]�H��l������ ������#��G�2�k� V���z����������� ���p*<N�� �l������ �#5GY}h ����v�b��>� // /V/D/z/h/�/ �/�/�/�/�/�/?
? @?.?d?R?t?v?�?�? �?�?�?O�?*OO:O `ONO�OrO�O�O��O �O�O_&__J_8_n_ \_�_�_�_�_�_�_�_ �_�_oFo4ojo|o�o �oZo�o�o�o�o�o�o B0fT�x� ������,�� P�>�`�b�t�����Ώ �������&�L��O d�v���2�����ȟʟ ܟ� �6�$�Z�l�~� ��N�����دƯ��  �2��B�h�V���z� ����Կ¿����.� �R�@�v�dϚψϪ� �Ͼ�������<�*� L�N�`ߖ߄ߺߨ��� �ߚ�������\�J� ��n��������� �"���2�X�F�|�j� �������������� .TBxf�� �����> ,bP�t��� ��/�(//8/:/ L/�/�ߚ/�/�/h/�/ �/�/$??H?6?l?Z? �?�?�?�?�?�?�?O �?ODOVOhO"O4O�O �O�O�O�O�O
_�O_ @_._d_R_�_v_�_�_ �_�_�_o�_*ooNo <oro`o�o�o�o�o�o �o�o&�/>P�/ ������� ��4�F�X��(��� |�����֏����Ə 0��@�B�T���x��� ��ҟ������,�� P�>�t�b��������� ������:�(�^� L�n�������2d� ����̿�$�Z�H�~� lϢϐ��������Ϻ�  ��0�2�D�zߌߞ� ��j����������
� ,�.�@�v�d���� ����������<�*� `�N���r��������� ����&J\� t��B���� ��F4j|� �^����/��  2 6# �6&J/6"�$TBJ�OP_GRP 2���� � ?�X,i#��p,� �_xJ� �6$��  �< ��� �6$ @�2 �"	 �C��} �&b  Cق'<�!�!>���
55�9>�0+1�33�=�CL� f�ff?+0?�ff�B� J1�%Y?d7�.���/>��2\�)?0�5���;���hCY� � � @� �!B�  �A�P?�?�3EC�  D�!�,�0*B�Oߦ?�3JB��
:���Bl�0���0�$�1�?O6!A�ə�AДC�1D9�G6�=q�E6O�0�p��B�Q�;�A�� �o��@L3D	�@��@__�O�O>B��\JU�OHH�1ts>�A@33@?1� C�� �@�_�_&_8_�>��D�UV_0�xLP�Q30<{�zR� @�0�V�P!o3o�_ <oRifoPo^o�o�o�o Ro�o�o�o�oM( �ol�p~��p4�6&�q5	V�3.00�#m61c�$*(��$1!�6�A� Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,IR�CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;S@�;Q��|8�`�rz@/&�8�6&�<��1�w�^$ESTPARS  *(�{ _#HR��ABL/E 1�p+Z�6#�|�Q� � 1�|�B|�|�5'=!|�	|�E
|�|�˕6!|��|�|���RD	I��z!ʟܟ� ��$���O������¯�ԯ�����S��x#  V���˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������U-���� ĜP�9�K�]�o��-��?�Q�c�u���6�NUoM  �z!� >  Ȑ����_CFG ������!@b IMEBF_TT����x#���a�VER��b�w��a�R 1�p+
 �(3�6"1 ��   6!���������� � 9�$�:�H�Z�l�~��� ������������^$R��_��@x�
b MI_CHANm�� x� kDBGL�V;0o�x�a!n E�THERAD ?U�� �y�$�"�\&n ROUT6��!p*!*~�SNMASK�|x#�255.h��fx^$OOLO_FS_DI��[���	ORQCTRL �p+;/��� /+/=/O/a/s/�/�/ �/�/�/��/�/�/!?���PE_DETA�I��PON_S�VOFF�33P_?MON �H�v��2-9STRTCH/K ���42�VTCOMPAT�a8�24:0FPRO�G %�%M�ULTIROBO�TTO!O06�PL�AY��L:_INSWT_MP GL7�YDUS���?�2LC�K�LPKQUICK�MEt �O�2SCR�E�@�
tps��2�A�@�I���@_Y���9�	SR_GRP 1��_ ���\� l_zZg_�_�_�_�_�_�^�^�oj�Q'ODo /ohoSe��oo�o�o �o�o�o�o!W E{i�������	12345C67��!���X�E�1�V[
 �}�ipnl/a�gen.htmno����𤏶�ȏ~�Pa�nel setup̌}�?��0�B�T�f� ��񏞟�� ԟ���o����@� R�d�v������#�Я �����*���ϯů r���������̿C�� g��&�8�J�\�n�� ���϶���������u� �ϙ�F�X�j�|ߎߠ� ���;�������0��B��*NUALRM�b@G ?��  [������������  ��%�C�I�z�m��������v�SEV  �����t�ECFG Ձ=]/B�aA$   B�/D
 ��/C�W i{�������� PRց;� �To\o�I�6?K0(%����0� ����//;/&/ L/q/\/�/�/�/l�Dc �Q�/I_�@HIST 1ׁ9�  (  ���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1 Ec0p?�?8�?�?/C�� >?P=962n?�?
OO.O�?�?�136c?|O�O �O�OAOSO�?�O__ 0_�O�O_Lu_�_�_�_ :_�/�_�_oo)o;o �__oqo�o�o�o�oHo��o�o%7I~� �a81�ou���� ��o���)�;�M� �q���������ˏZ� l���%�7�I�[�� �������ǟٟh��� �!�3�E�W������ ����ïկ�v��� /�A�S�e�Pb���� ��ѿ������+�=� O�a�s�ϗϩϻ��� ����ߒ�'�9�K�]� o߁�ߥ߷������� �ߎ�#�5�G�Y�k�}� ������������� ��1�C�U�g�y���v� ����������	� ?Qcu��(� ���)�M _q���6�� �//%/�I/[/m/ /�/�/�/D/�/�/�/ ?!?3?�/W?i?{?�? �?�?�����?�?OO /OAOD?eOwO�O�O�O �ONO`O�O__+_=_ O_�Os_�_�_�_�_�_ \_�_oo'o9oKo�_ �_�o�o�o�o�o�ojo �o#5GY�o}�������?���$UI_PANE�DATA 1������?  	�}�0�`B�T�f�x��� )�� ��mt�ۏ����#� 5���Y�@�}���v��� ��ן�������1���U�g�N������ �1��Ïȯگ��� �"�u�F���X�|��� ����Ŀֿ=����� �0�T�;�x�_ϜϮ� ���Ϲ������,ߟ�M��j�o߁ߓߥ� �������`��#�5� G�Y�k��ߏ����� ����������C�*� g�y�`���������F� X�	-?Qc�� ��߫���� ~;"_F�� |�����/� 7/I/0/m/�����/�/ �/�/�/�/P/!?3?� W?i?{?�?�?�??�? �?�?O�?/OOSOeO LO�OpO�O�O�O�O�O _z/�/J?O_a_s_�_ �_�_�O�_@?�_oo 'o9oKo�_oo�oho�o �o�o�o�o�o�o#
 GY@}d��&_ 8_����1�C�� g��_��������ӏ� ��^���?�&�c�u� \�������ϟ���ڟ �)��M������� ����˯ݯ0����� 7�I�[�m�������� ��ٿ�ҿ���3�E� ,�i�Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#� ������ ��$�6�� Z�A�~�e�w����� �������2��V�h��O�����v�p��$U�I_PANELI�NK 1�v��  � � ��}1234567890�� ��	-?G ��� o�����a���#5G�	��h��p&���  R �����Z�� $/6/H/Z/l/~//�/ �/�/�/�/�/�/
?2? D?V?h?z??$?�?�? �?�?�?
O�?.O@ORO dOvO�O O�O�O�O�O �O_�O�O<_N_`_r_�_�_�0,���_�X �_�_�_ o2ooVoho Ko�ooo�o�o�o�o�o �o��,>r}�� �������� ��/�A�S�e�w�� ������я���tv� z����=�O�a�s� ������0S��ӟ��� 	��-���Q�c�u��� ����:�ϯ���� )���M�_�q������� ��H�ݿ���%�7� ƿ[�m�ϑϣϵ�D� �������!�3�Eߴ_ i�{�
�߂����߸� �����/��S�e�H� ���~��R~'�'�a ��:�L�^�p����� ���������� �� 6HZl~��� #�5��� 2D ��hz����� c�
//./@/R/� v/�/�/�/�/�/_/�/ ??*?<?N?`?�/�? �?�?�?�?�?m?OO &O8OJO\O�?�O�O�O �O�O�O�O[�_��4_ F_)_j_|___�_�_�_ �_�_�_o�_0ooTo fo��o��o��o�o �o,>1bt ����K��� �(�:����{O�� ����ʏ܏�uO�$� 6�H�Z�l��������� Ɵ؟����� �2�D� V�h�z�	�����¯ԯ ������.�@�R�d� v��������п��� ϕ�*�<�N�`�rτ� �O�Ϻ�Io������� ��8�J�-�n߀�cߤ� �����߽����o1� �oX��o|������ �������0�B�T� f�������������� S�e�w�,>Pbt ��'���� �:L^p�� #���� //$/ �H/Z/l/~/�/�/1/ �/�/�/�/? ?�/D? V?h?z?�?�?�???�? �?�?
OO.O��ROdO �߈OkO�O�O�O�O�O �O_�O<_N_1_r_�_�g_�_7OM�m��$UI_QUICKMEN  ��_Aob�RESTORE �1�  �|��Rto�o�im�o�o�o�o �o:L^p�% ������o�� ��Z�l�~�����E� Ə؏���� �ÏD� V�h�z���7������� /���
��.�@��d� v�������O�Я��� ��ßͯ7�I���m� ������̿޿���� &�8�J��nπϒϤ� ��a�������Y�"�4� F�X�j�ߎߠ߲��� ���ߋ���0�B�T��gSCRE`?�#mu1sc�o`u2��3��4���5��6��7��8<��bUSERq�v�2��Tp���ks����U4��5��6��7���8��`NDO_C�FG �#k  �n` `PDAT�E ����NonebSEU�FRAME  �TA�n�RTOL_ABRTy�l���ENB����GRP� 1�ci/aCz  A�����Q��  $6HRd���`U�����MS�K  �����N&v�%�U�%����bVISCAND�_MAX�I����FAIL_ISMG� �PݗP#���IMREGNU�M�
,[SIZl�n`�A�,V?ONTMOU���@���2��a��a����FR:\ �� MC:�\�\LOG�B@F� !�'/!�+/O/�Uz �MCV�8#UDM1r&EX{+�S�P>PO64_��0�'fn6PO���LIb�*�#V����,f@�'�/�w =	�(SZV�.w����'WAI�/�STAT ߄���P@/�?�?�:$�?�?��2DWP�  ��P G<@+b=��� H��O_JMPER�R 1�#k
  ��2345678901dF�ψO{O�O �O�O�O�O_�O*__�N_A_S_�_
� ML�OWc>
 �_T�I�=�'MPHASE  ���F��PSHIF�T�1 9�]@<�\�Do�U#oIo�o Yoko�o�o�o�o�o�o �o6lCU� y����� ���	�V�-�e2����	�VSFT1�2	�VM�� �5ԑ1G� ���%Aȯ  B8̀̀�"@ pكӁ˂�у��Fz�ME@�?�{�\�!c>&%�aM1�i�k�0�{ �$`0TDINEND��\�O� �z�����S��w��P���ϜRELE�Q��Y����\�_ACTI�V��:�R�A ���e���e�:�RD�� ���YBOX c�9�د�6��0�2���19o0.0.�83�;�254��QF�	 �X�j���1�rob�ot���   �p�૿�5pc��̿�����7�𼻲�-�f�ZABC
�����,]@U��2ʿ �eϢωϛϭϿ��� �� ���V�=�z�a�Hs߰�E�Z��1�Ѧ