��   D�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b  �CLM�LIy@   $TYPES�INDEXS�$�$CLASS  ����lq�����apVIRTU�ALi{q'61IO�N  �����q�t+ UP�0 �u�qSt�yle Sele?ct 	  ��r��uReq. /E�cho���yAc�k�s�sIni�tiat�p�r�s"�t@�O�a�p���Y	��  ����V;p �����q��������q��sOp�tion bit+ A��B����}C�Decis��cod;��zTry�out mL��Path segJ�_ntin.�II��yc:��Task� OK��!�Man�ual opt.%r�pAԖBޟԖ�C�� decsn� ِ�Robot� interlo��"�>� isol3��C��i/�"�z�ment��z�ِ�����_�statu�s�	MH Fa�ult:��ߧAl�er��%��p@r 1�z L��[��m�+�; LE_CO�MNT ?�y�   ��䆳�Ŀ ֿ�����0�B�T� g�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼������������U������ �  ��ENAB  ���u���������ꐵMEN�U>�y��NAME� ?%��(%$* 4���D��p2�k�V��� z������������� 1U@Rdv� ������ *<u`���� ����/;/&/_/ J/f/n/�/�/�/�/�/ ?�/%??"?4?F?X? j?�?�?�?�?�?�?�? �=