��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ? � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1�� GPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|~GRG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"GSB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3��B�2���AX�D�#
 d �$CARD_E�XIST4$FSSB_TYP~!AHKBD_SNB֒1AGN Gn �$SLOT_N�UM�APREV4DEBU� g1G �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��U0LETE_O�K�BUS�P_CR�A$;4AV� 0/LACIw1�Rp�@k �1$@MEN�@$D�V�Q`Pv�VA{'�BLv� OU&R ,AЧ0�!� B� LM�_O�
eR�"CAsM_;1 xr~$ATTR4��@� ANNN@5I�MG_HEIGH|�AXcWIDTH4�VT� �UU0F_�ASPEC�A$�M�0EXP�.@A�X�f�CF�D ?X $GR� � �S�!.@B�PNFL�I�`�d� UIREx 3T!GITCH+Cj�`N� S�d_LZ`2AC�"�`EDp�dL� J�4S�0� <z�a�!p;G0 �� 
$WARNM�0f�!�@� -s�p�NST� CORN��"a1FLTR{uT�RAT� T}p ? $ACCa1�pp��|{�rORI�Pl�C�kRT0_S~B�\qHG,I1 E[ T�`�"3I�pCTYD�@*2 3`�#@� �!�B*HD�DcJ* Cd�2_�3�_�4_�5_�6_�7�_�8_�94�CO�$ <� �o�op�hK3 1#`O_Mc@�AC t � E�#6NGPvABA � �c1�Q8��`,��@Bnr1�� d�P�0�e�]p� cvnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"Q@�PC�P_*0OFS&R; @� RO_K8T��aIT�3T�NOMI_�0�1p�3�;CP�D �� Ќd@��hPV��mEX�p�� �0g0ۤ�p�r
�$TF�2C$MDM3i�TO�3�0U� ^F� ��Hw2JtC1(�Ez�g0#E�{"F�"F�40CPh@�a2 �@$�P�PU�3N)�ύRևAX�!DU���AI�3BUFp�F��@1 |pp����pPIT� PP�M�M�y��}F�SIMQSI �"ܢVAڤT�	��x' T�`(zM��P��B�qFACTb�@EW�P1�BTvv?�MC� ��$*1JB`p�*1DEC��F��������� �H0CHN�S_EMP1�$G��8��@_4�3�p2|@P��3�TCc�(r /�0-sx��ܐ� MB0i��!����JR� i�_SEGFR��Iv *�aR�TpN�C�ӗPVF4?�bx &��f{uJc !�Ja��� !28�ץ�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb���q@�۽�н����L�83�B���CRC�e�3CCp����c��m cҞb�1J�cѿ�.���*�D$ICb�Cq�5r��ե��@v�'���EVT���zF��_��F,p)N��ܫ�?�4�0A�! �r���h �Ϩ��p�2�͕a��� �د��R�Dx Ϗ��o"27��!ARV�O`C�$L	G�pV�B�1�P��@��t�aA�0'�|�+0Ro�� MEp`"1 �CRA 3 AZ�V�g6p�O �FCCb�`�`F��K������ADI��a�A �bA'�.p��p�`�c¢`S4PƑ�a�AMP$��-`Y�3P�M�]p�UR��QUA1  $.@TITO1/S@S��!����"0�DBP�XWO��B0!5��$SK���2�D�Bq�!"�"�PR�� 
� =����!g# S q1$2�S$z���L�)$�/H���� %�/�$C�!9&?�$ENE�q.c'*?�Ú RE�p�2(H ��O��0#$L|3$$@�#�B[�;���FOs_D��ROSr��#������3RIG7GER�6PApS��>��ETURN�2�c�MR_8�TUw�\�0EWM��M�cGN�P���BLAH��<E���P��&$�P� �'P@T�3�CkD{��DQ���4�1�1��FGO_AWA�Y�BMO�ѱQ#!� CS_�)  �PIS� I gb @{s�C��A��[ �B�$�S��AbP�@�EW�-�TNTVճ�BV �Q[C�(c`�UWr�P��J��P�$0��SAF�E���V_SV�bEOXCLU��n'ONL<зSY�*a�&�OT�a'�HI_�V�4��B���_ #*P0� 9�_z��pg �"�@SG�� +nrr�@6Acc *b��G�#@E�V.iHb>?fANNUN$0.$�fdID�U�2�S�C@�`�i�a��j�f:\�!�pOGI$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6�a�"MS�W�E. 8Q�KE3YI5���TM�10s�qA�vIN��#��"���/ D��HOST_P!�rT��t�a��tn��tsp�pEM�ӰV�����pLc U}LI�0  8	�=ȳ#��!Tk0�!1� � $S��ESAMPL��j�۰f爒�f���I�0��[ $SUB�k�#0�Cp��T�r#a�SAVʅ ��c���C��P�f�P$n0E�w YN�_B#2 0Q�D�I{dlpO(��9#�$�R_I�� �ENC2_S� 3  5�C߰�f�- �SpU����!!4�"g�޲�1T���5X�j`ȷg��0��0K�4�AaŔAV�ER�qĕ9g�DSP�v��PC��r"�(���ƓVALU�ߗHE�ԕM+�I�Pճ��OPP ���TH��֤��P�SH� �۰F��df��J� �q�'T�E�T+6 H�bLL_DUs�~a3@{�0�3:���OTX"����s�"�0NOAUkTO�!7�p$)�H$�*��c4�(�C�%8�C, �"�a&��L�� 8H *8�LH <6����c "�`, `Ĭ�kª�q���q��sq��~q��7*��8��9��0����U1��1̺1ٺ1�U1�1 �1�1ʥ2(�2����2̺2�ٺ2�2�2 �2��2�3(�3��3T��̺3ٺ3�3�U3 �3�3�4(��#�T�?��!9 < �9�&�z��I��1���M��QFE@'@� �: ,6��Q? �@P?9��5�E9�E�@A�b���A�� ;p$TP~�$VARI:��Z���UP2�P< ���TDe���K`�Q�����BAC��"= T�p��e$)�_,�bn�kp+ IFI@G�kp�H  ��P��"F@`�!>t� ;E��sC�ST�D� D���c�<� 	C��{��_����l���R  ���F?ORCEUP?b���FLUS�`H�N�>�F ���RD_CM�@E������ ��@v\MP��REMr F�Q���1k@���7Q
Kr4	NJ�5EFFۓ�:�@IN2Q��OV�O�OVA�	TR3OV���DTՀ�DTMX� ��@ �
ے_PH"p��CL��_TpE�@�p2K	_(�Y_T��v*(��@A;QD� ������!0tܑ0RQ���_�a����M�7�CL�dρR�IV'�{��EAR6ۑIOHPC�@��2��B�B��CM9@����R �GCLF�e!DYk(M�ap#5TuDG��� ��%�aFSSD �s?C P�a�!�1���PQ_�!�(�!1��E�3�!3�+5�&�GR)A��7�@��;�P�W��ONn��EBUG_SD2H�P{�_E A �p|�=��TERM`5�Bi5$Z �OR�I#e0Ci5Y�SM�_�P��e0D�6 ��TA�9E�6 ��UP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1젎4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ3Q�E�p %B`�'EC����@R$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"��A��?���ERV��XQ�Y�� mG>@�BN��U\���R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`� 0SMT6�G�3�GR��13�aPA�L@���`�q�uH �� ���TOC�A�`P	P�`$O�P����p�ѡ�`�0O��RE�`R�4C�AO�p낎Be��`R�Eu�h�A��eo$PWR�IMu��RR_�cN��q=B �I&2H���p_A�DDR��H_LE�NG�B�q�q�q$�Rj��S�JڢSS��SKN��u\��u̳�uFٳSE�A�jrS��[MN�!K���0��b����OLX���p����`ACRO 3pJ�@��X�+��Q���6�OUP3�b_"�IX��a�a1��}� ������(��H��D���ٰ��氋�IO
2S�D�����	�7�L $d��`Y!�_OFFr��PR�M_����HTT�P_+�H:�M (�|pOBJ]"�p��-$��LE~Cd����N � ��֑AKB_�TqᶔS�`lH�LVh�KR"~uHITCOU��[BG�LO�q����h�����`��`S9S� ���HW�#A�:�Oڠ<`INC�PU2VISIO W�͑��n��to��to�~ٲ �IOLN��P 8��R��r��$SLob PU�T_n�$p��P�& ¢��Y F_AS:�"Q��$L�������Q  U�0	P4A0��^���ZPHY��-���/��UOI �#R `�K����$�u�"pPpk����$������0UJ5�S�-���NE6WJOG�KG̲DIS����K�p���#T (�uAV8F�+`�CTR�C
��FLAG2��LG�dU ���؜�13?LG_SIZ����`b�4�a��a�FDl�I`�w� m�_�{0a� ^��cg���4�����������{0��� SCH�_���a7�N�d�V
W���E�"����4�"�UM�Aљ`LJ�@�7DAUf�EAU�p��d|�r�GH�b�����BOO��WL ?�6 IT��y0��REC��SCR� ܓ�D
�\���MARGm�!��զ ���d%�����S����Wp���U� �JGM[��MNCHJ���FN�KEY\�K��PR�G��UF��7P��F�WD��HL��STP��V��=@��А�RS��HO`����C�9T��b ��7�[�U L���6�(RD� ����Gt��@PO������z��MD�FOCU���RGEX��TUI��I��4�@� L�����P����`���P��NE��CAN�A��Bj�VAIL�I�CL !�UDCS�_HII4��s�O��(!�S���S��!��BUFF��!X�?PTH$m���v`��D���AtrY�?P��j�\3��`OS1Z2Z�3Z��� Z � ��[aEȤ��Ȥ�IDX�dPSRrO����zA�STL�R�}�Y&�� Y$E�C���K�&p&�1���![ LQ� �+00�	P���`#qdt�
�U�dw<���_ \ ?�4Г�\���t�#\0C4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#�1D���'B�LD�%�$�%ORGڰ5�2�P VŇVY8�s�T�r�$}d^ ���$6��$�%�S�`T� �B0�4>�6RCLMC�4]?0o?�9�9MI�p}dg_ d=њRQ�=�DSTB�p�c ;F�HHAX�R� JHdLEXCE�Sr1!BM!p�a`� /B�TE��`5a�p=F_A7Ji���KbOtH� K�db q\Q���v$MBC��LI|�)SREQU�IR�R�a.\o�AXD�EBUZ�ALt M��c�b�{P����2�ANDRѧ`�`d0;�2�ȺSDC��N�INl�K�x`��X� �N&��aZ���UP�ST� ezrL�OC�RIrp�E�X<fA�p�9AAOwDAQ��f XY�3OND��"MF,� �f�s"��}%�e/� �v�AFX3@IGG�� g ��t"���ܓs#N�s$R�a% ��iL��hL�v�@�ODATA#?pE��%�tR��Y�Nh �t $MD`qI�}�)nv� ytq�ytH�P`�Pxu��(�zsAN�SW)�yt@��yuD�+�)\b���0o�i -�@CUw�V�p 0�XeRR2��j D�u�{Q��7Bd$CA�LIA@��G��2N��RIN��"�<E�'NTE��Ck�r^��آXb]���_N�ql@k���9�D���Bm��7DIVFDH�@��:�qnI$V,��S�$�����X��o�*����o�H �$BELT|�u!ACCEL�q.�~�=�IRC��� ���D�T�8�$SPS�@�"L�@Ѐr��#^�S�Eы T�P�ATH3���I���3x�p�A_W��ڐ���2nC��4�_MG�$DD��T���$FW�Rp9���I�4��DE7�PP�ABN��ROTS�PEE�[g�� J���[�C@4��@$OUSE_+�VPi�F�SYY���1 q�YN!@A�ǦOF�F�qǡMOU��N�G���OL����INC�tMa6��HB�<�0HBENCS+�8q`9Bp�4�FDm�IN��Ix�]��B��VE���#�y�23_UP�񕋳LOWL� ��p� B���Du�9B #P`�x ���BCv�r��MOSI��BMO�U��@�7PERCH  ȳOV��â
� �����D�ScF� @MP����� Vݡ�@y�j�LUk��Gj�p��UP=ó���ĶTR�K��AYLOA �Qe��A��x�����N`�F�RTI�A$��MOUІ�HB�BS0�p7D5���ë�Z��DUM2ԓS_BCKLSH_Cx� k����ϣ���=���ޡ �	ACLAL�"q��1м@��CH�K� �S�RTY@��^�%E1Qq_�N޴_UM�@�C#���SCL0�r�LM?T_J1_L��9@H�qU�EO�p�b�p_�e�k�e�SPC�0�u���N�PC�N�!Hz \P��C�0~"sXT��CN_:�1N9��I�SF!�?�V���U�/���x�T�2��CB!�SH�:� �E�E1T�T����y����T��PA ��_	P��_� =�����P�!����J6 L�@���OG�G�TO7RQU��ONֹ���E�R��H�E�g_W2���_郅����I�I�I��F�f`xJ�1�~1�VEC3�0BD:B�1p�@SBJRK�F9�0DBL_S�M��2M�P_DL2GRV������fH_��d����COS���LNH������@��!*,�aZ����fMY�_(�T�H��)THET0��NK23���"郶�CB�&CB�C AA�B�"��!��!�&�SB� 2�%GTS�Ar�CIMa������,4#97#$DU ���H\1� �:Bk62�r:AQ(rSf$NE�D��`I��B+5��$̀�!A�%�5�7���LPH�E�2���2SC%C%�2-&PFC0JM&̀V�8V�8T߀LVJV!KV/KUV=KVKKVYKVgIH�8FRM��#X!KUH/KH=KHKKHYKUHgIO�<O�8O�Y�NOJO!KO/KO�=KOKKOYKOM&F��2�!+i%0d�7SP�BALANCE_lo![cLE0H_�%SPc� &�b&�b&PFULC�h�b�gخb%p�1k%�UT�O_��T1T2�i/�2N��"�{�t�#�Ѱ`�0�*�.�T��OÀ<�v INSsEG"�ͱREV4v�Ͱl�DIF�ŕ�1�lzw��1m�0OB0pq�я?�MI{���~nLCHWARY�涢AB��!�$MECH�!o ��q�AX��P����7Ђ�`n 
�d(�U�7ROB��CRr�H�����'�MSK�_f`�p P 
�`_��R/�k�z�����1S�~�|�z�{����z��qINUq�M?TCOM_C� �q  ���pO�?$NOREn��y��pЂr 8p �GRe�uSD�0A�B�$XYZ_�DA�1a���DEBaUUq������s z`�$��COD�� �L���p�$BUFINDX|�w  <�MORm�/t $فUA��ր����r�<��rG���u � $SIMUL  S�*�Y�<̑a�OBJE�`̖�ADJUS�ݐA'Y_IS�D�3�܎��_FI�=��Tu 7�~�6�'��p@} =�C�}p�@b�D���FRIr��T��RIO@ \�E}��y��OPWOYq�v}0Y�SYSBU/@v�$SOPġd����ϪUΫ}pPRUN,����PA��D���r\ɡL�_OUo��q�$)�IMA�G��w��0P_qIM��L�INv�K�?RGOVRDt�梄X�(�P*�J�|��0L�_�`]��0�RB�1�0��M��E�D}��p ��N�PMdֲ��c�w�SL�`�q�w x $OwVSL4vSDI��DEX����#�$��-�V} *�N4�\@#�B�2�G�B�_�M��y�q�E� �x Hw��p��AT+USW���C�0o��s���BTM�ǌ�I
�k�4��x�԰q�y Dw�E&���@E�r��7��жЗ�EXE��ἱ���8��f q�z @w���3UP'��$�pQ�XN����������� �PG΅{ h? $SUB�����0_���!�MPW�AIv�P7ã�LO�R���F\p˕$R�CVFAIL_C���BWD΁�v��DEFSP!p | Lw���Я�\���UNI+�����bH�R�p}_L\pAP��x�t���p�}H��> �*�j�(�s`~�NN�`KETB�%�J�PE Ѓ~��J0SIZE����X�'����S�OR��FORMAT�`��c ��WrEM�t��%�UqX��G��PLI��~p�  $ˀP_SWI�pq�J�_PL��AL_ S�����A��B���� C��D�$E���.�C_�U��� � � ���*�J3K0�����TIA4��5��6��MOM������h���ˀB��AD����������PU� NAR������1H���m��� A$PI�6q��	��� ��K4�)6�U��w|`��SPEEDgPG��������Ի� 4T�� � @��SAMr`��\�]��MOV_�_$�@npt5��5���1���2��������'�2S�Hp�IN�'� @�+����4($<4+T+GAMMWf�1>'�$GET`�p����Da���

pLI�BR>�II2�$H�I=�_g�t��2�&E�;��(A�.� �&LW �-6<�)56�&]��v��p��V��$�PDCK���q��_?�����q�&����7��4���9+� ��$IM_SR��pD�s�rF��r�rL	E���Om0H]��0�-�pq��P~JqUR_SCRN��FA���S_SAV�E_D��dE@�NOa�CAA�b�d@�$q� Z�Iǡs	�I� �J�K � ����H�L��> �"hq������ɢ �� bW^US�A����M4���a�� )q`��3�WW�I@v�_��q�.MUAo�� �� $PY+�3$W�P�vNG�{� �P:��RA��RH��RO�PL�����q� ��sJ'�X;�OI�&�Zxe8 ���m�� p��ˀ�3s�O�O�O�O�Ot�aa�_т� |�� q�d@��.v��.v��d@���[wFv��E���% �-r;B�w�t|�tP���PMA��QUa ��Q�8��1�QTH�H{OLG�QHYS��3ES��qUE�pZB���Oτ�  ـP�ܐ(�A����v�!�t�O`�q��u�"���8FA��IROG�����Q2���o�"��p�^�INFOҁ�׃hV����R���OI���� (�0SLEQ ������Y�3����Á��P0Ow0��5�!E0NU���AUT�A�COPAY�=�/�'��@Mg��N��=�}1������ ���RG��Á���X_�P�$;ख�`
��W��P��@��������EXT_CY�C bHᝡRpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�H�SdB����2�$��F�p���GPLeAdA
�TAR��Б@���P����裔d� ,�0F1L`�o@YN��K��M��Ck��PWR�+�9ᘐ��DELiA}�dY�pAD�a��RQSKIP4�� �A�$�OB`NT2����P_$�M� ƷF@\bIpݷ�ݷ� ݷd����빸��Š��Ҡ�ߠ�9���J2R� ��� 46V�EX� TQQ�� ��TQ������ ��`����RDC�V� �`��X)�R�p������r��m$RGEA�R_� IOBT�2FcLG��fipER��DTC���Ԍ���2T�H2NS}� 1����G T\0 ����u�M\Ѫ`I��d�QREF�1�Á� l�h��ENsAB��cTPE�0 4�]����Y�]��ъQ n#��*��"�������2�Қ�߼���������3�қ'�9�K�]�o��P��4�Ҝ�������������5�ҝ!�3�E�W�i�{�
�6�Ҟ��������(�����7�ҟ-�?Qcu�8�Ҡ��������SWMSKÁ�l��aڝ�EkA/��MO[TE6�����@0�݂TQ�IO}5��ISTP����POW@��� �pJ�����p����E�"$�DSB_SIGN�1UQ�x�C\�TP��/S232���R�i�DEVICEUS��XRSRPARIT|��4!OPBIT�Q�I�OWCONT�R+�TQ��?SRCU�� MpSUXTAS�K�3N�p�0p$TATU�PE#�0������p_XPC)��$FREEFRO�MS	pna�GET\�0��UPD�A�2ΙqRSP� :���� !$US�AN�na&����ER1I�0_�RpRYq5*"�_j@_�Pm1�!�6WRK9KD���6��~QFRIEND�Q��RUFg�҃�0TO�OL�6MY�t$�LENGTH_VT\�FIR�pC�@�ˀE> +IUFINt-RM��RGI�1�ÐAITI�$GX�ñ3IvFG2v7G1`���p3�B�GPR�p�1F�O_n 0��!�RE��p�53҅U�T�C��3A�A�F �G((��":���e1n! ��J�8�%���%]���%�� 74�X TO0�L��T�3H&���8���%b453GE�W$�0�WsR�TD�����T��M����Q�T]�=$V 2����1��а91�8�02�;2
k3�;3�:ifa�9�-i�aQ��NS��ZR$)V��2BVwEV�	V�B;�����&�S��`��F�"�k�@�2a�P5S�E��$r1C���_$Aܠ6wP!R��7vMU�cS�t p'��529�� 0G�DaV`��p�d`���P50�@��-�
25S�/� ��aRW�����B�&�N�AX�!�A:@LAh��r/THIC�1I���X�d1TFEj��q�u�IF_CH�3�qI0܇7�Q�pG1RxV�Ч�]��:�u�_J�F~�PRԀƱ�R�VAT��� �`�`���0RҦ�DOfEΦ�COUԱ��AX�I���OFFSE׆TRIGNS���c@����h�����H�<Y��IGMA0PA��pJ�E�ORG_�UNEV�J� ��S�����d ��$CА�J�GROU����TOށ�!��wDSP��JOGӐL�#��_Pӱ�"O�qp����@�&KEP�#IR��ܔ�@M}R��AP�Q^�Eh0���K�SYS�q"K�PG2�BRK�B��߄�pY�=�d����`�AD������BSO�C���N��DUM�MY14�p@SV��PDE_OP�#S�FSPD_OVR�-���C��ˢΓOIR٧3N]0ڦF�lڦ��OV��SF��p���F+�r!���C�C��1q"LCHDL>��RECOVʤc0���Wq@M������R�O�#��Ȑ_+���s @0�e@VER��$OFSe@CV/ �2WD�}��XZ2���TR�!����E_FDO�MOB_CM���B���BL�bܒ#��adtV@QR�$0p���G$�7�AM5��� eŤ��_M;��"'����8$CA��'�E�8�8$HBK(1����IO<�����QPPA������
��Ŋ�����DVC_DB hC;��#"<Ѝ�r!SՑ1[ڤ�S�3[֪�ATIOq 1q� ʡqU�3���CABŐ �2�CvP��9P^�B����_� �SUBCP	U�ƐS�P �MĀ)0NS�cM�"r�$HW_C��U��S�@��SA�A�pl$U�NITm�l_�AT����e�ƐCYCL�q�NECA���F�LTR_2_FI`O�7(��)&B�LPқ�/�.�_SCT�CF�_`�Fb�l���|�FqS(!E�e�CHA�1���4�D°"3�RSD���$"}����_T�b�PRO����� E%Mi_��a�8!�a� !�a��DI�R0�RAILAC4I�)RMr�LO��C���Qq��#q�դ�+PR=�S�A�p�C/�c 	��FUN9Cq�0rRINP�Q0�0��2�!RAC �B� ��[���[W3ARn���BL�AqA����DA`k�\���LD0 ���Q��qeq��TI"r��K�hPR�IA�!r"AF��P z!=�;��?,`�RK����MǀI�!�DFa_@B�%1n�LM�{FAq@HRDY�4_�P@RS�A�0� >�MULSE@�<��a ��ư�t��m�$�1$��1$1o���߰� x*�EG0wp����!AR���ӆ��09�2,%� 7�A�XE��ROB��WdpA��_l-��SY[�hW!‎&S�'WRU�r/-1��@�STR�������Eb� 	�%��J��AB� ���&X9�����OTo0 ;	$��ARY�s#2h��Ԓ�	ёFI@�~�$LINK|��qC1�a_�#��t�%kqj2XYZ�� t;rq�3�C1j2^8%'0B��'�4����+ �3FI���7�q0����'��_Jˑ��8�O3�QOP_�$;5���ATBA�QB�C��&�DUβ�&6��TURN߁"r�E`11:�p��9GFL�`@_���* �@�5�*7��^Ʊ 1�� KŐ	M��&8���"r��ORQ��a�( @#p=�j�g�#qXU�8����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb��T{� , ��@;�uQ���P\� i��UuQ�We�e�S�ERʑe	��E� O���UdAas��4�S�/7����AX ��B�'q��E1�e�� �i��irp�jJ@�j�@ �j�@�jP�j@ �j�! �f��i��i��i� �i��i�y�y��'y�7yTqHyDEBU8�$32���q`Ͳf2G + AB�����رnSVS�7� 
#�d��L�#�L��1 W��1W�JAW��AW��A W�QW�@!E@?D2.�3LAB�29U4�xAӏ��C # o��ERf�5� � i$�@_ A��!�PO��à�0#�
��_MRAt�� d� � T��ٔER1R����;TY&����I��V�0�cz�TO	Q�d�PL[ �d�"��� ?�w�! � �pp`T)0���_VA1Vr�aӔ����2ٛ!2�E����@�H�E����$W�����V!��$�P��oЩcI��aΣ	 HE�LL_CFG!�� 5��B_BASq�SR3��� a#Sb���U1�%��2��3��U4��5��6��7��8���RO����I0f�0NL�\CAB+�����ACK4������,�\@2@�&�?�_P�U�CO. U�OUG�P~ ����m��������TPհ_KAR��[@_�RE*��P8���|�QUE����uP����CSTOPI_AL7�l�k0��ph��]�l0SEM�d4�(�M4�6�TYN�3SO���DIZ�~�pA�����m_TM�MANRQ��k0E�����$KEYSWITCH���m����HE��BEAT4��|�E- LE~���
��U��F!Ĳ���B�_O_HOM=OG7REFUPPR&��(y!� [�C��O��-�ECOC��Ԯ0_I�OCMWD
�a�p	�m��� � Dh1$���UX���M�β<gPgCFORC���� ��OM.  �� @�5(�U��#P, 1��, 3���45	�NPXw_ASt�� 0���ADD���$S�IZ��$VAR\���TIP/�.�
�A�ҹM�ǐ��/�H1�+ U"S�U!Cz����FRIF��J�S0���5Ԓ�NF�� ܍� � xp`SIƗ�TE�C���CSG%L��TQ2�@&���x�� ��STMT��2,�P �&BWuP���SHOW4���S�V�$�� �Q�A00�@Ma}����� �����&���5���6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G�� 0G���0G���@GP��PG��1	1	U1	1+	18	1E	U2��2��2��2��U2��2��2��2��U2��2��2	2	U2	2+	28	2E	U3��3��3��3��U3��3��3��3��U3��3��3	3	U3	3+	38	3E	U4�4��4��4��U4��4��4��4��U4��4��4	4	U4	4+	48	4E	U5�5��5��5��U5��5��5��5��U5��5��5	5	U5	5+	58	5E	U6�6��6��6��U6��6��6��6��U6��6��6	6	U6	6+	68	6E	U7�7��7��7��U7��7��7��7��U7��7��7	7	U7	7+	78	7Ev��VP��UPDs��  �`NЦ��
�SYSLO>t�� � L��0d���A�aTA�0d��|�ALU:ed�~��CUѰjgF!aID�_L�ÑeHI�jI~��$FILE_����d��$2�
�cS�A>�� hO��`E_BLCK��b$�>�hD_CPUyM� yA��c�o�d�b�����R �Đ
PWl��!� oqLA���S=�ts�q~tRUN �qst�q~t���q�st�q~t �T��A�CCs��X ;-$�qLEN;��t�H��ph�_�I��ǀL�OW_AXI�F)1�q�d2*�MZ���ă��W�Im�ւ�aR�GTOR��pg�D�<Y���LACEk�ւp�pV�ւ~�_MA2�pv�������TCV��؁��T��ي����� t�V����V�Jj�R��MA���J��m�u�b����q2j�#�U��{�t�K�JK��VK�;���H���3��J0l����JJ��JJ��AAL��ڐ��ڐԖe4Օ5���N1��P�ʋƀW�LP�_(��g����pr�� =`�`GROUw`����B��NFLIC���f�REQUIRE3�EBU��qB���w�2����p���q�5�p�� \��A�PPR��C}�Y�
vްEN٨CLO7��S_M��H���u�y
�qu�� �`��MC�����9�_M	G��C�Co��`M��ܲ�N�BRKL�NO�L|�N�[�R��_L!INђ�|�=�J����Pܔ������������������6ɵ�̲8�k�+��q���� ��
��q)��7�PATH3�L�B�L���H�wࡠ�J�CN��CA�Ғ�ڢB�I�N�rUCV�4a��C!�UM��Y,�����aE�p����ʴ���PAYLOA��J{2L`R_AN�q�Lpp���$�M��R_F2LSHR��N�LOԡ�Rׯ�|`ׯ�ACRL_G� �ŒЛ� ��Hj`߂�$HM���FLE�Xܣ�qJ�u� :��������������1�F1 �V�j�@�R�d�v�������E����ȏڏ� ���"�4�q���6�M� ��~��U�g�y�ယ	T��o�X��H����� �藕?�����ǟِ ݕ�ԕ����%�7���JJ�� � `V�h�z���`AT��l��@�EL�� Sj��J|�Ŝ�JEy�gCTR��~�TN���FQ��HAND_�VB-���v`�� $��F2M�����ebSW�q�'���� $$MF�:�R g�(x�,4�%��0&�A�`�=��aM)F�A(W�Z`i�Aw�A��X �X�'pi�Dw�D��P2f�G�p�)STk��!4x��!N��DY�pנ M�9$`%Ц�H��H׀c�׎���0� ��P ѵڵ������������ ���1���R�6��QASYM$vř���v��J���cі�_SH>��Ǻ� ��ED����������J�İ%��C�IDِ�_VI�!X�2PV_UNIX�FThP�J��_R�5_Rc�cT z�pT�V��@���İ��ȷ��U ���Ӥ'��T��Hqpˢ���aEN�3�D	I����O4d�`J��� x g"IJAA ȱz�aabp�coc�`a��pdq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a��iT�@<� $�DUMMY9Q�o$PS_��RFC�s  S�v �p8���Pa� XƠ����STE���SB}RY�M21_VF�8$SV_ERF�qO��LsdsCLRJtEA��Odb`O�p� � D $�GLOBj�_LO ���u�q�cAp�r�@awSYS�qADR`�`�`TCH  �� ,��ɩb�W_NA���7���SR���l ���
*?�&Q�0" ?�;'?�I)?�Y)��X� ��h���x������)�� Ռ�Ӷ�;��Ív�?���O�O�O�D�XSCSRE栘p����3ST��s}y`�����/_HAΗq� TơgpTYP�b���G�aG�j��Od0IS_�䓀d�UEMd�# ����ppS�qa�RSM_�q*eUNEXCEP)fW�`S_}pM�x���g�z�8����ӑCOU��S��Ԕ 1�!�UE�&��Ubwr��PRO�GM�FL@$CUgpPO�Q��5��I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp��OUS�� �� @6p�v$BU�TTp�RpR�CO�LUMq�e��SE�RV5�PANE|H�q� � �@'GEU���Fy��?)$HELPõ)B/ETERv�)ෆ� ��A � ��0`��0��0ҰIN簊�c�@N��IH�1��_� �v��LN�r� �qprձ_ò=�$H���TEXl����F�LA@��RELVB��D`��������M��?,�ű�m�����"�USRVwIEW�q� <6p�`U�`�NFI<@;�FOCU��;�7PRI� m�`�Q�Y�TRIP�qm��UN<`Md� x#@p�*eWARN)e�6�SRTOL%���g��ᴰONCOR�N��RAU����T����w�VIN�Le�� $גPA�TH9�גCACH���LOG�!�LI�MKR����v���HwOST�!�bz�R��OBOT��d�IM>� �� ����Zq�Zq;�V�CPU_AVAIYL�!�EX	�!AN���q��1r��1r���1 �ѡ�p� � #`C����@$�TOOL�$��_wJMP� ���e$SS���Ea�VSHIF��Nc߃P�`ג�E�ȐR�����OSUR��Wk`RADILѮ��_�a��:�9a��`a�r���LULQ$OUTPUT_BM����IM�AB �@�r�TILSCO��C7����� ��&��3��A��@�q���m�I�2G���1V�pLe�}��yD�JU��N�WA�IT֖�}��{�%�! NE�u�YBO��� �� �$`�t�SB@T;PE��NECp�Jp^FY�nB_T��R�І�a$�[Yĭc	B��dM���F� `�p�$�pb�OP?�wMAS�_DO�!QT�pD��ˑ#�%��p!"DELAY�:`7"JOY�@(� nCE$��3@ �xm��d�pY_[�!"�`�"��[���P? ��1ZABC%�� � $�"R��
�ϐ�$$CLAS>������!pxE`� � VIRT]ќ�/ 0ABS����1� 5� < �! F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $�6HZi{0-�AX�L�p��"�63  ��{tIN��qztP#RE�����v�p�u�LARMRECO�V 9�rwtN�G�� .;	 �A   �.�0PoPLIC��?5��p�Ha�ndlingTo�ol o� 
V�7.50P/23~-�  �Pf���
��_SWt� �UP�!� x�F�0��t���A0v�� 864�� �it�y� r�2 7D�A5�� �� �Qf@��o�Ngoneisͅ˰ ��T���!�LAex>�_�l�V�uT��s9�U�TO�"�Њt�y��HGAPON
0g�1z��Uh�D 1581����̟ޟxry����Q 1���p�,�蘦����;�@��q_��"=2 �c�.��H���D�HTTHKYX��"�-� ?�Q���ɯۯ5���� #�A�G�Y�k�}����� ��ſ׿1�����=� C�U�g�yϋϝϯ��� ��-���	��9�?�Q� c�u߇ߙ߽߫���)� ����5�;�M�_�q� �������%���� �1�7�I�[�m���� ������!����- 3EWi{��� ���)/A Sew����/ ��/%/+/=/O/a/ s/�/�/�/�/?�/�/ ?!?'?9?K?]?o?�? �?�?�?O�?�?�?O#O]���TO�E�W��DO_CLEAN���7��CNM  � �__/_�A_S_�DSPDR3YR�O��HIc��M@�O�_�_�_�_oo +o=oOoaoso�o�o���pB��v �u���a�X�t������9�PL�UGG���G��U�P�RCvPB�@���_�orOr_7�SEGF}�K[mwxq �O�O�����?rqLAP�_�~q�[� m��������Ǐُ�����!�3�x�TOT�AL�f yx�USE+NU�p�� �H����B��RG_STR�ING 1u�
_�Mn�S5��
ȑ_ITEM1Җ  n5�� � �$�6�H�Z�l�~��� ����Ưد���� ��2�D�I/O �SIGNAL̕�Tryout �ModeӕIn�p��Simula�tedבOut���OVERR~�P = 100֒�In cycl���בProg OAbor��ב���StatusՓ	�Heartbea�tїMH Fa�ul��Aler '�W�E�W�i�{ύϟ�p�������� �C Λ�A����8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|���WOR{pΛ��(ߎ� ���� ��$�6�H�Z� l�~�������������p�� 2PƠ �X ��A{��� ����/A Sew�����SDEV[�o� #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1?�C?U?g?y?PALTݠ1��z?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_�?GRI�`ΛDQ�? _l_~_�_�_�_�_�_ �_�_o o2oDoVoho@zo�o�o�o2_l�R� �a\_�o"4FX j|����������0�B�T��oPREG�>�� f��� Ə؏���� �2�D� V�h�z�������ԟ����Z��$ARG�_��D ?	����;��  	$Z�W	[O�]O��Z��p�.�SBN_CONFIG ;�ꎱ����CII�_SAVE  �Z�����.�TCE�LLSETUP �;�%HOM�E_IOZ�Z�%�MOV_��
�R�EP�lU�(�UTOoBACKܠ���FRA:\�z� \�z�Ǡ'�`�z���ǡi�I�NI�0z���~n�MESSAG����ǡC���ODE_!D������%�O�4��n�PAUSX!�~;� ((O>� �ϞˈϾϬ������ ����*�`�N߄�r��߶�g�l TSK � wͥ�_�q�UP3DT+��d!�AſWSM_CF���;���'�-�GRgP 2:�?� N��BŰA��%�XSC�RD1�1
7� 	�ĥĢ�������� ��*�������r��� ��������7���[� &8J\n��*�>t�GROUN�UϾ�UP_NA��:�	t��_ED��17�
 �%�-BCKEDT�-�2�'K�`D���-t�z�q�Yq�z���2t1�����q�k�8(/��ED3/���/�.a/�/;/M/ED4�/t/)?�/.?8p?�/�/ED5`??��?<?.�?O�?�?ED6O�?qO�?.MO8�O'O9OED7�O`O�_�O.�O\_�O�OE�D8L_,�_�^�-�_ oo_�_ED9�_�_]o�_	-9o�oo%oCR_ �9]�oF�o�k� � N�O_DEL��GE_UNUSE���LAL_OUT� ����WD_ABORﰨ~���pITR_RTNz��|NONSk����˥CAM_�PARAM 1�;�!�
 8
S�ONY XC-5�6 234567w890 ਡ�@���?��( А\�
���{�u���^�HR5q�8̹��ŏR57ڏ��Aff��KO�WA SC310�M
�x�̆�d @<�
���e� ^��П\����*��<��`�r�g�CE__RIA_I�!�5=�F��}�z�� ��_LIU��]�����<��F�B�GP 1��Ǯ�M�_�q�0��C*  ����C1*��9��@��G����CR�C]��d��l���s��R�����[�Դm��v���������� C����b(�����=�HE�`�ONFIǰ�B�G_PRI 1�{V���ߖϨϺ�����������CHKPwAUS�� 1K� ,!uD�V�@�z� dߞ߈ߚ��߾����� �.��R�<�b��ҍO��������_�MOR�� �<6��� 	 ��� ��*��N�<����䡑��?��q?;�;�����K��9�P��|�ça�-:���	�

��M��@�pU�ð��<��,~���DB���튒)�
mc:cpmi�dbg�f�:����u�	p�/�&�H�
� �,s>܋�Q��?��g(�/��f�M/�w�O/�
DEF �l��s)�< b?uf.txts/��t/��ާ�)�	`z�����=L���*[MC��1����X?43��1��t�~īCz  BHH�ދ�B�$�y6��y��.�4D��Y�D���/�4E�CeYF��Y��,�'w�1���s�U��.�p�����1�BDw�M@x8�K�cCҨ��0fADȷ0�0E��8EX��EQ�EJP �F�E�F� �G��=F^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE d��
Q��;�(PG  B_<_��R�����	op6C4P�Y
s@ ]AQ�2s@�C�0B3�MaC�@�*cw��UT�pFP?ROG %�z�o�oigI�q���v��ld�KEY_TBL � �&S�#� �	
��� !"�#$%&'()*+,-./01i��:;<=>?@A�BC� GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������vq���͓���������������������������������耇����������������������p`LCK�l4�p`��`STAT ��S_AUTO_DO����5�INDT_'ENB!���R�Q?��1�T2}�^�STO�Pb���TRLr`L�ETE��Ċ_S�CREEN ~�Zkcsc���U��MMENU �1 �Y  <�l�oR�Y1�[��� v�m���̟�����ٟ �8��!�G���W�i� �������ïկ��4� ��j�A�S���w��� ��迿�ѿ����T� +�=�cϜ�sυ��ϩ� ��������P�'�9� ��]�o߼ߓߥ���� ����:��#�p�G�Y� ����������$� ���3�l�C�U���y� ���������� ��	�VY)�_MANU�AL��t�DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[/ , 
�odP�&/~&lMZ�IdP�x@P@#ONTImMه� d�`&�
�e�MOTN�END�o�REC�ORD 1(�[8g2�/{�O��!�/ ky"?4?F?X?�(`? �?�/�??�?�?�?�? �?)O�?MO�?qO�O�O �OBO�O:O�O^O_%_ 7_I_�Om_�O�_ _�_ �_�_�_Z_o~_3o�_ Woio{o�o�_�o o�o Do�o/�oS�o L�o����@� ��+�yV,�c�u� �������Ϗ>�P�� ���;�&���q���� ����P�ȟ�^���� ��I�[����� ����$�6�������jTOLERENCwsB���L�͖ �CS_CFG �)�/'dMC�:\U�L%04dO.CSV�� c���/#A ��CH��z� //.ɿ��(S��RC_OUT �*���SGN� +��"��#��27-JAN-�20 21:53�015l�10:5�1+ P/V�t�ɞ�/.��f�p�a�m��PJ�PѲ��VERS�ION Y�V2.0.84,�EFLOGIC {1,� 	:�ޠ=�ޠL��PR?OG_ENB��".p�ULSk' �����_WRSTJN�K ��"fEMO_�OPT_SL ?�	�#
 	R575/#=������0�B����TO � �ݵϗ��V_VF EX�d�%��PATH AYʇA\�����5+IkCT�Fu-��j�#eg�S�,�STBF_TTS�(�	d���l#!:w�� MAU��z�.^"MSWX�.��Q4,#�Y�/�
!J �6%ZI~m���$SBL_FA�UL(�0�9'TD�IA[�1<�� ����1234?567890
��P��HZl~� ������/ /@2/D/V/h/�� P� ѩ�yƽ/�� 6�/�/�/??/?A? S?e?w?�?�?�?�?�?p�?�?�,/�UMP��f�� �ATR��8��1OC@PMEl�OO�Y_TEMP?�Ç��3F���G�|DU�NI��.�YN_B�RK 2_�/�E�MGDI_STA���]��ENC2_S_CR 3�K7 (_:_L_^_l&_�_�_`�_�_)��C�A14_ �/oo/oAoԢ�B�T5�K�ϋo~o l�{_�o�o�o' 9K]o���� �����#�5��/ V�h�z��л`~����� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T��� x���������ү��� ��,�>�P�b�t��� ������ο���� (�f�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������:� �2�D�V� h�z���������� ��
��.�@�R�d�v� ������������� *<N`r�� �����& 8J\n����� �����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?��?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__�NoETMODE �16�5�Q �d�X
X_j_|Q��PRROR_PR�OG %GZ%��@��_  �UTAB_LE  G[�?�oo)oRjRRSE�V_NUM  <�`WP�QQY`��Q_AUTO_ENB  �eOS�Tw_NOna 7G[��QXb  *�*�`��`��`��`d`�+�`�o�o�o�dHI�SUc�QOP�k_AL�M 18G[ �2A��l�P+�ok@}�����o_Nb.�`  G[�a�R�
�:PTCP_VE/R !GZ!�_��$EXTLOG_7REQv�i\��SIZe�W�TOL�  �QDzr��A W�_BWD��p��xf́t�_DIn�� 9�5�d��T�QsRֆSTEP���:P�OP_D�Ov�f�PFAC�TORY_TUN�wdM�EATUROE :�5̀rQ�Handl�ingTool ��� \sfm�English �Dictiona�ry��roduAA Vis�� Master��ީ�
EN̐nalog I/O��ީ�g.fd̐ut�o Softwa�re Update  F OR��matic Ba�ckup��H59�6,�ground Editޒ�  1 H5�Camera�F���OPLGX�elyl𜩐II) X�7ommՐshw���7com��co����\tp���pan}e��  opl���tyle sel�ect��al C�nJ�Ցonit;or��RDE���tr��Relia�b𠧒6U�Dia�gnos(�푥�5�528�u��he�ck Safet�y UIF��En�hanced Rob Serv%��q ) "S�r�U?ser Fr[������a��xt. D�IO �fiG� �sŢ��endx�Ekrr�LF� pȐ�ĳr됮� ���� � !��FCTN /Menu`�v-�ݡ|���TP Inې�fac�  ER_ JGC�pב_k Exct�g���H558��igh�-Spex�Ski~1�  2
P���?���mmunic�'�ons��&�l�uqr�ې��ST Ǡ���conn��2ި�TXPL��nc=r�stru�����"FATKA�REL Cmd.� LE�uaG�54�5\��Run-T�i��Env��d�
!���ؠ++�s�)�S/W��[�LicenseZ��� 4T�0�ogB�ook(Syڐm�)��H54O�MA�CROs,\�/O�ffse��Loa��MH������r,� k�MechStop Prot����� lic/�MiвShif����ɒ�Mixx��)���x�StS�Mode �Switch�� �R5W�Mo�:�.�� 74 ����g��K�2h�ult�i-T=�M���LN (Pos�Regiڑ������|d�ݐt Fun��⩐.�����Numx~����� lne�|�ᝰ Adjup������  - W���tatuw᧒T��RDMz�o}t��scove U�9���3Ѓ�uest 492�b*�o�����62;�?SNPX b ����8 J7`���Li3br��J�48����"�� �Ԅ�
�6O��� Parts i�n VCCMt�3�2���	�{Ѥ�J9�90��/I� 2� P��TMILI�B��H���P�A�ccD�L�
TE�$TX�ۨ�ap1�S�Te����pke�y��wգ�d���Unexcep=tx�motnZ���������є�� qO���� 90J��єSP CSXC`<�f��Ҟ� Py�sWe}���PRI��>vr�t�menz�� ��iPɰ�a�����vGri=d�play��v���0�)�H1�M-�10iA(B20�1 �2\� 0\}k/�Ascii��l�Т�ɐ/�Col���ԑGuar� �
�� /P-�ޠ"Kv��st{Pat �:�!S�Cyc��΂�orie��IFn8�ata- quҐ��� ƶ��mH57m4��RL��am����Pb�HMI D�e3�(b����PC�Ϻ�Passwo�+!��"PE? Sp�$�[���tp��� vKen��Tw�N�p��YELLOW B�OE	k$Arc��v�is��3*�n0W�eldW�cialh�7�V#t�Op�����1y� 2F�a�portN�(�p�T1�T� �� �ѳxy]�&TX��t�w�igj�1� b� �ct\�JPN �ARCPSU P�R��oݲOL� S;up�2fil� &�PAɰאcro�� �"PM(����O$SuS� eвtex�ԣ r���=�t�s'sagT��P���P@�Ȱ�锱�rt�W��H'>r�dpn��n1
t�!�� z ��ascbi?n4psyn��+A}j�M HEL��NCL VIS �PKGS PLOA`�MB �,�4�VW�RIPE �GET_VAR {FIE 3\t���FL[�OOL: �ADD R729.FD \j8'�iCsQ�QE��DVvQ��sQNO WTW�TE��}PD  ��^��biRFOR ���ECTn�`��ALSE ALAfP�CPMO-130�  M" #h�D�: HANG F�ROMmP�AQfr���R709 DR�AM AVAIL?CHECKSO!���sQVPCS SU��@LIMCHK �Q +P~dFF PO�S��F�Q R59�38-12 �CHARY�0�PR�OGRA W�SwAVEN`AME�P�.SV��7��$E�n*��p?FU�{�TR}C|� SHADV0�UPDAT KC|JўRSTATI�`~�P MUCH y��1��IMQ MO?TN-003��}��ROBOGUIDE DAUGH�a8���*�tou�����I� Šhd�ATH|�PepMOVET��ǔVMXPACK� MAY ASS�ERT�D��YCL�fqTA�rBE C�OR vr*Q3rA�N�pRC OPToIONSJ1vr̐PSH-171Z@-x�tcǠSU1�1`Hp^9R!�Q�`_T�P���'�j�d{tb�y app wac 5I�~d�PHI����p�aTEL�MX?SPD TB5bLu� 1��UB6@�qEN�J`CE2�61��p���s	�may n��0� R6{�R� >�Rtraff)��� 40*�p��fr���sysvar ?scr J7��cNj`DJU��bH �V��Q/�PSET �ERR`J` 68���PNDANT �SCREEN U�NREA��'�J`D��pPA���pR`IgO 1���PFI�p}B�pGROUN�P�D��G��R�P�QnRS�VIP !p�a�PD�IGIT VER�S�r}BLo�UEW~ϕ P06  �!��MAGp�abZV��DI�`� SS�UE�ܰ�EPL�AN JOT` D�EL�pݡ#Z�@D�͐CALLOb�Q �ph��R�QIPN�D��IMG�R7{19��MNT/�PWES �pVL�c���Hol�0Cq���tP�G:�`C�M�caynΠ��pg.v�S�: 3D mK�v_iew d�` �p���ea7У�b� o�f �Py���ANN�OT ACCESGS M��Ɓ*�t47s a��lok��Flex/:�Rw�!mo?�PA?�-�����`n�pa S�NBPJ AUTO-�06f����TB���PIABLE1q �636��PLN:Y RG$�pl;pNW7FMDB�VI���t�WIT 9x�0@o���Qui#0�ҺPN� RRS?pUSB��� t & remov�@ )�_��&�AxEPFT_=� �7<`�pP:�OS�-144 ��h qs�g��@OST� �� CRASH �DU 9��$�P�pW� .$��L/OGIN��8&�J���6b046 issue 6 Jg���: Slow ��st��c (HCos`�c���`IL`�IMPRWtSPO�T:Wh:0�T�S�TYW ./�VMGqR�h�T0CAT��hos��E�q���� �O�S:+pRSTU' k�-S� ����E:��pv@�2�N� t\hߐ��m ���all��0�  �$�H� WA͐��3 CNT0 T��� WroU�alacrm���0s�d � @�0SE1���r R{�OMEBp���K� �55��REàSEs�t��g    } �KANJI��no���INIS?ITALIZ-p�d�n1weρ<��dr�� lx`�SCI�I L�fail�s w�� ��`�YSTEa���o��PvЧ IIH���1W�G�ro>Pm ol\�wpSh@�P��Ϡn� cflxL@АW{RI �OF Lq���p?�F�up��d�e-rela�d� "APo SY�c}h�Abetwe:0IND t0$gb#DO���r� `��GigE�#ope�rabilf  P�AbHi�H`��c�le{ad�\etf�P8s�r�OS 030��&: fig��GL�A )P ��i��7�Np tpswx�B��If�g�������5aE�a EXC�E#dU�_�tPCLO�S��"rob�NTdpFaU�c�!����PNIO V750�Q1��Qa��'DB ��P M�+Pv�QED�DET���-� \rk��ON�LINEhSBUG�IQ ߔĠi`Z�IB�S apABC �JARKYFq� ����0MIL�`� R��pNД �p0GAR��D*pR��P�"'! jK�0cT�P��Hl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P��`WIBPK05��!FȐB/��BUSY RUNN��C "�򁐈��R-p��LO�N�DIV�Y�CUL��fsfoaBW�p����30	V��ˠIT�`�a505.�@O=F�UNEX�P1bҬaf�@�E��SVwEMG� NMLq�� D0pCC_SA�FEX 0c�08"qD. �PET�`N@�#'J87����RsP�TA'�M�K�`K��H GUNCHG^۔MECH�pMcz� T�  y, g@��$ ORY LE�AKA�;�ޢSP�Em�Ja��V�tGR�Iܱ�@�CTLN�TRk�FpepR��j50�EN-`IN�����p �`�Ǒ�k!��T3/dqo�SKTO�0A�#�L�pA �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`D	U��aO�supk�t4� � P�F� Bnf��Q�PSVGN-18��V�SRSR)J�UP�a2�Q�#D�q� l O��QBRKCTR5Ұ�|"-��r�<pc�j!INVP�D ZO� ��T`�h#�Q�cHset,x|D��"DUAL� �w�2*BRVO117 A]�TNѫt�+bTa2473��q.?���sAUz�i�B�complete���604.� -^�`hanc�U�� F��e8��  ��npJtPd!q��`��w� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP��R�R(}\xPe� aʰ�I���E��1��p�� j  �� xSt�^t �A�AxP�q �5 sig��a��"AC;a��
�bCe�xPb_p��.pc�]l<bHbcb_cicrc~h<n�`tl1� ~`xP`o�dxP�b]o2�� �cb�c�ixP�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`�cptlibxzxP�l�cr�xrxP\�blpsazEdxP_fm�} gcxP�x���o|sp�or�mc(��ob_jzo"p�u6�wf��t���wms�1q��sld�)��jmc�o\�n�b�nuhЕ��|st�e���>�pl�qp�iwc1k���uvf0uߒ<��lvisn�CgoaculwQ
E �F  ! Fc.f9d�Qv�� qw����Data Acq/uisi��nF�|1��RR631`��TR��QDMCM �2֝P75H�1�P58�3xP1��71��559`�5�P57<PxP�Q����(���Q���o pxP!daq�\�oA��@�� �ge/�etdms�"�DMER"؟,�p#gdD���.�m���-��qaq.<᡾xP#mo��h���f{�u��`13��MACRO�s, SksaffP�@z����03�SR�QT(��Q6��1�Q9ӡ��R�ZSh��PxPJ6+43�@7ؠ6�P�@�PRS�@���e �Q��UС PIK�Q5?2 PTLC�W���xP3 (��p/O ��!�Pn �xP5���03\sfmn�mc "MNMCPq�<��Q��\$AcX�FM���ci,Ҥ�X�����cdpq+�
�sk��SK�xP�SH5�60,P��,�y�r�efp "REF�p�d�A�jxP	�of��OFc�<gy�to��TO_����ٺ����+je�u��caxis2�xPE�\�}e�q"ISDTc�|�]�prax ���MN��u�b�is�de܃h�\�w�xP!� isbasic���B� P]��QA7xes�R6�������.�(Ba�Q�ess��xP���2�pD�@�z�atis�� ��(�{�����~��m��FMc�u�{�
���MNIS��ݝ�� ��x����ٺ��x�� j75��Dev�ic�� Inte�rfac�RȔQJ�754��� xP�Ne`��xP�ϐ2��б����dn� "�DNE���
tpodnui5UI��ݝ	bd�bP�q_rsofOb
?dv_aro��u�����stchkc��z	 �(}�onl��G!ff L+H�J(��"l"/��n�b��z�haSmp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!2���xpc_2pcch=m��CHMP_�|8бpevws��2�ΌpcsF��#C �SenxPacro0�U·�-�R6�Pd�@xPk�����p��gT�L��1d M�2`��8��1c4ԡ�3 qem��GEM,\i(��Dgesnd�5���H0{�}Ha�@sy���c��Isu�xD��Fmd ��I��7�4���u���AccuCal�P��4� ��ɢ7ޠB0���6+6f�6��9!9\aFF q�S(�U��2�
X�p�!Bd�ѳcb_�SaUL�� � �� ?�ܖto���otplus\tsrnغ�qb�W�p��t���1��To�ol (N. A�.)�[K�7�Z�(P��m����bfclls� k94�"K4p���qtpap� �"PS9H�stpswo��p�L7��t\�q����D�yt5� 4�q��w�q��� �Mz�uk��rkey�����s��}t�sfe7atu6�EA��� cf)t\Xq�����df�h5���LRC0�md�!�587���a�R�(����2V��8lc?u3l\�pa3}@H�&r-�Xu���t,�� �q "�q�Ot��~ ,���{�/��1c�}����y�p�r��5����S�XAg�-�y���Wj�874�- iR�Vis���Queu�� Ƒ�-�6�1$���(����u����tӑ����
�tpv�tsn "VTS�N�3C�+�� v\pR�DV����*�prd�q\�Q�&�vst�k=P������nmx&_�դ�clrqν���get�TX��Bd���aoQϿ�0q�str�D[� ��t0�p'Z����npv��@�enlIP0��D!0x�'�|���sc ߸��tvo/��2�q���vb����q����!���h]��(� Control�PRAX�P5��5�56�A@59�P5-6.@56@5A��J69$@982 �J552 IDVR7�hqA���16�Hx���La�� ���Xe�frlparwm.f�FRL��am��C9�@(F �����w6{���A���QJ643�� 5}0�0LSE
_p�VAR $SGS�YSC��RS_UNITS �P�2�4�tA�TX.$VN�UM_OLD 5`�1�xP{�50+��"�` Funct ���5tA� }��`#@�`E3�a0�cڂ��9����@H5נ� �P���(�A����۶}�����ֻ}��bPR�b�߶~ppr4�TP�SPI�3�}�r�10�#;A� t�
`���1���96�����%C�� Aف��J�bIncr�	����\�`��1o5qni4�MNINp	xP�`����!��Hour_  � 2�21 �A�AVM���0 ���TUP ��?J545 ���6162�VC�AM  (��CLIO ���R6�N2�MSC� "P ��STYL�C�28�~ 13\�NRE� "FHRM S�CH^�DCS}U%ORSR {b��04 �E�IOC�1 j 5742 � os| �? egist��Ի��7�1�oMASK�934"�7 ��OCO ���"3�8��2���� 0 HB��ڢ 4�"39N� R�e�� �LCHK�
%OPLG%��3�"%MHCR.%MCd  ; 4? ��6 d�PI�54�s� D[SW%MD� pQ�K!637�0�0p"�Y1�Р"4 �6<2?7 CTN K � +5 ���"7��<2�5�%/�T�%FRD�M� �Sg!��9�30 FB( NBA��P� ( HLB  7Men�SM$@jB�( PVC ��290v��2HTC�C?TMIL��\@?PAC 16U�hA�J`SAI \@ELN���<29s�UE�CK �b�@FRM� �b�OR���I�PL��Rk0CSXsC ���VVFna}Tg@HTTP �N!26 ��G�@~obIGUI"%�IPGS�r� H863 qb�!�07r�!�34 �r�84 �\so`! Qx`CC3� Fb�21�!969 rb!51 ���!S53R% 1!s3!���~�.p"9js V{ATFUJ775"���pLR6^RP�WS�MjUCTO�@xT5�8 F!80���1X�Y ta3!770 ���885�UOL�  GTSo
�{` L�CM �r| TSS��EfP6 W�\@CPgE `��0VR� �l�QNL"��@00�1 imrb�c3� =�b�0���0�`6� w�b-P- R-��b8n@5EW�b9 �Ґa� ���b�`ׁ~�b2 2000���`3��`4*5�`5 !�c�#$�`7.%�`�8 h605? U�0�@B6E"aRp76� !Pr8 t�a�@�tr2 iB/d�1vp3�vp5 ȂRtr9Σ�a4@-pN�r3 F��r5&0�re`u��r7 ��r�8�U�p9 \h7�38�a�R2D7�"�1f��2&�7<� �3 7iC���4>w5Ip�Or60� C�L�1bEN�4 I�pyL�uP��@N�&-PJ8�N�8NeN�C9 H�r`�E�b7]�|���8�ВࠂG9 2��a`0�q�Ђ5�%U097 �0��@1�0���1� (�q�3 5R ���0���mpU���0�0�7*�H@(q��\P"RB6�q124�b;��@���@�06� x�3 pB�/x�u ��x�6 H606�a1� ��7 6 ���p��b155 ����7>jUU162 ��3 g��4*�65 2e "_��P�4#U1`���B1���`=0'�174 �q���P�E186 R L��P�7 ��P�8&��3 (�90 B�/�s191����@2s02��6 3���A�RU2� d��O2 b2h`��4��b��2�4���19v RQ�2��u2d�Tpt)2� ��H�a2hP�$2�5���!U2�p�p"
�2�p��@5�0-�@��8 @�9��T�X@�� �e5�`rb	26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0@�gqGA���a�52ѐ�Ḳ6�6�0ہ5� ׁ2��84�E��9�EU5@ٰE\�q5hQ`S�2ޖ5�p\w�۲�pJ �4-P��5�p1\t�H�-4��PCH�7j��phiw�@��P�x��?559 ldu� P �D���Q�@�������A �`.��P>��8�g581�"�q58�!�AM۲T�A iC�a589��@�x���F�5 �a��12׀ 0.�1���,�2�����,�!P\h8��Lp ���,�7��6�084�0\� ANRS 0C}A��p��{��sran��FRA�� �Д�е���A%�� �ѹ�Ҍ�����(�� ��Ќ���З���������ь����$�G��1��ը��������� xS�`�q�  �����`6�4��M��iC/50T-H������*��)p46��� C��xN����m75s֐�� Sp��b46���v����ГM-7�1?�7�З����4A2������C��-��F��70�r�E��/h����O$��rlD���c7c7C� q��Ѕ���L��/���2\imm7c7�g������`���(��e�����"� �������a r��&c�T,�Ѿ�"��,��� ��x�Ex�m7�7t����k���5������)�iC��-HS-� B
_� >���+�Т�7U�]P���Mh7�s��a7������-9?�?/260L_������Q�������]�9pA/@���q�S�х��^�h621��c��92������.�)92c0�g$�@������)$��5$���pcylH"O"
�21�8��t?�350� ���p��$�
�� F�350!���0�x�9�U/0\m9��M9A3��4%�� s��3M$��X%u<���"him98J3����� i d�"m4~��103p�� ����h�794̂�&R���H �0����\���g�5A U��՜��0���*2� �00��#06�а�Ճ�է!07{r  ��������kЙ@�����EP�#�������?��#!�;&0s7\;!�B1P��@�A��/ЁCBׂ2�!��:/��?�ҽCD25�L����0�"l�2BL
#��B��\20�2_�r�re� ��X��1��N����A@��z��`C�pU��`��04��Dy	A�\�`fQ��s�U���\�5  ��� p�^t��<$85���+P=�ab1l��1LT��lA8�!uDnE(�.20T��J�1 e�bH85���b�Ռ�5[�16Bs��������d2��x��m6t!`Q����b�ˀ���b#�(�6iB ;S�p�!��3� ���b�s��-`�_�W80�_����6I	$�X5�1�U85��R�p6S����/�/+q�!@�q��`�6o��5m[o)�m6sW��Q�|�?��set06p h��3%H�5��10p$@����g/�JrH��?  ��A��856����F�� ���p/2��h�܅�✐)�5��̑v�𘜐(��m6��Y�H�ѝ̑m�6�Ҝ��ae6�DM����-S�+��H2�����Ҽ� � �r̑��✐��l���p1���F����2�\t6h T6H����Ҝ�'Vl ���ᜐ�V7ᜐ/�(���;3A7��p ~S��������4�`堜��V���!3��2��PM[��%ܖO�chn��vel5���8�Vq���_arp#���̑�.���2l_h�emq$�.�'�6415���5���?����F�����5g�L�ј�[���1��𙋹1<����M7NU�Р���eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h������ u���㜐��ZS0�!ܑ4���M-����S�$̑�ք �� 0���<�����07shJ�H�v�À�sF� �S*󜐳���̑���vl�3�A�T�#��Q�0��Te��q�pr����T@75j�5�dd�̑ 1�(UL�&�(�,���0��\�?���̑�a�� xSt���a�eD�w�2��(�	�2�C��A/���\�+p�<����21 (ܱ�CL S����B̺@��7F���?�<�lơ1L����c� ���u19�0����e/q���O���9�K��r9 (��,�Rs�ז�5�<G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O���M1!41w���2T@� _std��G�y�� �ң�H� jdgm����w0\� �1L� ��	�P�~�W*�b���t 5������3�,���E{���d���L��5\L��3�L�|#~���~!���4�#��O����h�L6A�������a2璥���44������[6\j4s ��·���#��ol�E"w�8Pk�����?0x j�H1�1Rr�>��]�2a�2Aw�P ��	2��|41�8��ˡ��@{� �%�A<��� +� ?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R�� ˑb�W���Fs���) �ѐ�!���a�1�����5��16�16C���C����0\imBQ��d����b��\Be5�-���DiL����O�_�<ѠPEtL �E�RH�ZǠPgω�am1l��u���̑�b@�<����<�$�T� ̑�F����Ȋ�DpbĜ�X"�ᒢ��pĻ ���^t��9��0\� j971\�kckrcfJ�F�s�����c��e "CTME�r�����!|�a�`main.[�8�g�`run}�_vc�#0�w�1Oܕ�_u����bctme���Ӧ�`ܑ�j73�5�- KARE�L Use {�U���J��1���p� Ȗ�9�B@���L�9��7j[�atk208 "K��(Kя��\��9��a���̹����cKRC4�a�o ��kc�qJ� &s�����Grſ�fs�D��:y��s��A1X\�j|хrdtB�, L��`.v�q�� �spǑIf�Wfj52��TKQuto Seut��J� H5K7536(�932���-91�58(�9�BA��1(�74O,A$�(TCP Ak���/�)Y� �\tpqtool.v���v���! con�re;a#�Cont�rol Re�b{le��CNRE(� T�<�4�2���D�)���NS�552��q(g�� (򭂯4X�cOux~�\sfuts�UTS`�i�栜���At�棂��? 6�T�!�SA OO+D6���������,!��6c+� igt�t6i��I0�T�W8 ���la��vo58�o�bFå򬡯i��Xh��!Xk�0Y!8�\m6e�!6EC���v��6���������<16�A���A�6s����U�g�T|�,����r1�qR����Z4�T�����,#�eZp)g����<ONO0���uJ��tCR;��F<�a� xSt�f���prdsuchk� �1��2&&?���t��*D%$�r(�✑ �娟:r��'�s�qO��<scrc�C�\At�trldJ"o��\�V����Pay�lo�nfirm�l�!�87��7��A�3ad�! �?@ވI�?plQ��3���3"�q��x pl��`���d7��l�calC�uDu���;���mov�����initX�:s8O��a8�r4 ��r67A4|��e Genera#tiڲ���7g2q$g R� (S�h��c ,|�bE��$Ԓ\�:�"���4��4�4�. sg��5�F$d6"�e�!p "SHA�P�TQ ngcr pGC�a(�&"� ���"GDA¶��r�6�"aW�/�$d�ataX:s�"tp�ad��[q�%tput;a__O7;a�o8�1�yl+s�r�?�:�#$�?�5x�?�:c O�:Ay O�:�IO�s`O%g�qǒ�?�@0\ۜ�"o�j92;!�Pp�l.Collis�QSkip#��@5� �@J��D��@\ވ�C(@X�7��7�|s}2��ptcls�#LS�DU�k?�\_� ets�`�< �\�Q��@���`dcKLqQ�FC;��J,όn��` (��4eN����T�{���' j(�c�q���/IӸaȁ<��̠H������зa�e\mcc�lmt "CLM��/��� mate\v��lmpALM�?>p7qmc?�����2vm�q��%�3s��_�sv90�_x_msu�2L^v_� K�o��{in�8(3r<�c_logr��r�trcW� �v_3�~yc��d�<�ste��der$c;Ce� Fiρ��R��Q�?�l�enter߄|��(�Sd��1�TX�+fZK�r�a99sQ9+��5�r\tq\� _"FNDR����STDn$�LANG�Pgui��D⠓�S������csp�!ğ֙uf䟀ҝ�s����$�����e +�=����������������w�H�r\fn�_�ϣ��$`x�tcp�ma��- TCP������R638 aR�Ҡ��38��M7p,���Ӡ�$Ӡ��8p0Р�VS,�>�tk��99�a��B3���P�զԠ��D�2�����UI��t���hqB���8���������p���re8�ȿ��exe@4π��B���e38�ԡG�r�mpWXφ�var @�φ�3N�����v�x�!ҡ��q�R�BT $cOP�TN ask E�0��1�R MAS�0�H593/�96g H50�i�480ԅ5�H0��m�Q�K(��7�0�g�Pl�h�0ԧ�2�ORDP���@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`am��b��7�.f���u�d��r��splayD�E���1wПUPDT Ub��8o87 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60�q��B����qs�can��B���aAd@�������q`� �䗣�#��К�`2�� vlv��Ù�$�0>�b���! S���Easy/К�Ut�il��룙�511# J�����R7 ���Nor֠��inc�),<6Q�� �`c��"4�[���986(FVRx So����q�nd6����P��4� a\ (��
  ������"�d��K�bdZ����men7���- Me`tyFњ�Fb��0�TUa�577?i3R��\�5�au?��!� n����f������l\m�h�Ц�űE|h#mn�	��<\O�$��e�1�� l!���y��Ù�\|p�����B���Ћmh �@��:.aG!�� �/�t�55�6�!X��l�.us��Y/k)eOnsubL���eK�h�� �B\1;5g?�y?�?�?D��?*rmx�p�?Ktbox O�2K|?�G��C?A%das���?1ӛ#� � TR��/��P�4B�`�U@�P�V�P"�Q�P0�U �PO��P�"�T3�U�P �f�Pk"�2}�4�T�P �f�P2�"�Q5�S�Q@���R?Ă�Q3t.�PF׀al��P+O�n�P517��IN0a���Q(}g��PES	Tf3ua�PB�l�i�g�h�6�aq��P �� xS��` � n�0mbump�P�Q969g�69�Qq��P0�baAp�@>Q� BOX��,�>vche�s�>ve�tu㒣=wffse�3���]�;u`aW��:zol�sm<u�b�a-��]D�K�ib�Q�c����Q<twaǂ �tp�Q҄Taror Recov�br�O�P�642�����a�q��a⁠QErǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>��pjot��PXc��C��1�adb -�ail���nag���b�QR629�a�Q��b�P�  �
 � �P��$$CL~[q ����������$�PS?_DIGIT���"�!�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��������*璬1:P�RODUCT�Q0�\PGSTK�bV�,n�99�\����$FEAT_INDEX���~�� �搠ILECOM�P ;��)���"��SETUPo2 <��?�  N !��_AP2BCK �1=�  �)}6/E+%,/i/��W/�/~+/�/O/ �/s/�/?�/>?�/b? t??�?'?�?�?]?�? �?O(O�?LO�?pO�? }O�O5O�OYO�O _�O $_�OH_Z_�O~__�_ �_C_�_g_�_�_	o2o �_Vo�_zo�oo�o?o �o�ouo
�o.@�o d�o���M� q���<��`�r� ���%���̏[���� ���!�J�ُn����� ��3�ȟW������"� ��F�X��|����/� ��֯e������0��� T��x������=�ҿ �s�ϗ�,ϻ�9�b�t� P/ 2) *.VRiϳ�!�*���������Ɲ�PC�7�!�F'R6:"�c��χ��T��߽�Lը����x���*.F���>� �	N�,�k�x�ߏ��STM �⠸���Qа���!��iPendant? Panel���H��F���4������GIF�������pu����JPG&�P��<����	�PANEL1.D	T��������2�Y�G��
3w�����//�
4�a/��O///�/�
TP�EINS.XML�/���\�/�/�!�Custom T?oolbar?��PASSWOR�D/�FRS:�\R?? %Pa�ssword Config�?��? k?�?OH�6O�?ZOlO �?�OO�O�OUO�OyO _�O�OD_�Oh_�Oa_ �_-_�_Q_�_�_�_o �_@oRo�_voo�o)o ;o�o_o�o�o�o*�o N�or��7� �m��&���\� ����y���E�ڏi� �����4�ÏX�j��� �����A�S��w�� ���B�џf������� +���O��������� >�ͯ߯t����'��� ο]�򿁿�(Ϸ�L� ۿpς�Ϧ�5���Y� k� ߏ�$߳��Z��� ~�ߢߴ�C���g��� ��2���V����ߌ� ��?����u�
��� .�@���d������)� ��M���q�����< ��5r�%�� [�&�J� n��3�W� ��"/�F/X/�|/ /�/�/A/�/e/�/�/ �/0?�/T?�/M?�?? �?=?�?�?s?O�?,O >O�?bO�?�OO'O�O KO�OoO�O_�O:_�O ^_p_�O�_#_�_�_Y_��_}_o�_�_Ho)f��$FILE_DG�BCK 1=���5`��� ( �)
S�UMMARY.DyGRo�\MD:�o��o
`Diag� Summary��o�Z
CONSLOG�o�o�a
J�a�ConsoleO logK�[�`�MEMCHECK�@'�o�^qMe�mory Dat�a��W�)>�qHADOW����P��sShad�ow Chang�esS�-c-��)	FTP=��9�����w`qmmen�t TBD׏�W0�<�)ETHERNET̏�^�q��Z��aEther�net bpfiguration[���P��DCSVRF�ˏ��Ïܟ�q%��� verify� allߟ-c1P{Y���DIFFԟp��̟a��p%��diffc���q���1X�?�Q�� �����X��CH�GD��¯ԯi��px��� ���2`�G�Y��� ��� �GAD��ʿܿq��p���Ϥ�FY3h�O�aώ�� ��(�GAD������y��p�����0�UPDAT�ES.�Ц��[FORS:\�����a�Updates �List���kPS�RBWLD.CM�.��\��B��_pP�S_ROBOWEL���_����o��,o !�3���W���{�
�t� ��@���d�����/ ��Se����� N�r� =� a�r�&�J� ��/�9/K/�o/ ��/"/�/�/X/�/|/ �/#?�/G?�/k?}?? �?0?�?�?f?�?�?O �?OUO�?yOO�O�O >O�ObO�O	_�O-_�O Q_c_�O�__�_:_�_ �_p_o�_o;o�__o �_�o�o$o�oHo�o�o ~o�o7�o0m�o � ��V�z� !��E��i�{�
��� .�ÏR���������� .�S��w������<� џ`������+���O� ޟH������8���߯�n����$FIL�E_��PR����������� �MDONL�Y 1=4�� 
 ���w�į�� 诨�ѿ�������+� ��O�޿sυ�ϩ�8� ����n�ߒ�'߶�4� ]��ρ�ߥ߷�F��� j�����5���Y�k� �ߏ���B�����x� ���1�C���g���� ��,���P����������?��Lu�VI�SBCKR�<�a��*.VD|�4 OFR:\��4 �Vision VD file�  :LbpZ�# ��Y�}/$/� H/�l/�/�/1/�/ �/�/�/�/ ?�/1?V? �/z?	?�?�???�?c? �?�?�?.O�?ROdOO �OO�O;O�O�OqO_ �O*_<_�O`_�O�__�%_�_�MR_GR�P 1>4�L~�UC4  B�P�	 ]�ol`��*u����RHB ��2 ���� ��� ���He�Y�Q`ork bIh�oJd�o�Sc�o��oE�� LQ�hJ��F�;5U�aR���V�o�!}B���A��b �Q6���;�o{0  =�s�lqhr�G�xq~�o� F@ �r��d�aX}J��NJ�k�H9�H�u��F!��IP�sX}?�`�.�9�<9��896C'�6<,6\b� X1�,.�g�R���v�A�PA�����|�ݏ x���%��I�4�F� �j�����ǟ���֟���!��E�`r�UBH�P�c������ů��R
6�P;�kP;�˯R��e�Q �cB��P5���@�33@���4�m�,�/@UUU��U�~w��>u.�?! x�^��ֿ���3���=[z�=�̽�=V6<�=��=�=$q���~��@8�i�7G��8�D��8@9!�7�ϥ�@Ϣ���cD��@ D�� CϬ����C��P��P' �6��_V� m�o��To ��xo�ߜo������ A�,�e�P�b���� ����������=�(� a�L���p��������� ��������*��N9 r]������ ��8#\nY �}������� /ԭ//A/�e/P/�/ p/�/�/�/�/�/?�/ +??;?a?L?�?p?�? �?�?�?�?�?�?'OO KO6OoO�OHߢOl��� �ߢ��O�� _��G_bO k_V_�_z_�_�_�_�_ �_o�_1ooUo@oyo dovo�o�o�o�o�o�o Nu� �������� ;�&�_�J���n����� ��ݏȏ��%�7�I� [�"/�描�����ٟ �������3��W�B� {�f�������կ���� ���A�,�e�P�b� �������O�O�O� �O�OL�_p�:_���� �Ϧ��������'�� 7�]�H߁�lߥߐ��� ��������#��G�2� k�2��Vw������ �����1��U�@�R� ��v������������� -Q�u�� �r��6��) M4q\n�� ����/�#/I/ 4/m/X/�/|/�/�/�/ �/�/?ֿ�B?�f? 0�BϜ?f��?���/�? �?�?/OOSO>OwObO �O�O�O�O�O�O�O_ _=_(_a_L_^_�_�_ �_���_��o�_o9o $o]oHo�olo�o�o�o �o�o�o�o#G2 kV{�h��� ����C�.�g�y� `����������Џ� ��?�*�c�N���r� �������̟��)� �M�_�&?H?���?�� �?�?�?����?@�I� 4�m�X�j�����ǿ�� �ֿ����E�0�i� Tύ�xϱϜ������� ��_,��_S���w�b� �߭ߘ��߼������ �=�(�:�s�^��� ��������'�9�  �]�o����~����� ��������5 Y DV�z���� ��1U@y d��v�����/ Я*/��
/�u/��/ �/�/�/�/�/�/?? ;?&?_?J?�?n?�?�? �?�?�?O�?%OOIO 4O"�|OBO�O>O�O�O �O�O�O!__E_0_i_ T_�_x_�_�_�_�_�_ o�_/o��?oeowo�o P��oo�o�o�o�o +=$aL�p� ������'�� K�6�o�Z������ɏ ��폴� ��D�/  /z�D/��h/ş��� ԟ���1��U�@�R� ��v�����ӯ����� �-��Q�<�u�`��� `O�O�O���޿�� ;�&�_�J�oϕπϹ� ���������%��"� [�F��Fo�ߵ����� �o��d�!���W�>� {�b���������� ����A�,�>�w�b� ���������������=��$FNO ���\��
F�0l q  FLA�G>�(RRM_�CHKTYP  �] ��d ��] ��OM� _MsIN� 	���� ��  XT SS�B_CFG ?�\ �����OT�P_DEF_OW�  	��,I�RCOM� >�$�GENOVRD_�DO��<�lT[HR� d�dqo_ENB] q�RAVC_GRP� 1@�I X (/ %/7//[/B/ /�/x/�/�/�/�/�/ ?�/3??C?i?P?�? t?�?�?�?�?�?OO OAO(OeOLO^O�Oo�ROU�F\� ��,�B,�8�?���O�O�O�	__���  D�E_�Hy_�\@@m_B��=�vR/��I�O�S+MT�G�SUo�o&oRHOSTC��1H�I� �\�zMSM�l[�bo�	12�7.0�`1�o  e�o�o�o#z �oFXj|�l60s�	anonymous��������4ao�&�&� �o�x��o������ҏ �3��,�>�a�O� ���������Ο�U%� 7�I��]����f�x� �������ү���� +�i�{�P�b�t����� �������S�(� :�L�^ϭ�oϔϦϸ� �����=��$�6�H� Zߩ���Ϳs������ ����� �2���V�h� z��߰��������� 
��k�}ߏߡߣ�� �߬���������C� *<Nq�_��� ���-�?�Q�c�e J��n���� ���/"/E�X/ j/|/�/�/�% '/?[0?B?T?f?x? ��?�?�?�?�??E/�W/,O>OPObO�KDaE�NT 1I�K sP!�?�O  �P�O�O�O�O�O#_�O G_
_S_._|_�_d_�_ �_�_�_o�_1o�_o go*o�oNo�oro�o�o �o	�o-�oQu 8n������ ��#��L�q�4��� X���|�ݏ���ď֏�7���[���B�QUICC0��h�z�۟��1ܟ��ʟ+����2,���{�!ROUTER|�X�j��˯!PCJOG�̯��!192�.168.0.1�0��}GNAME �!�J!ROB�OT�vNS_CF�G 1H�I ��Auto�-started^�$FTP�/�� �/�?޿#?��&�8� JϏ?nπϒϤ�ǿ�� [������"�4ߵ&�� ��������濜����� �����'�9�K�]�o� ������������� �/�/�/G���k��ߏ� ������������ 1T���Py��� ��"�4�	H-|� Qcu�VD�� ��/�;/M/_/ q/�/����/
/�/ >?%?7?I?[?*/? �?�?�?�/�?l?�?O !O3OEO�/�/�/�/�? �O ?�O�O�O__�? A_S_e_w_�O4_._�_ �_�_�_oVOhOzO�O �_so�O�o�o�o�o�o �_'9Kno�o �����o*o<o NoP5��oY�k�}��� ��pŏ׏����0����C�U�g�y���_�T_ERR J;������PDUSIZW  ��^P�����>ٕWRD ?�z���  guest����+�=�O�a�s�*�S�CDMNGRP �2Kz�ÐC��۠\��K��� 	P01.1�4 8�q   �y��B  �  ;�����{ �����������������������~ �ǟI�4�m�X��|��  i  �  
����� ����+��������
��k�l�.x�����"�l�ڲ۰s�d��������_GR�OU��L�� ���	��۠07K�Q?UPD  ���YPČ�TYg������TTP_AU�TH 1M�� �<!iPend�an���<�_��!KAREL:q*�����KC%��5�G��VISI?ON SETZ���|��Ҽߪ���� �����
�W�.�@���d�v���CTRL CN�������
��FFF9E3����FRS:D�EFAULT��FANUC W�eb Server�
������q��������������WR�_CONFIG ;O�� ����IDL_CPU_kPC"��B���= �BH#MIN�.�BGNR_I�O��� ���% NP�T_SIM_DO�s}TPMOD�NTOLs �_�PRTY�=!O�LNK 1P�� �'9K]o>�MASTEr ��|���O_CFG�ƟUO����CY�CLE���_A�SG 1Q���
 q2/D/V/h/z/ �/�/�/�/�/�/�/
?�?y"NUM�x��Q�IPCH���£RTRY_C�N"�u���SCRQN������ ���R����?���$J23_DS/P_EN����~�0OBPROC�3ܷ�JOGV�1S�_�@��8�?р';ZO'??0CPO�SREO�KANJI_�Ϡu�A#��3T ���E�O�ECL_LM B2e?�@�EYLOGGINʭ������LA�NGUAGE ,_�=� }Q���LG�2U�����J �x�����PC �� �'0������MC:\RS�CH\00\˝L�N_DISP �V�������TOYC�4Dz\A�S�OGBOOK W+��o���o�o���Xi�o�o�o�o�o�~}	x(y��	�ne�i�ekElG_BUFF 1X�	��}2����Ӣ ������'�T� K�]�����������ɏ ۏ���#�P��Ëq�DCS Zxm =���%|d1h`�ฟʟܟ�g�IO ;1[+ �?'����'�7�I�[�o�� ������ǯٯ���� !�3�G�W�i�{�����б�ÿ׿�El TM  ��d��#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g��yߋߝ߈t�SEVt�0m�TYP΁� ��$�}�AR�S"�(_�s�2FL 31\��0�������������5�T�P<P���DmNGNAM�4�U�f�7UPS`GI�5�A��5s�_LOAD�@G %j%;DF��GI6����MAXUALRM B7�P8��y���3�0Q]&q��Ca]s�@3�~�� 8@=@^+� طv	���V0+�P�A5d�1r���U�� ����E(i Ty������ �/ /A/,/Q/w/b/ �/~/�/�/�/�/�/? ?)?O?:?s?V?�?�? �?�?�?�?�?O'OO KO.OoOZOlO�O�O�O �O�O�O�O#__G_2_ D_}_`_�_�_�_�_�_ �_�_o
ooUo8oyo do�o�o�o�o�o�o�o��o-��D_LDX�DISA^�� �M�EMO_APX�E� ?��
  �0y�����������ISC 1_�� �O�� ��W�i�����Ə�� ���}��ߏD�/�h� z�a����������� ���@���O�a�5� �����������u�� ׯ<�'�`�r�Y���� ��y�޿�ۿ���8� ��G�Y�-ϒ�}϶ϝ� ����m�����4��X��j�#�_MSTR �`��}�SCD 1as}�R���N��� �����8�#�5�n�Y� ��}���������� ��4��X�C�|�g��� ������������	 B-Rxc��� ����>) bM�q���� �/�(//L/7/p/ [/m/�/�/�/�/�/�/ ?�/"?H?3?l?W?�?�{?�?�?�?n�MKC_FG b���?~��LTARM_�2�cRuB ��3WpTNBpMETsPUOp�2�����NDSP_CMN�TnE@F�E�� 	d���N�2A�O�D��EPOSCF�G��NPSTOL 1�e-�4@�<#�
;Q�1;UK_YW7_Y_ [_m_�_�_�_�_�_�_ o�_oQo3oEo�oio�{o�o�a�ASING_CHK  �M^AqODAQ2CfO��7J�eDEV }	Rz	MC:'|�HSIZEn@�����eTASK %�<z%$123456789 ��u�gTRIG 1g�� l<u%���3`���>svvYPaq���kEM_INF� 1h9G �`)AT&�FV0E0(���)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏP� �t�������]�ί�� ���(�۟�^�� #�5�����k�ܿ� � ��ů6��Z�A�~ϐ� C���g�y�������� 2�i�C�h�ό�G߰� �ߩ��ߙϫ������ ��d�v�)ߚ��߾�y� ��������<�N�� r�%�7�I�[������ 9�&��J[��g��>ONITO�R�@G ?;{  � 	EXEC�1�3�2�3�4��5��p�7�8
�9�3�n�R� R�RRR R(R4R@RL�R2Y2e2q2�}2�2�2�2��2�2�3Y3�e3��aR_GRP_SV 1it�z�q(�5�
��5o��۵MO~q�_DCd~�1PL_NAME !<u�� �!Def�ault Per�sonality� (from FwD) �4RR2k!� 1j)TEX)�TH��!�AX d �?>?P?b?t?�?�?�? �?�?�?�?OO(O:O�LO^OpO�O�O�Ox2 -?�O�O�O__0_B_T_f_x_�b<�O�_�_ �_�_�_�_o o2oDo�Voho&xRj" 1o��)&0\�b, ��9��b�a @D7�  �a?��c�a�?�`�a�aA'�6x�ew;�	l�b�	 �x7Jp��`�`�	p �< ��(p� �.r� K��K ��K�=*�J���J?���JV��kq`q�P�x�|� �@j�@T;f�r�f�q�acrs��I�� ��p����p�r�ph}�3���´  ���>��ph�`z���꜖"�Jm�q� H�N��ac���$�dw��  _�  P� Q� }�� |  а��m�Əi}	'� �� �I� ��  ����:��È�È=̣��(��#�a	����I  �n �@H�i~�ab�Ӌ�b��$w���"N0�� � 'Ж�q�p@2?��@����r�q�5�C�pC0C�G@ C����`O
�A1]w@B�UV~X�
nwB0"h�A��p�ӊ�p@����aDz���֏����Я	�pv�( �� -���I��-�=��A�a��we_q�`�p �?�ff ��m��>� ����ƼЇ!@ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`�� <
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC��������#/*/c/N/�wi�����v/C�`� CHs/`
=$�p��<!�!��ܼ�'��3A�A�AR�1AO�^?�$��?���±�
=ç>�����3�W
=�#��]�;e��?������{�����<�>(��B�u��=�B0�������	R��zH�F��G���G���H�U`E����C�+��}I#��I��HD��F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*OO NO9OrO]O�O�O�O�O �O�O�O_�O8_#_\_ G_�_�_}_�_�_�_�_ �_�_"oooXoCo|o go�o�o�o�o�o�o�o 	B-fQ�u �������,� �P�b�M���q����� Ώ���ݏ�(��L� 7�p�[������ʟ�� �ٟ���6�!�Z�E��W���#1( ���9�K���ĥ ������Ư!3�8����!4Mgs8��,�IB+8�J���a���{� d�d�����ȿ���ڼJ%P8�P�=:�GϚ�S�6�h�z���R�Ϯ����������  %�� ��h�V� ��z߰�&�g�/9�$�������7����pA�S�e�w�  ������������2� F�$�&Gb	��������!C���@���8���~��F� DzN���� F�P DC�������)#B��'9K]o#?̯��@@v
4$R8�8��8�.
 v��� !3EWi{��p��:� ������1��$MS�KCFMAP  ���� ����(.�ON�REL  ��!9��EXCFENBE'
#7%^!�FNCe/W$JOG_OVLIME'dO �S"d�KEYE'��%�RUN�,��%�SFSPD�TY0g&P%9#SI�GNE/W$T1MO�T�/T!�_CE_GRP 1p��#\x��?p��? �?�?�?�?O�?O BO�?fOO[O�OSO�O �O�O�O�O_,_�OP_ _I_�_=_�_�_�_�_��_oo�_:o�T�COM_CFG 1q	-�vo�o�o}
Va_ARC_b"��p)UAP_C�PL�ot$NOCH�ECK ?	+ �x�%7 I[m���������!�.+NO_WAIT_L 7l%S2NT^ar	+z�s�_ERR_1s2s	)9�� ,o̏ޏ��x���&�^�dT_MO��t��, J*oq�9�_PARAM��u	+��a�ß'g{��� =?�345678901��,� �K�]�9�i�������0ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDSP��c#6p(OFFSE?T_CART�o���DISƿ��PEN_FILE尨!�a�i��`OPTION�_IO�/��PWO_RK ve7s# ��V�ؤ!!�8p�4�p�	 ���p���<���RG_D?SBL  ��P#���ϸ�RIEN�TTOD ?�C�� !l�UT_S/IM_D$�"����V��LCT �w}�h�iĜa[�1�_�PEXE�j�RAATvШ&p%� ��2^3�j)TEX)TH}�)�X d3� ������%�7�I�[� m�����������@���!�3�E���2�� u���������������c�<d�ASe w���������Ǎ�^0OUa0o�(��(�����u2, ����O H @D� M [?�aG?��cc�D][�Z��;�	ls��xJ���������<w ��� ���2�H(��H3k�7HSM5G�2�2G���Gp
1͜�'f�/-,�2�CR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t�!�/ �/�"t�32����/6  ���P%�Q%��
%�|T��S62�q?'e	'� � �2�I� �  ���+==���г?�;	�h	�0�I�  �n @@�2�.��Ov;��ٟ�?&gN�]O  '�'�uD@!� C�C�A@F#H!�/�O�O sb�
���@�@"��@�e`0B�QqA�0Yv: �13Uwz$oV_�/z_e_��_�_	��( ?�� -�2�1 �1ta�Ua�c���:A�r���.  �?��ff���[o"o�_U�`oXÜQ8���o�j�>�1  Po�V( ���eF0�f�Y���^L�?����xb��P<
6b<���;܍�<����<� <�&�,/aA�;r�@|Ov0P?fff?�0�?&ip�T@�.�{r�J<?�` �u#	�Bdqt�Yc� a�Mw�Bo��7� "�[�F��j������� ُ����3�����,���(�E�� �E��3G+� F��a��ҟ�����@,��P�;���B�pAZ�>��B��6�<Oί D���P��t�=���a��s�����6j�h��<7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�%?��?���������#	Ę��P �N|F|CH���Ŀ�������@I�_�'��3A�A�AR�1AO�^?��$�?��� ����
=ç>�����3�W
=�s#� U��e���B���@��{�����<���(��B�u���=B0�������	�b�H�F��G���G���H�U`E����C�+��I�#�I��H�D�F��E���RC�j=[�
�I��@H��!H�( E<YD0߻��� ������� �9�$�]� H�Z���~��������� ����#5 YD} h������� 
C.gR�� �����	/�-/ /*/c/N/�/r/�/�/ �/�/�/?�/)??M? 8?q?\?�?�?�?�?�? �?�?O�?7O"O[OmO XO�O|O�O�O�O�O�O��O�O3_Q(���ٙ��b��gUU���W_i_2�3��8��_�_2�4Mgqs�_�_�RIB+�_��_�a���{�miGo5okoYo�o�}l��P'rP�nܡ ݯ�o=_�o�_�[R?Q�u���  �p���o� �/��S��z
uүܠ�������ڱ����એ�����   /�M�w�e��������l�2 F�$��Gb��t��a�`�p�S�C�y�@p�5�G��Y�۠F� Dz��� F�P �D��]����پ���ʯܯ� ��~�?_���@@�?��K�K���K���
 �|����� ��Ŀֿ�����0��B�T�fϽ�V� ����{��1��$P�ARAM_MEN�U ?3���  �DEFPULSE�r�	WAITT�MOUT��RC�V�� SHE�LL_WRK.$�CUR_STYLv��	�OPT�N�PTB4�.�C�R_DECSN�� �e��ߑߣ������� ����!�3�\�W�i��{���USE_P�ROG %��%������CCR����e����_HOST7 !��!��:����T�`�V��/��X����_TIME���^��  ��GDEBUG\�˴��GINP_FLMSK����Tfp����WPGA  �����)CH����TYPE������� ���� -? hcu����� ��//@/;/M/_/ �/�/�/�/�/�/�/�/�??%?7?`?��WO�RD ?	=	�RSfu	PNeSUԜ2JOK��DRTEy�]TR�ACECTL 1�x3��� ��`�`&�?�3�6D/T Qy3�%@�0�D � �c2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�Z�.O|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��p����� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o� $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ������������(��$�PGTRACEL�EN  )�  ��(���>�_UP z/���m�u�Y��n�>�_CFG7 {m�W�(�En���PЬ� ���DEFSPD e|��'�P��>��IN��TRL �}��(�8��IPE_CONFI��}~m��m����Ԛ�>�LID����=�GRP� 1��W���)�A ���&f�f(�A+33D��� D]� C�O� A@1��Ѭ(��d�Ԭ��0�0�� 	 1��1���G ´�����B� 9����O�9�s�(��>�T?�
5�������� =��=#�
���� P;t_��������  Dz (�
H�X ~i������ /�/D///h/S/�/���
V7.10�beta1��  A�E�"�ӻ�A (�� ?�!G��!>��r�"����!���!oBQ��!A\� P�!���!2p����Ț/8?J?\?n?};� ���/��/�?}/ �?�?OO:O%O7OpO [O�OO�O�O�O�O�O _�O6_!_Z_E_~_i_ �_�_�_�_�_�_'o 2o�_VoAoSo�owo�o �o�o�o�o�o.�R=v1�/�#F@ �y�}��{m��y =��1�'�O�a��? �?�?������ߏʏ� �'��K�6�H���l� ����ɟ���؟�#� �G�2�k�V���z��� �����o��ίC� .�g�R�d��������� �п	���-�?�*�c� ����Ϯ���� ��B�;�f�x����� ��DϹ��߶������ ��7�"�[�F�X��|� �����������!�3� �W�B�{�f������� �� �����/S >wbt���� ��=Ozό� �ψ����ϼ� / .�'/R�d�v߈߁/0 �/�/�/�/�/�/�/#? ?G?2?k?V?h?�?�? �?�?�?�?O�?1OCO .OgORO�OvO�O�O�� �O�O�O__?_*_c_ N_�_r_�_�_�_�_�_ o�_)oTfx�to ���/�o/ >/P/b/t/mo�| �������3� �W�B�{�f�x����� Տ�������A�S� >�w�b����O��џ�� ����+��O�:�s� ^�������ͯ���ܯ �@oRodo�o`��o�o �o��ƿ�o���*< N�Y��}�hϡό� �ϰ��������
�C� .�g�Rߋ�v߈��߬� ����	���-��Q�c� N�ﲟ���l����� ���;�&�_�J��� n�����������,� >�P�:L������� �����(�:�3 ��0iT�x�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?a?s? ��?�?X?�?�?�?�? O'OOKO6OoOZO�O ~O�O�O�O�O*\ &_8_r���_�_���$PLID_K�NOW_M  ~�� Q��TSV ��]�P��? o"o4o�OXoCoUo�o� R�SM_GRP� 1��Z'0{`J�@�`uf�e�`
�5� �gpk 'Pe]o�� ��������S+MR�c��mT�EyQ}? yR�������� ��폯���ӏ�G�!� �-������������ ����ϟ�C���)� ����������寧����QST�a1 1�j�)���P0� A 4��E2�D�V� h�������߿¿Կ� ��9��.�o�R�d�v�@���ϬϾ����2�90� Q�<3��A3�/�A�S��4l�~ߐߢ��5���������6
��.�@��A7Y�k�}���8���������MAD � )��P�ARNUM  �!�}o+��SCH
E� S�
��f���S��UPDf�x�|�_CMP_�`�H�� �'�UE�R_CHK-�a��ZE*<RSr��_�Q_MOG����_�X�_RES_G��!���D� >1bU�y�� ���/�	/����+/�k�H/g/ l/��Ї/�/�/�	� �/�/�/�X�?$?)? ���D?c?h?����?x�?�?�V 1��U��ax�@c]�@t�@(@c\�@��@D@c[�*@���THR_INR�r�J�b�Ud2FMA�SS?O ZSGMN�>OqCMON_QU?EUE ��U�V� P~P X�N$ U�hN�FV�@END8�A��IEXE�O�E���BE�@�O�COP�TIO�G��@PR�OGRAM %��J%�@�?���BT�ASK_IG�6^O?CFG ��Oz���_�PDATA�c�.�[@Ц2=�Do Vohozo�j2o�o�o�o �o�o);M j�INFO[��m� �D������ ��1�C�U�g�y��� ������ӏ���	�dwpt�l )�QE ?DIT ��_i�>�^WERFLX	C��RGADJ M�tZA�����?נ�ʕFA��IORIT�Y�GW���MPD�SPNQ����U�G�D��OTOE@1��X� (!A�F:@E� c�Ч!�tcpn���!�ud����!i�cm���?<�XY_��Q�X���Q)�� *�1�5��P��]�@�L���p��� �����ʿ��+�=Ϡ$�a�Hυϗ�*��P�ORT)QH��P��E��_CART�REPPX��SK�STA�H�
SSA�V�@�tZ	25?00H863���_�x�
�'��X�@�swPtS�ߕߧ���/URGE�@B��x	WF��DO�F"[�W\�������WRU�P_DELAY ��X���R_HO�TqX	B%�c���R_NORMALq^xR��v�SEMI�������9�QSKIP�'��tUr�x 	7�1�1��X�j�|� ?�tU������������ ��$J\n4 ������� �4FX|j� ������/0/ B//R/x/f/�/�/�/�tU�$RCVTM�$��D�� DCR�'���Ў!=��Bv�4C �V�>�.>��z�6:e�:����������6��:�o?�� �<
6b<���;܍�>u.��?!<�&�?h?�?�?�@>��? O O2ODOVOhOzO�O �O�O�O�O�?�O�O_ _@_+_=_v_Y_�_�_ �?�_�_�_oo*o<o No`oro�o�o�o�_�o �o�o�o�o8J- n��_����� ��"�4�F�X�j�U ������ď���ӏ� ��B�T��x����� ����ҟ�����,� >�)�b�M��������� ���ïկ�Y�:�L� ^�p���������ʿܿ � ����6�!�Z�E� ~ϐ�{ϴϗ�����-� � �2�D�V�h�zߌ� �߰���������
��� .��R�=�v��k�� ���������*�<� N�`�r���������� ������&J\ ?������� �"4FXj|���!GN_ATC� 1�	; �AT&FV0E�0�ATDP�/6/9/2/9��ATA�,�AT%G1%�B960�+�++�,�H/,��!IO_TYPE'  �%�#t��REFPOS1 �1�V+ x�u/�n�/j�/
= �/�/�/Q?<?u??�?�4?�?X?�?�?�+2 1�V+�/�?�?\O��?�O�?�!3 1� O*O<OvO�O�O_�OS4 1��O�O�O�_�_t_�_+_S5 1�B_T_f_�_o	o|Bo�_S6 1��_��_�_5o�o�o�oUoS7 1�lo~o�o�o�H3l�oS8 1�%_����SMASK 1�V/  
?�M��'XNOS/�r�������!MOTE  �n��$��_CFG �����q���"PL_RANG������POWER �����SM_D�RYPRG %�o�%�P��TAR�T ��^�UME_PRO-�?�����$_EXEC_E�NB  ���GSPD��Րݘ��gTDB��
�RM�.
�MT_'�T�����OBOT_N�AME o�����OB_ORD_NUM ?��b!H863  �կ�����PC_TI�MEOUT�� xޚS232Ă1��� LTE�ACH PENDcAN��w��-���Maint�enance CGons���s�"��~�KCL/Cm�Ț

���t�ҿ No Use-p��Ϝ�0�NPO�\򁋁��.�oCH_L�������q	��s�MAVGAIL�����糅���SPACE1 ;2��, j�߂ �D��s�߂� �{~S�8�?�k� v�k�Z߬��ߤ��ߚ � �2�D���hߊ�|� ��`��������� � �2�D��h��|� ��`���������y���2����0�B��� f�����{���3);M_ ������/� /44FXj |*/���/�/�/?(??=?5Q/c/u/ �/�/G?�/�/�?O�? $OEO,OZO6n?�? �?�?�?dO�?�?_,_@�OA_b_I_w_7�O �O�O�O�O�_�O_(o�Ioo^oofo�o8 �_�_�_�_�_�oo6o Ef){����G �o� t���
M� � ��*�<�N�`�r����� ��w���o�収���d.��%�S�e�w� ����������Ǐَ�� �Θ8�+�=�k�}��� ����ůׯ͟���� %�'�X�K�]������� ��ӿ������#��E�W� `� @�������x�����\�e���������� �R�d߂�8�j߬߾� �ߒߤ���������� 0�r���X�����������8����
��ύ�_MODE�  �{��S E��{|�2�0�����3�	S|)�CWORK_AD޳�0��+R  �{�`� �� _INTVAL����d���R_OPT�ION� ���H VAT_GRPw 2��upG(N�k |��_���� �/0/B/��h�u/T�  }/�/�/�/�/�/�/ ?!?�/E?W?i?{?�? �?5?�?�?�?�?�?O /OAOOeOwO�O�O�O �OUO�O�O__�O=_ O_a_s_5_�_�_�_�_ �_�_�_o'o9o�_Io oo�o�oUo�o�o�o�o �o�o5GYk- ���u���� �1�C��g�y���M� ����ӏ叧�	��-� ?�Q�c����������� ����ǟ�;�M��_����$SCAN�_TIM��_%�}�R �(�#�((�<04Wd d 
�!D�ʣ��u��/�����U�"�25���@�d5�P�g��]	����������dd�x�  P~���� ��  8� ҿ�!���D��$�M�_�q� �ϕϧϹ��������8ƿv��F��X��/� ;�o�b��pm��t�_DiQ̡  � l�|�̡ ĥ�������!�3�E� W�i�{�������� ������/�A�S�e� ]�Ӈ����������� ��);M_q ������� r���j�Tfx� ������// ,/>/P/b/t/�/�/�/p�/�/�%�/  0�� 6��!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O *�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo �O�OJ�o�o�o�o�o �o�o 2DVh z�������
�7?  ;�>�P� b�t���������Ǐُ ����!�3�E�W�i��{�������ß � ş3�ܟ��&�8�J��\�n�������������ɯ����,�� �+�	12�345678��W 	� =5���@f�x���������� ���
��.�@�R�d� vψϚ�៾������� ��*�<�N�`�r߄� �Ϩߺ��������� &�8�J�\�n�ߒ�� �����������"�4� F�u�j�|��������� ������0_�T fx������ �I>Pbt �������! /(/:/L/^/p/�/�/ �/�/�/�/�2�/�?�#/9?K?]?�i�Cz  Bp˚ /  ��h2��*��$SCR_GR�P 1�(�U8�(�\x�d�@ � ��'�	 ?�3�1 �2�4(1*�&�I3�Fp1OOXO}m��CD�@�0ʛ)���H�UK�LM-10�iA 890?�9�0;��F;�M61�C D�:�CP��1

\&V�1	�6F� �CW�9)A7Y	(R�_��_�_�_�_�\���0i^�oOUO>o Po#G�/���o'o�o��o�o�oB�0ƐrtAA�0* C @�Bu&Xw?���ju�bH0{UzAF?@ F�`�r� �o�����+�� O�:�s��mBqrr����������B�͏b�� ��7�"�[�F�X���|� ����ٟğ���N��� AO�0�B�CU
L���xE�jqBq=��Ҕ��$G@�@pϯ BȆ��G�I
E�0E�L_DEFAUL�T  �T���E��MI�POWERFL � 
E*��7�WF�DO� *��1E�RVENT 1����`(�� L�!DUM_EI�P��>��j!AF_INE�¿C�O!FT�����r�!o:� ���a�!RPC_M'AINb�DȺPϭ�Nt�VIS}�Cɻ�����!TP��PU��ϫ�d��E�!
P�MON_PROX	YF߮�e4ߑ��_��f����!RD�M_SRV�߫�g��)�!R�IﰴYh�u�!
v�M���id���!RL�SYNC��>�8|���!ROS��4��4��Y�(�}��� J�\����������� ��7��["4F� j|����!��Eio�ICE_�KL ?%� �(%SVCPRG1n>���3��3���4//�5./3/�6V/[/��7~/�/��D�/�9�/�+�@��/�� #?��K?��s?�  /�?�H/�?�p/�? ��/O��/;O��/ cO�?�O�9?�O� a?�O��?_��?+_ ��?S_�O{_�)O �_�QO�_�yO�_� �Os����>o�o }1�o�o�o�o�o�o�o ;M8q\� �������� 7�"�[�F��j����� ��ُď���!��E� 0�W�{�f�����ß�� �ҟ���A�,�e� P���t��������ί��y_DEV ���MC:���_!�OU�T��2��RE�C 1�`e�j�; �	 ������˿���ڿ��
 �`e���6�N�<� r�`ϖτϦ��Ϯ��� ����&��J�8�n߀� bߤߒ��߶������� "��2�X�F�|�j�� ������������� .�T�B�x�Z�l����� ��������,P >`bt���� ��(L:\ �d����� / �$/6//Z/H/~/l/ �/�/�/�/.��/?�/ 2? ?V?D?f?�?n?�? �?�?�?�?
O�?.O@O "OdORO�OvO�O�O�O �O�O�O__<_*_`_ N_�_�_x_�_�_�_�_ �_oo8oo,ono\o �o�o�o�o�o�o�o �o "4jX�� �������� B�$�f�T�v������� �����؏��>�,��b�P�r���p�V 1��}� P
�ܟ� yA��TYPE\���HELL_CF�G �.�F�͟ � 	�����RSR������ӯ���� ���?�*�<�u�`�������������_�  �%Ϡ3�E��Q�\����M�o�p��d��2���d]�K�:�HK ;1�H� u��� ����A�<�N�`߉� �ߖߨ������������&�8��=�OMM� �H���9�FT?OV_ENB&��1�OW_REG_�UI���IMWA�IT��a���OU�T������TIM������VAL|����_UNIT���K�1�MON_AL�IAS ?ew� ( he�#���� ����������); M��q����d ��%�I[ m�<���� ��!/3/E/W//{/ �/�/�/�/n/�/�/? ?/?�/S?e?w?�?�? F?�?�?�?�?�?O+O =OOOaOO�O�O�O�O �OxO�O__'_9_�O ]_o_�_�_>_�_�_�_ �_�_�_#o5oGoYoko o�o�o�o�o�o�o�o 1C�ogy� �H����	�� -�?�Q�c�u� ����� ��ϏᏌ���)�;� �L�q�������R�˟ ݟ�����7�I�[� m��*�����ǯٯ� ���!�3�E��i�{� ������\�տ���� �ȿA�S�e�wω�4� �Ͽ����ώ����+� =�O���s߅ߗߩ߻� f�������'���K� ]�o���>������ ����#�5�G�Y���}���������n��$�SMON_DEF�PRO ������ �*SYSTEM*  d=���RECALL ?�}�� ( �}���>Pbt��  ,����� ;M_q��(� ���//�7/I/ [/m//�/$/�/�/�/ �/�/?�/3?E?W?i? {?�? ?�?�?�?�?�? O�?/OAOSOeOwO�O O�O�O�O�O�O__ �O=_O_a_s_�_�_*_ �_�_�_�_oo�_9o�Ko]ooo�o�o&d&c�opy mc:d�iocfgsv.�io md:=>�inspiron:2260�o�o�o�	n0�bfrs:�orderfil�.dat vir�t:\temp\@�o`r��)a(.v*.dBTxW����k
xyzra?te 61 �� �n�����%e.�O}@H�Z�����"h3.~@xmpbackNpb�t����� }*�cdb�p*C�U�Y������!i.x.�:\ ��8�R�ݟn�����%e/.�a6�H�Z�_�� ��'���˯ݯn����������3400  H�Z�����"�4��� ��a�sυϗϪ�EϽ� Y�����ߡ�.�@U�992 ��o߁ߓ�&d'�H�Z�V����� ��0�����e�w��n��W�G�Y������!i2.�@�O�`�r�����)a)��I���X����� �-.�A�T� ��m�$���G�� ]� %�7����� l~�������Y� �/!3�Wh/z/ �/��B/��/�/
? /ASd?v?�??��H?��?�?OO ��$SNPX_A�SG 1�����9A� �P 0 '%�R[1]@1.Y1O �?�#�%dO �OsO�O�O�O�O�O�O  __D_'_9_z_]_�_ �_�_�_�_�_
o�_o @o#odoGoYo�o}o�o �o�o�o�o�o*4 `C�gy��� ����	�J�-�T� ��c�������ڏ��� ��4��)�j�M�t� ����ğ������ݟ� 0��T�7�I���m��� �����ǯٯ���$� P�3�t�W�i������� �ÿ����:��D� p�Sϔ�wω��ϭ���  ���$���Z�=�d� ��sߴߗߩ�������  ��D�'�9�z�]�� ��������
���� @�#�d�G�Y���}��� ����������*4 `C�gy��� ���	J-T �c������ /�4//)/j/M/t/ �/�/�/�/�/�/�/?�0?4,DPARAM� �9ECA ��	��:P�4��0$HOFT_K�B_CFG  �p3?E�4PIN_S_IM  9K�6��?�?�?�0,@RVQSTP_DSB�>��21On8J0SR ���;� & �=O{Op0�6TOP�_ON_ERR � p4�9�APT�N �5�@�A�BRINGo_PRM�O J0�VDT_GRP �1�Y9�@  	 �7n8_(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2Dkhz��� ����
�1�.�@� R�d�v���������Џ �����*�<�N�`� r���������̟ޟ� ��&�8�J�\����� ������ȯگ���� "�I�F�X�j�|����� ��Ŀֿ����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�tߛߘߪ߼����� ����(�:�a�^�p� ����������� � '�$�6�H�Z�l�~���������������3VP�RG_COUNTƛ6��A�5EN�B�OM=�4J_�UPD 1��;8  
p2�� ���� )$6 Hql~���� �/�/ /I/D/V/ h/�/�/�/�/�/�/�/ �/!??.?@?i?d?v? �?�?�?�?�?�?�?O OAO<ONO`O�O�O�O �O�O�O�O�O__&_ 8_a_\_n_�_�_�_YSDEBUG" ʇ �Pdk	�PSP�_PASS"B�?�[LOG �V�m�P�Xξ_  �g�Q
�MC:\d�_b_MPCm��o�o��Qa�o �vfSA/V �m:dUb��U\gSV�\T�EM_TIME �1�� (�P@�TNu]qT1SV�GUNS} #'�k�spASK_OPTION" �g�ospBCCFGg ��| �b��z`����4� �X�C�|�g�����ď ֏������	�B�-� f�Q�c���������� ϟ��,�>�)�b��YR���S���ƯA��� ��� ��D��nd��t 9�l���������ڿȿ �����"�X�F�|� jϠώ��ϲ������� ��B�0�f�T�v�x� ���ߦؑ������� (��L�:�\��p�� ���������� �6� $�F�H�Z���~����� ��������2 V Dzh����� ����4Fdv ������/ /*/�N/</r/`/�/ �/�/�/�/�/�/?? 8?&?\?J?l?�?�?�? �?�?�?�?�?OO"O XOFO|O2�O�O�O�O �OfO_�O_B_0_f_ x_�_X_�_�_�_�_�_ �_oooPo>otobo �o�o�o�o�o�o�o :(^Lnp� ����O��$�6� H��l�Z�|�����Ə ؏ꏸ����2� �V� D�f�h�z�����ԟ ����
�,�R�@�v� d���������ίЯ� ��<��T�f����� ��&�̿��ܿ��&� 8�J��n�\ϒπ϶� �����������4�"� X�F�|�jߌ߲ߠ��� ��������.�0�B� x�f��R��������� ���,��<�b�P��� ����x��������� &(:p^�� ����� 6 $ZH~l��� �����/&/D/V/ h/��/z/�/�/�/�/��&0�$TBCS�G_GRP 2���%� � �1 
 ?�  /?A?+?e?O? �?s?�?�?�?�?�;2�3�<d, ��$A?1	 HC{���6>��@E~�5CL  B�'2�^OjH4J��B�\)LFY  A��jO�MB��?�IBl��O�O�@�JG_�@�  D	�15_ __�$YC-P{_F_`_j\��_�]@0�>�X�Uo �_�_6oSoo0o~o�o��k�h�0	V�3.00'2	mw61c�c	*�`0�d2�o�e>�JC0(�a�i ,p�m-w  �0����o�mvu1JCFG [��% 1 #0vz��rBr�|�|����z� � %��I�4�m�X���|� �������֏���3� �W�B�g���x����� ՟��������S� >�w�b�����'2A �� ʯܯ������E�0� i�T���x���ÿտ� �����/��?�e�1 �/���/�ϜϮ����� ���,��P�>�`߆� tߪߘ��߼������ ��L�:�p�^��� ���������� �6� H�>/`�r�������� �������� 0V hz8����� �
.�R@v d������� //</*/L/r/`/�/ �/�/�/�/�/�/�/? 8?&?\?J?�?n?�?�? �?�?���?OO�?FO 4OVOXOjO�O�O�O�O �O�O__�OB_0_f_ T_v_�_�_�_z_�_�_ �_oo>o,oboPoro to�o�o�o�o�o�o (8^L�p� ������$�� H�6�l�~�(O����f� d��؏���2� �B� D�V�������n���� ԟ
���.�@�R�d�� ��v��������Я� ��*��N�<�^�`�r� ����̿���޿�� $�J�8�n�\ϒπ϶� ��������ߊ�(�:� L���|�jߌ߲ߠ��� �������0�B�T�� x�f���������� ����,��P�>�t�b� �������������� :(JL^�� ���� �6 $ZH~l��^� ��dߚ //D/2/ h/V/x/�/�/�/�/�/ �/�/?
?@?.?d?v? �?�?T?�?�?�?�?�? OO<O*O`ONO�OrO �O�O�O�O�O_�O&_ _6_8_J_�_n_�_�_ �_�_�_�_�_"ooFo ��po�o,oZo�o�o �o�o�o0Tf x�H����� ��,�>��b�P��� t���������Ώ�� (��L�:�p�^����� ��ʟ���ܟ� �"� $�6�l�Z���~����� دꯔo��&�ЯV� D�z�h�������Կ¿ ��
��.��R�@�v�8dϚτ�  ����� �������$�TBJOP_GR�P 2ǌ���  ?�������������xJ�BЌ��9� �<� �X����� @���	 ��C�� t�b  �C����>��1͘Րդ�>̚й���33=�C�Lj�fff?��?�ffBG��ь������t�ц�>��(�\)�ߖ�E����;��hCY�j��  @h��B�  A����f�~��C�  Dh�8��1��O�4�N�����
:���Bl^��j�i�l�l�����Aə�A��"��D��֊=qqH���нp�h���Q�;�A}�j�ٙ�@L��D	2�������$�6�>B�\��T���Q��tsx�@33@���C���y�x1����>��Dh�����������<{�h�@i�  ��t��	��� K&�j�n| ���p�/�/(:/k/�ԇ���!��	V3.00J��m61cI�*� IԿ��/�' �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I��!CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;��;Q�T,8�4` *�ϴ?�2���3\�X/O���ESTPARS c ��	���HR@ABLE 1���I�0��
H�7 8��9
G
H
H����*
G	
H

H
HYE���
H
H
HN6FRDIAO�XO@jO|O�O�O�ETO"_�4[>_P_b_t_�^:BS _� �JGoYoko}o �o�o�o�o�o�o�o 1CUgy�� ��`#oRL�y�_�_�_ �_�O�O�O�O�OX:B~�rNUM  �ū�P��� �V@P:B_CFG �˭�Z�h�@��IMEBF_TT%ApU��2@�VERS��q��R 1̞��
 (�/����b� ����J�\��� j�|���ǟ��ȟ֟� ����0�B�T���x��������2�_���@��
��MI_CH�AN�� � ��DOBGLV����������ETHERA�D ?��O��������h�����R�OUT�!��!�������SNMA�SKD��U�25�5.���#�����O�OLOFS_DI�%@�u.�ORQC?TRL ����� }ϛ3rϧϹ������� ��%�7�I�[�:����h�z߯�APE_D�ETAI"�G�PON_SVOFF=����P_MON ��֍�2��STRTCHK �^������VTCOM�PAT��O�����FPROG %^��%  BCKED�T-Q��9�PLA�Y&H��_INST+_Mް �������US�q��LCK����QUICKM�E�=���SCRE�Z�G�tps� ���u�z�����_��@@n�.�SR_�GRP 1�^�/ �O���� 
��+O=sa�쀚�
m���� ��L/C1g U�y����� 	/�-//Q/?/a/�/�	123456�7�0�/�/@Xt�1����
 �}i�pnl/� gen.htm�? ?2?�D?V?`Pan�el setupZ<}P�?�?�?�?�?�? �??,O>OPO bOtO�O�?�O!O�O�O �O__(_�O�O^_p_ �_�_�_�_/_]_S_ o o$o6oHoZo�_~o�_ �o�o�o�o�o�oso�o 2DVhz�1 '���
��.�� R��v���������Џ|G���UALRM��oG ?9� � 1�#�5�f�Y���}��� ����џן���,���P��SEV  �����ECFG ��롽��A�� ��Ƚ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �(�� ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1�����(�:�� ����962�߆��`���K�]�o�36u� 
��.�@���W�i�{� ��������R����� /A��ew�� ��N��+ =O�s��������f��f// '/9/K/]/`�/�/�/ �/�/�/j/�/?#?5? G?Y?�/�/�?�?�?�? �?�?x?OO1OCOUO gO�?�O�O�O�O�O�O tO�O_-_?_Q_c_u_ _�_�_�_�_�_�_� �)o;oMo_oqo�o�_ �o�o�o�o�o�o% 7I[m� � ������3�E� W�i�{������ÏՏ �������A�S�e� w�����*���џ��� ��ooO�a�s��� ������ͯ߯��� '���K�]�o������� ��F�ۿ����#�5� ĿY�k�}Ϗϡϳ�B� ��������1�C��� g�yߋߝ߯���P��� ��	��-�?�*�<�u� ������������ �)�;�M�������� ��������l�% 7I[����� ��hz!3E Wi������ �v////A/S/e/�P���$UI_P�ANEDATA �1�����!�  	�}w/�/�/�/�/?? )?>?��/i?{? �?�?�?�?*?�?�?O OOAO(OeOLO�O�O �O�O�O�O�O�O_&Y� b�>RQ?V_ h_z_�_�_�__�_G? �_
oo.o@oRodo�_ �ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_� �!�3�E�W��{��_ ����ÏՏ���`�� /��S�:�w���p��� ��џ������+�� O�a���������ͯ ߯�D����9�K�]� o��������ɿ��� Կ�#�
�G�.�k�}� dϡψ����Ͼ���n� ��1�C�U�g�yߋ��� ����4�����	��-� ?��c�J����� �����������;�M� 4�q�X��������� ��%7��[�� �����@� �3WiP� t�����/� //A/����w/�/�/�/ �/�/$/�/h?+?=? O?a?s?�?�/�?�?�? �?�?O�?'OOKO]O DO�OhO�O�O�O�ON/ `/_#_5_G_Y_k_�O �_�_?�_�_�_�_o o�_Co*ogoyo`o�o �o�o�o�o�o�o-�Q8u�O�O}���������) �>��U-�j�|����� ��ď+��Ϗ��� B�)�f�M��������� �����ݟ�&�S�K��$UI_PAN�ELINK 1��U  ��  ��}�1234567890s���������ͯ դ�Rq����!�3�E� W��{�������ÿտDm�m�&����Qo�  �0�B�T�f�x� �v�&ϲ��������� ߤ�0�B�T�f�xߊ� "ߘ����������� ��>�P�b�t���0� ������������$� L�^�p�����,�>�������� $�0, &�[gI�m�� �����>P 3t�i��Ϻ � -n��'/9/K/]/ o/�/t�/�/�/�/�/ �/?�/)?;?M?_?q? �?�UQ�=�2"��? �?�?OO%O7O��OO aOsO�O�O�O�OJO�O �O__'_9_�O]_o_ �_�_�_�_F_�_�_�_ o#o5oGo�_ko}o�o �o�o�oTo�o�o 1C�ogy��� ��B�	��-�� Q�c�F�����|����� ��֏�)��M�� �=�?��?/ȟڟ� ���"�?F�X�j�|� ����/�į֯���� �0��?�?�?x����� ����ҿY����,� >�P�b��ϘϪϼ� ����o���(�:�L� ^��ςߔߦ߸����� ��}��$�6�H�Z�l� �ߐ���������y� � �2�D�V�h�z�� ��-���������
�� .RdG��} ����c���< ��`r����� ���//&/8/J/� n/�/�/�/�/�/7�I� [�	�"?4?F?X?j?|? ��?�?�?�?�?�?�? O0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�__�_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o ��6H�l ~a������ ��2��V�h�K��� ����1�U
�� .�@�R�d�W/������ ��П������*�<� N�`�r��/�/?��̯ ޯ���&���J�\� n�������3�ȿڿ� ���"ϱ�F�X�j�|� �Ϡϲ�A�������� �0߿�T�f�xߊߜ� ��=���������,� >���b�t����� +������:�L� /�p���e��������� �� ��6����ۏ��$UI_Q�UICKMEN � ����}��RESTO�RE 1٩��  � 
�8m3\ n���G��� �/�4/F/X/j/|/ '�/�/�//�/�/? ?0?�/T?f?x?�?�? �?Q?�?�?�?OO�/ 'O9OKO�?�O�O�O�O �OqO�O__(_:_�O ^_p_�_�_�_QO[_�_ �_I_�_$o6oHoZolo o�o�o�o�o�o{o�o  2D�_Qcu �o������� .�@�R�d�v�������Џ⏜SCRE�� ?�uw1sc� u2�U3�4�5�6��7�8��USE�R����T���k�s'���4��5��6ʆ�7��8��� ND�O_CFG ڶ�  �  � P�DATE h��None��SEUFRAME�  ϖ��R�TOL_ABRT8����ENB(��?GRP 1��	�Cz  A�~� |�%|�������į֦!��X�� UH�X�~7�MSK  K�4S�7�N�%uT��%�����VISCAND_MAXI��I�3���FAI�L_IMGI�z ��% #S���IMRE/GNUMI�
���gSIZI�� �ϔ�,�ONTMOiU'�K�Ε�&�����a��a���s�FR:�\�� � �MC:\(�\LO�Gh�B@Ԕ !�{��Ϡ�����z? MCV����oUD1 �EX	��z ��PO64�_�Q��n66��PO!�LI�O�䞶e�V�N�f@�`�I�� =	_�S�ZVmޘ��`�W�AImߠ�STAT' �k�% @��4�F�T�$#�x �2�DWP  ���P G��=���͎���_JMPERR 1ޱ�
  �p2345?678901�� �	�:�-�?�]�c��� ��������������$�MLOW�ޘ���Ό�_TI/�˘'���MPHASE � k�ԓ� ��SoHIFT%�1 Ǚ��<z��_ ����F/ |Se����� ��0///?/x/O/ a/�/�/�/�/�/�����k�	VSFT]1\�	V��M+3� �5�Ք p��~��A�  B8[0[0�Πpg3a1Y21�_3Y�7ME��K��͗	6e���&%�J�M���b��	���$��TDINE#ND3�4��4OH�+�G1�OS2OIV I����]LRELE�vI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�YBOX �ǝf_\��b�2�TI190.0.�P�83p\�V25�4p^�Ԓ	 ��S�_�[b���robot84q_ ?  p�9o\�pc�PZoMh��]Hm�_Jk@1�o�ZWABCd��k�,�� �P\�Xo}�o0) ;M�q����@����>��aZ�b��_V