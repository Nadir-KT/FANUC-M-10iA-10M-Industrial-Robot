��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �)(�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�:  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"�SBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�� W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2����AXD�#
 �d $CARD�_EXIST4�$FSSB_TY�PuAHKBD_YS�B�1AGN Gn� $SLOT�_NUMJQPREV,DBU� g1� �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��AETE_OK�RUS�P_CR�Q$;4�V� 0LACIw1�RAP�k �1x@ME@$D�V�Q�Pv�Ah{oQL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa�!ip;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I�9�TY�D,P*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6���7��8��94�ACO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS�`�}Aw��"�tP_*0wOFSzR @� �RO_K8���aIT<�3��NOM_�0�1�ĥ3��TC �� $���AxP��K}EX�� �0g0I0x1��p�
$TFa�ކC$MD3��TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF�vF��40CPp@�a2 6
P$A`PU�3N�)#�dR*�AqX�!sDETAI�3�BUFV��p@1c |�p۶�pPIdT�� PP[�MZ�M�g�Ͱj�F[�SIMQSI�"0��A.���9��lw Tp|z�M��P�B�FAC5TrbHPEW7�P1�Ӡ��v��MCd�k �$*1JB�p<�*1DECHښ�H���(�c� � ~+PNS_EMP��G$GP���,P_���3�p�@Pܤ��TC ��|r��0�s��b�0��� �B���!
���JR|� ��SEGFR���Iv �aR�TkpN&S,�PVF���� &k�Bv�u �cu��aE�� !2��+�8MQ��E�SIZ�3�����T��P�����aRSINF����Ӏkq��������LpX�����F�CRCMu�3CClpG��p��� O}���b�1�������T2�V�DxIC��C����r����P��{� E�V �zF_��FR�pNB0�?���8���A�! �r� Rx����V�lp�2��aPR�t�,�g:�qRTx #�5�5H"2��uAR���`CX�'$LG�p��B�1 `s�P�t�aA�0{�Уb+0R���tME�`0!BupCrRA 3tCAZ�л�pc�OT�#FC�b�`�`FNp��8�1��ADI+�a %��b�{��p$�pSp�c�`S�P��a,Q�MP6�`Y�3��M�'�pU��aU � $>�TITO1��S�S�!��$�"0�D�BPXWO��!���$SK��FD�B�"�"@�PR8� 
� ���g# >�q1$��S$��+�L9$?H(�V�%@?R4C9&_?R4ENE��c'~?(�� RE�p�Y2(H �O�S��#$L�3$$@3R��;3�MVOks_D@!V�ROScr�r�w�S���CRIG7GER2FPA�S��>7�ETURN0B�c�MR_��TUː\[��0EWM%���cGN>`��RLA���Eݡ�P�&$�P�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWA�YRMO#�aw!�� CS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�o 
CdSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc �@Sp�i�a+ �j�f���ΰAPIx2,��$1F�b�$ѐOT�@A� $DUMMAY��Ft��Ft±� |6U- ` !�HE�|s��~bc�B�@ SUFFI���4PCA�Gs5rCw6dr�!MSWU�. 8!�KEYI��5�TM�1�s�qoA&�vINޱ�D, �/ D��HOST�P!4���<���<�0°<��p<�EM'����Z�� SBL� UL>��0  �	�����DT�01� � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0QSp�����#��SAV� ����c�S< 9�`�f�P$�0E!� YN�_B�#2 0�`D�I�d�pO|�m��#�$F�R_IC� �ENC2_Sd3  ��< 3�9���� cgp����!4�"��2�A��ޖ5���`ǻ�@�Q@K&D-!�a�AV�ER�q����DSP
���PC_�q��"��|�ܣ�VALU�3�HE�(�M�I�P)���OPPm ��TH�*��SH" T�/�Fb�;�d�����d D�q�16� H(rLL_DU ǀ�a�@��k���֠�OT�"U�/����R_NOAUT5O70�$}�x�~�@s��|�C� ���C� 2iaz�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|�8p�����9 <���z�ΓKI����H猡�BaFEq@{@:� ,��&a? �P_P?��>�����E�@��v�QQ���;fp$TP�$VARI����,�7UP2Q`< W�߃TD��g���`������%���BAC�"=# T2����$)�,+r8³�p IFI��p��� q M�P"�F�l@``>t ;h��6����ST� ���T��M ����0	��i���F����������kRt ����FOR�CEUP�b܂FL+US
pH(N��� ���6bD_CM�@E �7N� (�v�P��REM� Fa���@j���
K�	N���EFF/���@3IN�QOV���OVA�	TROV� DT)��DTMX:e �P:/���Pq�vXpCL�N _�p��@ ��	_�|��_T: �|�J&PA�QDI����1��0�Y0RQDm�_+qH���M���CL�d#�RIV�{�ϓN"EAR/�I�O�PCP��B�R��CM�@N 1b =3GCLF��!�DY�(��a�#5T��DG���� �%�r�SS� )�? PP(q1�1�`_1�"811�EC13zD;5D6�GRA�J��@�����PW��ON2EBUG��S�2���gϐ_E� A ��@a� �TERM�5B<�5 �ORIw�0yC�5���SM_-`T���0D�:A�9E�5����UP��F�� -QϒA��P�3�@B$SEG�GJ� EL�UUSE.PNFI��pBx���1@��4>DC$UF�P��$���Q�@"C���G�0T������SNSTj�PATxۡg��APTHJ�A�E*�Z%qB\`F�{E��F�q�pARxPY�aSHFT͢qA�AX_SHOR$�>��6% @$GqPE���GOVR���aZPI@P�@$U?r *aAYLO���j�I�"��A8ؠ��ؠERV��Q i�[Y)��G�@R��i�e��i�R�!P�uA�SYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C��%UP���P���WORڒ@M��k0SM5T��G��GR��3�aPA�@��5�'�_H � j�A�'TOCjA7pP]Pp$OPd�O��C��%�p�O!��R%E.pR�C�AO�?��Be5pR�EruIx|'QG�e$PWR) 3IMdu�RR_$s��\5��B Iz2H8��=�_ADDRH�H_LENG�B�q�qT:�x�R��So�J.�SS��SK�����0� ��-�SE*��ھrSN�MN1K�	�j�5�@r�֣O�L��\�WpW�Q�>pACRO�p���@H �����Q� ��OUPW3�b_>�I��!q�a1��������|�� ������-���:���ViIOX2S=�D��e��]���L $x��p�!_OFF[r�_�PRM_�^�aTTP_�H��wM (�pOBJ�"l�pG�$H�LE�C���ٰN � \9�*�AB_�T��b
�S�`�S��LV���KRW"duHITC�OU?BGi�LO�q����d� Fp�k�GpSS� ���HQWh�wA��O.��`�INCPUX2VISIO��!��¢.��á<�á-� �IO�LN)�P 87�R�'�[p$SL�b�d PUT_��$�dp�Pz �� F�_AS2Q/�$ALD���D�aQT U�0�]P�A���0��PH�YG灱Z���4�UO� 3R `F���H�@Yq�Yx�ɱvpP�S�dp���x��ٷZ ��UJ��S����N�E�WJOG�G �D{IS��$�KĠL��3T |��AV���`_�CTR!S^�FgLAGf2H�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_<��Dq �LN?���V��EE!2�C�D��n�U�����`L��n��DAU��EA��0Ġt����GHr���I�BOO)�WL3 ?`�� ITV����0\�REC�SCRf 0�a�D^�����MARG��`!P�)� T�/ty�?I�S�H��WW�I���T�JGM���MNCH��I�F�NKEY��K��PRG��UF��P��FWD��HL�STP��V��@�����RSS�H�` �Q�C�T1�ZbT�R ���U�����|R��t�i�2��G��8PPO��6��F�1�M��FOCU���RGEXP�TU%I��IЈ�c�� n��n����ePf����!p6�eP7�N���CA�NAI�jB��VAI�L��CLt!;eDCS_HI�4�.��O�|!�S �Sn�8��_BU�FF1XY��PT�$�� �v��f�QL6q1YY��Pp �����pOS1�%2�3���_�0Z �  ��aiE��*��IDX�dP��RhrO�+��A&S�T��R��Yz�<! _Y$EK&CK+����Z&m&KF�1[ L��o�0��]PL� 6pwq�t^����w��7�?_ \ �`�Р瀰�7��#�0C��]{ ��CLDP��>;eTRQLI�jd8.�094FLGz�0�r1R3�DM�R7��LqDR5<4R5ORG.� ��e2(`���V�8.��T8<�4�d^ �q�<4(��-4R5S�`T00m���0DFRCLM�C!D�?�?3I@��M9IC��d_ d����RQm�q�DSTB	�  �Fg�H�AX;b �H�LE�XCESZr�rBMup�a`��B;d���rB`��`a��F_�A�J��$[�O�H0K��db \��ӂS�$�MB��LIБ}SREQUIR�R>q�\<Á�XDEBU��oAL� MP�c�ba��Ph؃ӂ!BoAND�ф�`�`d�҆�c�cDC1��IN�����`@�(h?Nz�@q��o��R�QPST8� �e�rLOC�RI,�p�EX�fA�p���AoAODAQP�f� X��ON��[rMF�����f)�"I��%��e��T���FX�@I�GG� g ��q��"E�0��#���$R�a%;#7y��Gx��xVvCPi�DATAw��pE:�y��RFЭ�N�Vh t $MD�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?�uD�)�b�	@nÐi �@CU��qV�T0�eRR2Ňj Dɐ�Qނ�Bd�$CALI�@F�Gt�s�2�RIN��:v�<��NTE����kE���,��b����_Nl��ڂ��kDׄ�Rm�DIViFD�H�@ـn�$�V��'c!$��@������~�[���oH �$B�ELTb��!ACC�EL+��ҡ��ICRC�t����T/!���$PS�@#2L��q�Ɣ83������<� ��PATH����D����3̒Vp�A_� Q�.�4�B�Cᐈ��_MGh�$DDxQ���G�$FWh���p��m�����b�DE���PPABNԗR?OTSPEED����00J�Я8��@��~��$USE_�2�P��s�SY��c�ZA kqYNu@Ag���OFF�q�MO�UN�NGg�K�OL�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I(���4�\B�ݠVEO�w�Ͳ23�_UPE�߳LOWL���00����D���BwP��� �1RyCʀƶMOSIV��JRMO���@GPE�RCH  �OV ��^��i�<!�ZD <!�c��d@�P��!V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�(��<�1Ӣ`0 ��RTI$Qx�0 MO���МB@ R�0J��D��s�H�x���b�DUM2(��S_BCKLSH_C(���>�=�q�#��U��ԑ���2�t�]ACLALvŲ�1n�PN�CHK00'%SD�RTY4�k��y�1r�q_6#2�_UM$Prj�Cw�_�SCL���ƠLMT_J1_�LO��@���q��E������๕�幘S�PC��7������P	Co���H� �PU�m�C/@�"XT_�c�C�N_��N��e���S	Fu���V�&#�����9�(���=�C�u�SH6#��c����1�Ѩ��o�0�͑
��_�PALt�h�_Ps�W�_10���4�R�01D�VG�Jb� L�@J�OGW����TORQU��ON*�Mٙ�sRHљ�&�_W��-�_=��PC��I��I�I�%II�F�`�JLA.,�1[�VC��0�D�B�O1U�@i�B\J�RKU��	@DBOL_SMd�BM%`�_DLC�BGRV���C��I��H_p� �*COS+\�(LN�7+X>$ C�9)I�9)u*c,)b�Z2 HƺMY@!̳( "TH&-�)TH�ET0�NK23�I��"=�A CB6CB=�C�A�B(261C�616SBC�T25'GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t���B�6���AQ|r�f$NE�DpIB U�\B$5��$!��!A�%Ep(G%(!LPH$U�2׵�2SXpCc%pC�r%�2�&�C�J�&!�V�AHV6H3�YLVhJV�uKV�KV�KV�KV
�KV�IHAHZF`RXM���wXuKH�KH�KH��KH�KH�IO2LORAHO�YWNOhJOuKUO�KO�KO�KO�KO�&F�2#1ic%�d�4GSPBALANgCE_�!�cLEk0H_�%SP��T&�b�c&�br&PFULC��hr�grr%Ċ1k�y�UTO_?�jTg1T2Cy��2N&� v�ϰctw�g�p�0Ӓ~���T��O���� �INSEGv�!�R�EV�v!���DIF���1l�w�1m�
�OB�q
����M�Iϰ1��LCHW3AR����AB&u�?$MECH,1� X:�@�U�AX:�P��pY�G$�8pn 
Z���|���ROBR�C�R(���N�(��MSK_�`f�p WP Np_��R����΄ݡ�1��ҰТ`΀ϳ��΀"�IN�q��MTCOM_�C@j�q  �L��p��$NOR�E³5���$�r� 8� GR�E�S�D�0ABF�$XYZ_DA5A���DEBU�qI��Q��s �`$�COD��� ��k�F��f�$BUFIN�DXР  ��M{OR��t $-�U��)��r�B���(�����Gؒu � $SIMULT ৐~�� ���OBJ�E�` �ADJUS<>�1�AY_Ik���D_����C�_FIF�=�T� ��Ұ ��{��p� �����p�@:��D�FRI��ӥMT��RO� ��E�z{�͐OPWO��ŀv0��SYS�BU�@ʐ$SOP�����#�U"��pPgRUN�I�PA��DH�D����_OUb�=��qn�$}�/IMAG��ˀ�0�P�qIM����IN��q���RGOVR!Dȡ:���|�P~���Р�0L_6p���i⦄�RB���0��ML���EDѐF� ���N`M*����'��˱SL�`ŀw �x $OVSL�vSDI��DEX�m�g�e�9w�����V� ~�N���w�����țǖȳ�M�̐ ���q<��� x HxˁE�F�ATUS�Ѕ�C�0àǒ��BSTM����If����4����(�ŀy DBˀEz�g���PE�r������
���EXE ��V��E�Y�$Ժ ŀgz @ˁ��UP{�fh�$�p��XN����9�H� �P�G"�{ h $GSUB��c�@_��|01\�MPWAI��P����LO��<�F��p�$RCVF�AIL_C�f�B�WD"�F���DEF�SPup | L�ˀ`�D�� U�UCNI��S���R`Ь��_L�pP��&*@�P�ā}��� @B�~���|��`ҲN�`�KET��y���Pԙ $�~���0SI�ZE] ଠ{���S�<�OR��FORMAT/p � F���r�EMR��y�UX8����PLI7�ā�  $�P�_SWI��Ş_�PL7�AL_ )�ސR�A��B�(0uC��Df�$Eh�[���C_=�U� � � ����~�J3�0����TWIA4��5��6��MOM������4 �B�AD��*���* PU70NR W��W �U������ A$PI �6���	��) �4l�}69��Q���c�_SPEED�PGq� 7�D�>D�����>tMt[��SAM�`痰>��MOV���$��p�5���5�D�1�$2��������{�Hip�IN?,{�F( b+=$�H*�(_$�+�+�GAMM�f�1{��$GET��ĐH�D�����
^pLIBRt�ѝI��$HI��!_��Ȑ*B6E��*81A$>G086LW=e6 \<G9�686��R��ٰ�V��$PD#CK�Q�H�_����;"��z�.%�7��4*�9� ��$IM_SRO�D`�s"���H�"�LE�BO�0\H��6@�@��U� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_�D�E��NO��C gA�Ҷ��@�$����I ��	�I� %Z[� �� RX" ��m���"�q �'"�8�Hӱ�t�W�UpS��хDM��O㵐.'}q��C�g���@ʣ����S�M��AÂ� � $sPY��$WH`'�NGp���H`��Fb`��Fb��Fb��PLM�@��	� 0h�H�{�X��	O��z�Z�eT�M���G� pS��C���O__0_B_�a��_%�� |S����@	 �v��v �@���w�v���EM��%O�fr�B��ː��ftP��P�M��QU� ��U�Q��Af�QTH�=�HOL��QHY�S�ES�,�UE���B��O#��  -�P0�|�gAQ���ʠJu���O��ŀ�ɂ�v�-�A;ӝROG��a2D�E�Âv�x_�ĀZ�INFO&���+����bȆAO�I킍 ((@SLEQ/�#�����H�o���S`c0O�0��01EZ0NU�e�_�AUT�Ab�COPY��Ѓ�{��@M��N�����1�P��
� ��RGI���f��X_�Pl�$��(���`�W��P��j@��G���EXT_CYCtbR��pr����h�_NA�c!$�\�<�RO�`~]�� � m��POR�ㅣ����SRVt�)����DI �T_l���Ѥ{��ۧ��ۧ �ۧ5٩6J٩7٩8���AS�BZ쐒��$�F6����PL�A�A^�TAR��@E `�Z��p���<��d� ,(@cFLq`h��@YNL�ꟼM�C���PW�RЍ�쐔e�DE�LAѰ�Y�pAD�#q2w�QSKI�P�� ĕ�x�O��`NT!� ��P_x���ǚ@�b�p1� 1�1Ǹ�?� �?� �>��>�&�>�3�>�=9�J2R;쐷� 4��EX� TQ����ށ�Q���[�pKFд�w�RDCIf�� �U`�X}�R��#%M!*�0�)��$R�GEAR_0IO�TJBFLG�igpERa��TC݃����>��2TH2N���O 1�b��Gq �T�0 ����Mİ��`Ib���REuF�1�� l�h���ENAB��lcTPE?@���!(ᭀ ����Q�#�~�+2 (H�W���2�Қ���"�4�F�X�j�3�қ�{��������j�4�Ҝ��
��.�@�R�
j�5�ҝu�������(����j�6�Ҟ���(:Lj�7�ҟ�o�����j�8�Ҡ��"4F^j�SMSK������a��E�A��MO[TE������@0 "1��Q�IO�5"%)I��tRd�Wi@��  �����X�gp�i�쐤��Y"$DS?B_SIGN4A�Q�i�̰C��>%S23�2%�Sb�iDEVICEUS#�R�R�PARIT�!O�PBIT�Q��O?WCONTR��QXⱓ�RCU� M�S�UXTASK�3NxB��0�$TATU�P���RS@@쐦�F�6�_�PC}�$�FREEFROMqS]p�ai�GETN@.S�UPDl�ARB���SP%0���� }!m$USA��p�az9�L�ERI�0Lf��pRY�5~"_�@�f�P�1�!�6WRK���D9�F9ХF�RIEND�Q4bU�F��&�A@TOOL�HFMY5�$LENGTH_VT���FIR�pqC�@�E<� IUFIN�R����RGI�1�A'ITI:�xGX��I6�FG2�7G1a����3�B�GPRR�DA���O_� o0e�I1RE`R�đ�3&���TC��8�AQJV�G|�.2
���F��1�!d�9Z �8+5K�+5��E�y�L0>�4�X �0m�LN�T�3Hz��89�(�%�4�3G��W�0�W	�RdD�Z��Tܳ`��K�a3d��$cV 2���1��I�1H�02K2sk3K3Jci�aI�i�a`�L��SL��R$Vؠ
�BV�EVk�]V*R��� �,6Lc���9V`2F{/P:B��PS_�E��$rr�C�ѳg$A0��wPR���v�U�cSk�� {��8���� 0���VX`�!�tX`��0P��ꁂ
�5SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V��� �S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD��<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C���:c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQkfC��30=	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�qG �X��ȑ����$.A$�1$�c1Ó���� x~�EG� ݓ��q!AR����09p>B�%��AXE���ROB��W�A4�_�-֣SY���!6��&MS�'WR���-1���STR��5�9�E�� 	5B��=QB90�@6������kOT�0o 	$�ARY8�w20����	%�FI��;�$�LINK�H��1��a_63�5�q�2XYZ"��;�q�3�@��1�2�8{0B�{D��� CFI��6G��
�{�_J��6��3a'OP_O4Y;5�Q#TBmA"�BC
�z��DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ ��@�5<:7�� +1�?0K�Mc�6�8Cb�vrb�4�ORQ��X�>8�#op�� ����wq�Uf�����T'OVE�Q��M;�@E#�UK#�UQ"�VW�Z Q�W���Tυ� ;� ���QH�!`�ҽ��U�Q��WkeK#kecXER��	GE	0��S�dAWaǢ:D���7!�!AX�rB! {q��1uy-!y �pz�@z�@z6Pz \Pz� z1v�y �y�+y�;y�Ky �[y�ky�{y��y��q�yDEBU��$����L�!º2WG`  AB!�,��S9V���� 
w��� m���w����1���1�� �A���A��6Q��\Q����!�m@��2CLAB3B�U�����So ) ÐER��>�� � $�@� mAؑ!p�PO���Z�q0w�_�_M�RAȑ� d r T�-�ERR�L�ÏTYz�B�I�qV3@�cΑTOQ�d:`L� �d2�p ��|˰[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	V FZN_wCFG_!� 4�� ?º�|�ų����@�ȲW �'����\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(����$�!s�Q�g�P{RV �HELLĥ�� 56�B_BAS�!�RSR��ԣo ��#S��[��1r�%���2ݺ3ݺ4ݺ5*ݺ6ݺ7ݺ8ݷ���ROOI䰝0�0NLK!�CAB� ���ACK��IN��T�:�1�@�@ z�m�_�PU!�CO� ��OU��P� Ҧ) ��޶���TPFWD_�KARӑ��RE�~��P��(��QU�E�����P
��CSTOPI_AL������0&���㰑�0S#EMl�b�|�M��dЛTY|�SOK�}�D�I�����(���_�TM\�MANRQ�ֿ0E+�|�$K�EYSWITCH�&	���HE
�B�EAT����E� LQEҒ���U��FO������O_HOM��O�REF�PPARz��!&0��C+�9OA�ECO��B<�rIOCM�D8׆�� ���8�` �# D�1����U��&��MH�»P�CFOR�C��� ���O}M�  � @V�T�|�U,3P� 1-��`� 3-�4��N�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��C@�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fi�7s�VP�UP}D��  ��x|�԰��YSLOǢ� � z��и� ��o�E��`>�^t��А�ALUץ����CU����wFOqID_L��ӿuHI�zI�$FILE_���t�ĳ$`�JvSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_�TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅�%L~�_Vj����ޠ�� ` �GR�OU�pD��B�N�FLIC��RE�QUIREa�EB�UA��p����2��������c��{ \��APPR��iC���
�EN��CLOe��S_M� v�,ɣ�
���7� ���MC�&����g�_MG�q�C�� �{�9���|�BRKz�NOL��|ĉ R��_LI|��Ǫ�k�J����P
���ڣ������&���/���6���6��8��q��Ə� ��8�%�xW�2�e�PATHa׀z�p�z�=�vӥ�ϰ�6x�CN=�CA����l�p�IN�UC���bq��CO�UM��YZ������qE%���2�������PAYLO�A��J2L3pR_AN��<�L��F�B��6�R�{�R_F2LgSHR��|�LOG���р��ӎ���ACRL_u�������.���9H�p�$H{���FLEX
��J>�� :�/� ���6�2�����;�M�_�F16����n��� ������ȟ��Eҟ� ����,�>�P�b�� �d�{����������H��5�T��X�� v���EťmFѯ �������&�/��A�S�e�+p�x�� � ������j�4pcAT����n�EL S �%øJ���ʰ;JE��CTR�Ѭ��TN��F&��HA_ND_VB[
�ܤpK�� $F20{�6� �rSW	�D��U��� $$Mt�h�R��08��@<b 35��^6A�p3�k��qD{9t�A�̈p��A��AA�ˆ0��U���D�˕D��P��G��IS�T��$A��$AN��DYˀ�{�g4�5D��� v�6�v��5缧�^�@��P�����#��,�5�>�D�J�� &0�_�ER!V9�SQOASYM��] ��¤��x��ݑ���_SHl�������sT�(����(�:�JA���S�pcir��_VI�#�Oh9�``V_UN!I��td�~�J���b �E�b��d��d�f��n���������uN$���D��H����3��"CqEN� �pDI��>�Obt2DpNx�� ��2IxQA�q��q��-��s �p� s����� ��/OMME��r4r�QTVpPT�P ���qe�i����P�x� ��yT�Pj� $DUMMY9��$PS_��RF�q�0$:� ps���!~q� X�����K�STs�ʰS�BR��M21_V�t�8$SV_ER�t�O��z���CLR�x�A  O�r?p? O�ր � D �$GLOB���#LO��Յ$�o��P�!SYSADR��!?p�pTCHM0 �� ,����W7_NA��/�e��os�TSR��l (:]8:m� K6�^2m�i7m�w9m� �9���ǳ��ǳ���ŕ ߝ�9ŕ���i�L� ��m��_�_�_�TDџXSCRE�ƀӚ� ��STF����}�pТ6�1] _:v AŁ� T����TYP�r�K��u�!u���O�@I�S�!��t���UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��PO�*q��D�UI_�pH>;� � 8��N�_HE
p��Q��p?RY ?���,��J�*��;�OUS>�� � @d����$BUTT��R|@���COLUM��<�u�SERVc#=��PANEv Ł� w� �PGEU�!��F��9�)$HE�LP��WRETER��)״���Q�� ����@� P�P� �IN��s�PN(ߠw v�1�����o ���LN�'� ����_��k��$H��M TEX8�#����FLAn +/RELV��D4p��������M��?,@��ӛ$����P=�USRVIEWŁ�� <d��pU�p�0NFIn i�FOsCU��i�PRILP�m+�q��TRI}P)�m�UNjp�{t� QP��XuW�ARNWu<�SRT+OLS�ݕ������O|SORN��RA�Uư��T��%��V�I|�zu� =$�PATHg���CACHLOG6�O�LIMybM���x'��"�HOST6��!�r1�R�OgBOT5���IMl�	 ��C� g!��E��L���i�VCPU_�AVAILB�O�EX7�!BQNL�(��`�A�� Q��Q �\�ƀ�  QpC����@$TOOLz6�$�_JMP�� �I�u$S�S�!$1VSHI9F��|s�P�p��6�s���R���OS�URW�pRADIz��2�_�q�h�`g! �q)�LUza�$OUTPUTg_BM��IML��oR6(`)�@TILN<SCO�@Ce� ;��9��F��T�� a��o�>�3���$��w�2u�<qV�zu9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+Z�t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2$��2���5��`�? �'��ZABCS�� � $�2��J�
�  �$$CLA}S�����A���@'@@VIRT8��O.@ABS�$��1 <E�� <  *AtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@��R�d�v�����M@[�A�XLր�&A�dC  ���IN��ā��GPRE������LARMRECOV <I䂥��NG�� \K	 =#�
J�\�M@�PPLIC�?�<E�E�H�andlingT�ool �� 
�V7.50P/2{8 *A�Hy���
�_SW�� �UP*A� ��F�0ڑ����A@��� 20��*A��:�����FB 7DA�5�� '@�Iy@����No�ne������ ���T��*A4�9xx��P_���V����g�U�TOB�ค����HGAPON8@��LAz��U��D 1<EfA�����x����� Q 1שI Ԁ��Ԑ��:�i�n����#B=)B ���\��HE�Z�r�HTTHKY��$BI�[� m�����	�c�-�?� Q�o�uχϙϫϽ��� �����_�)�;�M�k� q߃ߕߧ߹������� �[�%�7�I�g�m�� ������������W� !�3�E�c�i�{����� ����������S/ A_ew���� ���O+=[ as������ �K//'/9/W/]/o/ �/�/�/�/�/�/�/G? ?#?5?S?Y?k?}?�? �?�?�?�?�?COOO 1OOOUOgOyO�O�O�O �O�O�O?_	__-_K_Q_��(�TO4�s����DO_CLEAN���e��SNM  9� �9oKo]o�oo�o�DSPDR3YR�_%�HI��m@&o�o�o#5G Yk}����"���p�Ն �ǣ�q�XՄ��ߢ��g�PL�UGGҠ�Wߣ��P�RC�`B`9���o�=�OB��oe�SEGF��K������ o%o����#�5�m���LAP�oݎ���� ������џ������+�=�O�a���TOT�AL�.���USE+NUʀ׫ �X����R(�RG_STR�ING 1��
_�M��Sc��
��_ITEM1 �  nc��.� @�R�d�v��������� п�����*�<�N��`�r�I/O �SIGNAL���Tryout �Mode�In�p��Simula�ted�Out���OVERR~�` = 100��In cycl����Prog OAbor����ĿStatus�	�Heartbea�t��MH Fa�ulB�K�Aler Uم�s߅ߗߩ߻���p������ �S ���Q��f�x��� ������������,� >�P�b�t�������,�WOR������V�� 
.@Rdv� ������p*<N`PO�� 6ц��o���� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/�DEV�*0�? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O�qO�O�O�OPALTB��A���O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o�OGRI�p��ra�O Lo�o�o�o�o�o�o *<N`r��@����`o��RB� ��o�>�P�b�t��� ������Ώ������(�:�L�^�p����PREG�N��.���� ����*�<�N�`�r� ��������̯ޯ����&����$ARG�_��D ?	����i��  	$��W	[}�]}�������\�SBN_CONFIG i�������CII�_SAVE  ��۱Ҳ\�TCE�LLSETUP �i�%HOM�E_IO�͈�%�MOV_�2�8�R�EP���V�UTOoBACK
�ƽ�FRA:\��� �Ϩ���'�`!��������� ����$�6�c�pZ�lߙ��Ĉ���� ���������!凞�� M�_�q����2��� ������%�7���[� m��������@��������!3E$��� Jo�������WINI�@��ε���MESSAG�����q��ODEC_D$���O,0�.��PAUS�!��i� ((O l��������  /�//$/Z/H/~/�l/�/�'akTSK�  q�����UgPDT%�d0~;WSM_CF°�i�еU�'1G�RP 2h�93 �|�B��A�/S�XS�CRD+11
1; ����/�?�? �? OO$O��߳?lO ~O�O�O�O�O1O�OUO _ _2_D_V_h_�O	_|X���GROUN0|O�SUP_NAL��h�	�ĠV_E�D� 11;
 ��%-BCKED�T-�_`�!oEo%�A��a��o����Y�ߨ���e2no_˔o�o�b���ee�o8"�o�oED3�o��o ~[�5GED4�n#�� ~�8j���ED5Z���Ǐ6� ~���}���ED6����k�ڏ ~G�8��!�3�ED7��Z���~� ~�V�şןE�D8F�&o��Ů�}����i�{�ED9ꯢ�W�Ư
}3�����CRo����π3�տ@ϯ����P�PN�O_DEL�_�RGE_UNUSE�_��TLAL_OUT� q�c�QWD_ABOR� �΢Q���ITR_RTNz����NONSe����CAM_�PARAM 1��U3
 8
S�ONY XC-5�6 234567w890�H � @���?��ҟ( АV�|[�r؀~�X�HR5�k�|U�Q�߿�R57�����Aff���KOWA SC3W10M|[r�̀�d @6�|V ��_�Xϸ���V��� ����$�6��Z�l��CE_RIA_I8�57�F�1���R|]��_LI�O4W=� ��P<z~�F<�GP 1�,���_GY<k*C*  ���C1� 9� @� G�� �CLC]� d*� l� s�R� ���[�m� v� �� �� �� C��� �"�|W��7�H=EӰONFI� ���<G_PRI 1�+P�m®/���������'CH�KPAUS�  1E� ,�>/P/ :/t/^/�/�/�/�/�/ �/�/?(??L?6?\?4�?"O�����H^�1_MOR��� ��PBZ?�<���5 	 �9 O �?$OOHOZK�2	���=9"�Q?55���C�PK�D3P��|����a�-4�O__|Z
�OG_�7@�PO�� ��6_��,xV��ADB���='�)�
mc:cpmi�dbg�_`��S:�  7;�P����U�p�_)o�S  Y�C@��	f�P��_mo8j�  �׏`�Oko�o9iU�)�I)�JOkg�o��o�l�`hOkf��oGq:I�ZDEFg f8��)�R�6pbuf.txt m�]n�@����# �	`)Ж�A=L�m��zMC�21�=���9���4�=��n׾�Cz  BH�BCCPUeB���CF�;.�<C���C5�rSZE@D�nyD�Q��D��>���D�;D�����F��>�F�$G}RB�Gzր���SY��!�vqGR���Em�)�.��)�)��<�q�G�Sx2��Ң �� fa�D�j���ES\�E@EX�EQ��EJP F�E��F� G��ǎ^F E��� FB� H,-� Ge��H3Y����  >�3�3 ���xV � n2xQ@��5Y���8B� A�AST<#�
� �_'�%�~�wRSMOFS����~2�yT1�0D�E �O@b 
��(�;�"�  (<�6�z�R���?��j�C4��SZm� �W��{�m�C��B�-G�Cu�@$�q���T{�FPROG� %i����c�I���� �Ɯ�f�KEY?_TBL  �vM��u� �	
��� !"#$%�&'()*+,-�./01c�:;<=>?@ABC�p�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������p��������������������������������������������������������������!j�L�CK��.�j���ST�AT���_AUT/O_DO���W/��INDT_ENB�߿2R��9�+�T2<w�XSTOP\߿2�TRLl�LETE�����_SCRE�EN i�kcsc��U��MMENU 1 i?  <g\�� L�SU+�U��p3g�� ����������2�	� �A�z�Q�c������� ��������.d ;M�q���� ��N%7] �m���/� �/J/!/3/�/W/i/ �/�/�/�/�/�/�/4? ??j?A?S?y?�?�? �?�?�?�?O�?O-O fO=OOO�OsO�O�O�O �O�O_�O_P_Sy�_MANUAL���n�DBCOU�RI�G���DBNUM��p��<���
�QP�XWORK 1!R�ү�_oO.o@o|Rk�Q_AWAY�S���GCP ��=��df_AL�P�dbB�RY�������X_�p� 1"�� , 
�^���o xvf`%MT�I^�rl@�:s�ONTIM���&���Zv�i
õ�cMOTNEND����dRECORD �1(R�a��ua�O��q��sb�.� @�R��xZ������� ɏۏ폄���#���G� ��k�}�����<�ş4� �X���1�C���g� ֟��������ӯ�T� 	�x�-���Q�c�u��� �������>���� )Ϙ�Mϼ�F�࿕ϧ� ����:�������%�s` Pn&�]�o��ϓ�~ߌ� ��8�J�����5� � ��k����ߡ��J��� ��X��|��C�U��� �������0������	��dbTOLER7ENCqdBȺb`�L�͐PCS_C�FG )�k)wd�MC:\O L�%04d.CSVd
�pc�)sA �+CH� z�p)~����hMRC_O_UT *�[�`�+P SGN +��e�r��#�10�-MAY-20 �08:57*V27�-JANj21:�48�k P;����)~�`�pa�m��P�JPѬVERSION SV2.0.��6tEFLOGIC� 1,�[ 	�DX�P7)�PF."PROG_ENB�o\�rj ULSew �T��"_WRSTJ�NEp�V�r`dEMO�_OPT_SL �?	�es
 	R575)s7)�/�??*?<?'�$TO�  �-��?&V�_@pEX�Wd�u��3PATH ASA\�?�?O/{�ICT�aFo`-��gdse�gM%&ASTBF_TTS�x�Y^C��StqqF�PMAU� \t/XrMSWR.�i�6.|S/�Z! D_N�O0__T_C_x_�g_�_�tSBL_F�AUL"0�[3wTDIAU 16M6p��A1234567890gFP?BoTofoxo �o�o�o�o�o�o�o�,>Pb�S�pP�_ ���_s� � 0`�����)� ;�M�_�q����������ˏݏ��|)UMP��!� �^�TRp�B�#+�=�PMEfE~I�Y_TEMP9 È�3@�3A v��UNI�.(YN_?BRK 2Y)�EMGDI_ST�A�%WЕNC2_�SCR 3�� 1o"�4�F�X�fv����������#��ޑ14 ����)�;�����:ݤ5����� x�f	u�ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� �P�b�t�� ��xߞ� ����������
��.� @�R�d�v����� ��������*�<�N� ��r������������� ��&8J\n �������� "`�FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/4?,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O?�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �O�O�o�o�o
. @Rdv���� �����*�<�N� `�r����o����̏ޏ ����&�8�J�\�n� ��������ȟڟ�����H�ETMODE� 16���+ ��ƨ
R�d��v�נRROR_P�ROG %A�%��:߽�  ��TA�BLE  A�������#�L�RRS�EV_NUM  y��Q��K��S���_AUTO_?ENB  ��I��Ϥ_NOh� 7�A�{�R�  *U�������������^�+��Ŀֿ迄�H�ISO���I�}�_A�LM 18A� e�;�����+鿀e�wωϛϭϿ��_\H���  A����|��4�TCP_V_ER !A�!�����$EXTLOGo_REQ��{��V�SIZ_�Q�TOoL  ��Dz���=#׍�XT_BWD����r����n�_DI�� 9��}�z���m���STEP����4��_OP_DO����ѠFACTORY�_TUN�dG�E�ATURE :�����l�H�andlingT�ool ��  -� CEngl�ish Dict�ionary��O�RDEAA �Vis�� Mas�ter���96 �H��nalog �I/O���H55�1��uto So�ftware Update  ���J��matic �Backup��P�art&�gr�ound Edi�t��  8\ap�Cameraz��F��t\j6R��ell���LOA�DR�omm��sh�q��TI" ��cyo��
! o����pane�� �
!��tyle select��H59��nD���o�nitor��48�����tr��Rel�iab���adi�nDiagn�os"����2�2 u�al Check� Safety �UIF lg\a���hanced �Rob Serv> q ct\��lUser FrU���DIF��Ext�. DIO ��f�iA d��en]dr Err L@���IF�r��  �П�90��FCT�N MenuZ v�'��74� TP �In��fac � SU (G�=�p��k Exc�n g�3��Hig�h-Sper Sk]i+�  sO�H9 ~� mmunic!��onsg�teurh� ����V����^conn��2��{EN��Incr�stru���5.�fdKARE�L Cmd. L�?uaA� O�R�un-Ti� EnIv����K� ��+%��s#�S/W��74���License|T�  (Au* �ogBook(S�y��m)��"
�MACROs�,V/Offse6��ap��MH� �����pfa5�Mec�hStop Pr3ot��� d�b =i�Shif���/j545�!xr ��#��,K�b o�de Switc]h��m\e�!oz4.�& pro��4��g��Mul�ti-T7G��n�et.Pos Regi��z�}P��t Fun����3 Rz1��Nu!mx �����9m�1>�  Adjuj��O1 J7�7�* ��<���6tatuq1EIKRDMt�ot��scove�� ��@By- }Ouest1�$Go� �� U5\SNPX b"���YA�"Libr����#b�� �$~@h�pd]0��Jts in VCCM�����0�q  �u!��2 R�0��/I�08��T�MILIB�M J�92�@P�Acc�>�F�97�TPT�X�+�BRSQelZ0�M8 Rm��q%��692��Une�xceptr mo�tnT  CVV�P���KC����+�-��~K  II)��VSP CSXC��&.c�� e�"�� =t�@Wew�gAD Q�8bvr �nmen�@�iP�� a0y�0�pfG�ridAplay !� nh�@*�3R�1�M-10iA(B�201 �`2V" y F���scii��load��83 �M��l����Gua=r�d J85�0�maP'�L`���stua�Pat�&]$Cyc8���|0ori_ x%oData'Pqu���ch�1��g`� mj� RLJam�5����IMI De�-B(\A�cP" #�^0C  etk}c^0asswo%q.�)650�ApU��Xnt��Pven��CTqH�5�0�YELLOW BqO?Y��� Arc�0�vis��Ch�W�eldQcial44Izt�Op� ��gs�` 2@�a��p�oG yRjT1� NE�#HT� xyWb��! �p�`!gd`���p\� =P���JPN ARCP�*PR�A�� �OL�pSup̂f�il�p��J�� ��cro�670�1C~E��d��SS�pe�t�ex�$ �P� Soz7 t� ssagN5� <Q�BP:� �9 �"0�QrtQC��P�l0dpn�笔�r�pf�q�e�ppm�ascbin4p�syn�' ptx�]08�HELNC�L VIS PK�GS �Z@MB �&��B J8@I�PE GET_V�AR FI?S (�Uni� LU�OO�L: ADD�@2/9.FD�TCm���E�@DVp���`A��ТNO WTWTOEST �� V�!���c�FOR ��E�CT �a!� AL�SE ALA`�CPMO-130���� b D: HAN?G FROMg���2��R709 D�RAM AVAI�LCHECKS �549��m�VPC�S SU֐LIM�CHK��P�0x�F_F POS� F��� q8-12� CHARS�ER>6�OGRA ��Z@wAVEH�AME��G.SV��Вאn$���9�m "y�TR}Cv� SHADP��UPDAT k�0>��STATI���? MUCH ����TIMQ MOTN-003��@�OBOGUIDE? DAUGH���b8��@$tou� �@�C� �0��PATH|�_�MOVET��� R64��VMX�PACK MAY ASSERTjS޴�CYCL`�TA���BE COR �71�1-�AN��R�C OPTION�S  �`��APSwH-1�`fix��2�SO��B��XO򝡆��_T��	�i��0j���du�byz p cwa��y�٠HI������U�pb XSP�D TB/�F� \�hchΤB0���EmND�CE�06\Q��p{ smay In@�pk��L ���traff#�	� ���~1from �sysvar s�cr�0R� ��d�DJU���H�!A���/��SET ER�R�D�P7����N�DANT SCR�EEN UNRE�A VM �PD�D���PA���R�I�O JNN�0�F�I��B��GROUNנD Y�Т٠��h�SVIP 5�3 QS��DIGI?T VERS��k���NEW�� P0�6�@C�1IMAG��ͱ���8� DIx`���pSSUE�5���EPLAN J=ON� DEL���1�57QאD��CALLI���Q��m����IPND}�IMG� N9 PZ�19޴�MNT/��ES� ���`LocR HCol߀=��2�Pn� �PG:��=�M��c�an����С: �3D mE2vie�w d X��e�a1 �0b�pof �Ǡ"HCɰ�AN�NOT ACCE�SS M cpite$Et.Qs a� {loMdFlex)a�:��w$qmo G
�sA9�-'p~0��h0�pa��eJ AU�TO-�0��!ip�u@Т<ᡠIABL�E+� 7�a FPL�N: L�pl lm� MD<�VI�����WIT HOCv�Jo~1Qui�t�"��N��USB�@��Pt & rem�ov���D�vAxi�s FT_7�PG�ɰCP:�OS-�144 � h s� 268QՐOST��p  CRASH� DU��$P��W�ORD.$�LOgGIN�P��P:	��0�046 iss�ueE�H�: Solow st��c�`6����໰I�F�IMPR��SPOT:Wh4���N1�STY��0VMGqR�b�N�CAT��-4oRRE�� � 58�1��:%�R�TU!Pe -M a�SE:�@pp���AGp�L��m@al�l��*0a�OCB �WA���"3 CN�T0 T9DWro>O0alarm�ˀm0d t�M�"0�2�|� o�Z@OME�<�� ��E%  #1�-�SRE��M�st�}0g     �5KANJI5n�o MNS@�I�NISITALI�Z'� E�f�we���6@� dr�@ f�p "��SCII� L�afails� w��SYSTaE[�i��  � tMq�1QGro8�m n�@vA����&���n�0q��RWR=I OF Lk���� \ref"�
�u�p� de-rel}a�Qd 03.�0�SSchőbet�we4�IND e�x ɰTPa�DOȬ l� �ɰGi�gE�soperawbil`p l,��aHcB��@]�le�Q0cflxz�Ð���OS {����v4pwfigi GLA�$��c2�7H� la�p�0ASB� Ifz��g�2 l\c�0��/�E�� EX'CE 㰁�P���$i�� o0��Gd`]���fq�l lxt��EFal��#0��i�O�Y�n�CLOSn��SRNq1NT^��F�U��FqKP�AN�IO V7/ॠ1p�{����DB �0ء�ᴥ�ED��DE�T|�'� �bF�N�LINEb�BUG�T���C"RLIB���A��ABC J�ARKY@��� r7key�`IL���P�R��N��ITGAR
� D$�R �Er�� *�T��a�U�0��h�[�ZE V� �TASK p.vr�P2" .�XfJ��srn�S谥dIB�P	c���B/��B�US��UNN�  j0-�{��cR'���LOE�DIVS�C�ULs$cb����BW!��R~�W`P���&��IT(঱tʠ�{OF��UNEXڠ�+���p�FtE��S�VEMG3`NML� 505� D*�C?C_SAFE�P*�p �ꐺ� PET��8'P�`�F  !���IR����c i S�>� K��K�H �GUNCHG��S^�MECH��M��T*�%p6u��tP�ORY LEAKr�J���SPEg�D��2V 74\G�RI��Q�g��CTLN��TRe @�_��p ���EN'�IN�������$���r��T�3)�i�STO�A$�s�L��͐X	����q��Y� ��TO2�J m��0F<�K�����DU�S��O��3$ 9�J F�&�����SSVGN-18#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRKC�TR/"� �q\j5���_�Q�S�qINVJ0D ZO�Pݲ�� �s��г�Ui ɰ̒�a��DUAL� J�50e�x�RVO1/17 AW�TH!�Hr%�N�247%�5q2��|�&aol ���R���at�Sd�cU8���P,�LER��i�x�Q0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�cб���{�U��RO�P 2�b�pB��ITP4M��b !�AUt c0< � pl�ete�N@� �z1^qR635 (�AccuCal2zkA���I) "�(ǰ�1a\�Ps��ǐ � bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etaca2��AT���PC�`��슰�_p�.pc�!Ɗ��:�circB���5�tl��Bɵ��:�fm+�Ί�V�b��ɦ�r�upfrma.����ⴊ�xed�8�Ί�~�pedA�D ��}b�ptlib0B�� �_�rt�߄	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆�D����c�Ӳ�5�j>ʌ����tcȐ��	�r(����mm 1��T�#sl^0��T�mѡ�&#�rm3��ub Y��q�std}��pl�;�&�ckv�=�r�vaf�䊰��9�vi������ul�`�0fp�q� �.f��� d�aq; i Data� Acquisi
��n�
��T`���1�89��22� DMCM RR[S2Z�75��9 ?3 R710�o�59p5\?��T{ "��1 (D�T� nk@���������E Ƒȵ��Ӹ�et3dmm ��ER����gE��1�q\mo?۳�=(G����[(

�2�` ! ��@JMACRO���Skip/Of�fse:�a��V�4�o9� &qR662����s�H�
 6�Bq8����9Z�4_3 J77� 6�J783�o ���n�"v�R5IK�CBq2 PTLC�Zg R�3 (�s, ��������03�	зJԷ\�sfmnmc "MNMC����ҹ�%wmnf�FMC"�Ѻ0ª etmcr�� �8����� ,K�DV��   874�\prdq>,jxF0���axisH�Process �Axes e�rol^PRA
�Dp� �56 J81j�5-9� 56o6� ��l�0w�690 98� �[!IDV�1��2(8x2��2ont�0�
 ����m2���?C���etis "I�SD��9�� FpraxRAM�P� D��defB�,�G�isbasicH�B�@޲{6�� 70U8�6��(�Acw: ������D
�/,��AMOX�� ��DvE��?�;T��>Pi� RAFM';�]�!PAM�V�W��Ee�U�Q'
bU�7y5�.�ceNe� �nterfaceh^�1' 5&!54�K<��b(Devam±��/�#���/<�Tane`"DNEWE���btpdnui �A�I�_s2�d_rsCono���bAsfj|N��bdv_arFv�f�xhpz�}w��hkH9xstc��gAp�onlGzv{�ff ��r���z�3{�q'Td>pcha�mpr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�!��pcchmp]aM�P&B�� �mpe�v�����pcs���YeS�� MacKro�OD��16Q! )*�:$�2U"_,��Y�(PC ��$_;�������o��J�geg{emQ@GEMSW�|~ZG�gesndy�<�OD�ndda��Sƕ�syT�Kɓ�su^Ҋ���n�m���L��O  ���9:p'�ѳ޲��spotplusp���`-�W�l�J�s��t[�׷p�key�ɰ�$��s��-Ѩ�m���\fea;tu 0FEAWD�oolo�srn '!2 p���a�As3���tT.� (N. A.)��!e!(�J# (j�,��o�BIB�oD -�.�n6��k9�"K��u[�-�_���p� "P�SEqW����wop "sEЅ�&�:� J������y�|��O8� �5��Rɺ���ɰ[� �X�������%�(
 ҭ�q HL�0k� 
�z�a!�B�Q�"(g�Q�����]�'� .�����&���<�!ҝ_�#��tpJ�H�~Z�� j�����y������2 ��e������Z����V� �!%���=�]�͂���^2�@iRV� on��QYq͋JF0� 8�ހ�`�	(^�dQueue���X\1����`�+F1tpvtsen��N&��ftpJ0v �RDV�	f���J1 Q���v�eyn��kvstk���mp��btkcl�rq���get�����r��`k�ack�XZ�st1rŬ�%�stl��~Z�np:!�`�� �q/�ڡ6!l�/Yr$�mc�N+v3�_`� ����.v�/{\jF��� �`�Q�΋ܒ�N50 (�FRA��+��͢f?raparm��Ҁ��} 6�J643�p:V�ELSE
�#�VAR $SG�SYSCFG.$��`_UNITS �2�DG~°@�4Jgfqr��4A�@FRL-� �0ͅ�3ې���L�0 NE�:�=�?@�8�v�9~Qx304��;�B�PRSM~QA�5T�X.$VNUM_�OL��5��DJ50�7��l� Functʂ"qwAP��琉�G3 H�ƞ�kP9jQ��Q5ձ� ��@jLJ zBJ[�6N�kAP�����S��"TPPRp���QA�prna�SV�ZS��AS8Dj5k10U�-�`cr�`8 ��ʇ�DJR`jYȑH  �Qm �PJ6�a21���48AAVM3 5�Q�b0 lB�`�TUP xbJ�545 `b�`61�6���0VCA�M 9�CLI�O b1�5 ����`MSC8�
rP� R`\sSTYL MNIN�`oJ628Q  �`�NREd�;@�`SC�H ��9pDCSU� Mete�`OR�SR Ԃ�a04 �kREIOC ��a5�`542�b9 vpP<�nP�a�`�R�`�7�`�MAS�K Ho�.r7 <�2�`OCO :��r�3��p�b�p���r0�X��a�`13\mn��a39 HRM"��q�q��LCH}K�uOPLG B��a03 �q.�pH�CR Ob�pCpP�osi�`fP6 i=s[rJ554�òp'DSW�bM�D�pqR��a37 }Rjr0 L�1�s4 �R6�7���52�r5 �2�r7� 1� P6���Re�gi�@T�uF�RDM�uSaq%�4�`930�uSNB�A�uSHLB̀\�sf"pM�NPI��SPVC�J5�20��TC�`"M�NрTMIL�I=FV�PAC W�poTPTXp6.%��TELN N M�e�09m3U�ECK�b�`UFR��`��VCOR��V�IPLpq89qSX9C�S�`VVF�J��TP �q��R62]6l�u S�`Gސ~�2IGUI�C���PGSt�\ŀH863�S�q�����q�34sŁ684`���a�@b>�3 :B抂1 T��96 :.�+E�51 y�q353�3�b1 ���b31 n�jr9 ���`�VAT ߲�q75� s�F��`�sAWSyM��`TOP u��ŀR52p���a809 
�ށXY q���s0 ,b�`885�QXрOLp}�"pE�v��tp�`LCMDў�ETSS���6� �V�CPE o�Z1�VRCd3
�NuLH�h��001m2�Ep��3 f��p��4� /165C��6�l���7PR��00�8 tB��9 -2[00�`U0�pF�1&޲1 ��޲2L"����p��޲4��5 �\hmp޲6 RB�CF�`ళ�fs�8� �Ҋ��~�J�7 OrbcfA�L�8\P0C����"�32m0u��n�K�Rٰn�5 5oEW
n�9 zΊ�40 kB��3 ��6ݲ�`00iB%/��6�u��7�u���8 µ������sU0��`�t �1 05\;rb��2 E��K���j���5˰��6A0��a�HУ`:�63�`jAF�_���F�7 ڱ�݀H�8�eHЋ��cUI0��7�p��1u��8u��9 73�������D7� ��5\t�97 ��8U�Q1��2��1�1:����h��1np�"��8�(�U1��\pyl���,࿱v ��B�85E4��1V���D�4��im��1�<���$>br�3pr�4@pGPr�6 B���цp���1����1�`͵15=5ض157 �2�у62�S����1�b��2����1Π"�2L���B6`�1<cf�4 7B�5 DR���8_�B/��18�7 uJ�8 06��90 rBn�1 �(��202 0E�W,ѱ2^��2��9�0�U2�p�2��2 �b��4��2�a"RiB����9\�U2�`xw�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`ڰR,:7 �2��V�2��5���2^��a^9���qr�����n�5����5᥁"�8Ha�Ɂ}�5B���5������`UA���� ��8�6 �6 S�0��5��p�2�#�529 ��2^�b1P�5�~�2`���&P5���8��5��u�!�5\��ٵ544��5��	R�ąP nB^z�c (�4�����SU5J�V�5��1�1@^��%�����5 �b21��gA��5m8W82� rb��95N�E�5890r�: 1�95 �"�� ����c8"a��|�L (���!J"5|6��^!"�6��B�"8�`#���+�8%�6B�AM�E�"1 iC��622�Bu�6V��d� �4��84�`ANR�SP�e/S� �C�5� �6� ��� \@� �6� �V� 3t��?� T20CA�R���8� Hf� 1DH��� AOE� ��w ,K|�� �0X\�� �!64K��ԓ�rA� �1 (M-7�!/50T�[PM��P�Th:1�C�#P�e� �3�0� 5`M�75T"� �D8p�! �0Gc� u�4��i1�-710i�1� S�kd�7j�?6�:-HS,� �RN�@�UB��f�X�=m75sA*A6an���!/CB�B2.6A �0;A�C�IB�A�2�QF1�UB2:�21� /70�S� �4����Aj1�3p����r#0 B2\m*A@C��;bi"i1K��u"A~AAU� imm7c7��ZA@I�@�Df�A�D5*A�E� #0TkdR1�35Q1�" *�@�Q�1�QC)P�1 *A�5*A�EA�5B�4>\77
B7=Q�D�2H�Q$B�E7�C�D/qA	HEE�W7�_|`jz@@� 2�0�Ejc7(�`�E"l7�@7�A
1��E�V~`�W2%Q�R9\ї@0L_�#��� �"A���b��H3s=rA/2�R5nR4�7�4rNUQ1ZU�A�s\m9
1M92L2�!F!t^Y�ps� 2ci��-?�qhimQ�t  w0 43�C�p2�mQ�r�H_ �H20�Evr�QHsXBFSt62�q`s����� ��Pxq350_�*A3I)�2�d�u0X�@� '4TX�0�pa3i1A3sQ25L�c��st�r�VR1%e�q0
��j1��O 2 �A�UEiy�.�‐� �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ�� qA!Pvs� 5	15aU ���?PŅ���ဝQG9A6�zS*�7�q�b5�1����Q��00	P(��V7]u�aitE1 ���ïp?7� !?�z���rbUQRB1P�M=�Qa9��H��QQ�25L�������Q���@L��8ܰ��y0�0\ry�"R2B�L�tN  ��w� �1DV��2�qeR�5���_bx�3�X]1m1lcqP!1�a�E�Q� 5F����!5���@M-16 Q�� f���r��Q�e�� ��� PN�LT_`�1��i1��9453�p�@�e�|�b1l>�F1u*AY2�
��R8`�Q����RJ�J3�D}T� 85
Qg�/0�� *A!P�*A�Ð𫿽�Y2ǿپ6t�6=Q����Pȓ��� AQ� g�*ASt]1^u�a jrI�B����~�|I��b��yI�\m�Qb�I �uz�A�c3Apa9q� B6S��S��m����}�85`N�N�  �(M���f1����6����161��5�s`�SC��U��A�����5\set036c����10�y�#h8��a6��6��9r�2HS ���Er���W@}�a��I�lB� ��Y�ٖ�m�u�C������5�B��B��h `�F���X0���A:���C�M��AZ��@��4��6i����� e�O�- 	���f1��F ������1F�Y	���T6HL3��U66~`���Ur�dU�9D20Lf0 ��Qv� ��fjq��N� �����0v
� ��i	��	��72lqQ2�������� \chngmove.V���d���@2l_arf	�f~�� 6������9C�Z��0�~���kr41 S���0��V��t����8��U�p7nuqQ%��A]��V�1\�Qn�BJ�2W�E�M!5���)�#:�648��F�e50S�\� �0�=�PV���e�� ����E������m7shqQSH" U��)��9�!A��(����� ,Ks��ॲTR1!�L��,�60e=�4F�d����2��	 R-�� ���������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2��"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D�� �5V��@2cVE��pȖ�T��pt갖�1L ~E�#�F�Q��9E�#Dce/��RT��59�� �	�A�EiR�������9\m20�20 ��+�-u�19r4�`� E1�=`O9`�1"ae��O�2��_$W}am41�4�3�/d?1c_std��1�)�!�`_T��r�_ 4\jdg�a�q�P J%!~`-�r�+bg8B��#c300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W �"PsA��e��� �t�i�P�W.�� c�FX.�e�kE1�4�44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�A Pf��coWo!\�[2a��2A;_2��QW2�bF�(�V11ă23�`��X5�Ra2�1�J*9�a:88�J9X�l5�m1a`첚��*���(85�& �������P6����R,52&A����,8fA9IfI50\u�z��OV
�v��}E֖J0���Y>� 16r�C �Y��;��1��L���A q�&ŦP1��vB)e��m�����1p� .�1DV��27�F��KAREL Us�e S��FCTN<��� J97�FA+�� (�Q޵�p%�L)?�Vj9F?(�j�R�tk208 "Km�6Q�y�j��iæP�r�9�s#��v�kr;cfp�RCFt3����Q��kcctme��!ME�g����6�mWain�dV�� ��Cru��kDº�c��0�o����J�dt�F9 �»�.vrT�f�����E%�!��5�FR�j73B�K���UtER�HJ�O  J��# (ڳF���F�q� Y�&T��p�F�z��19�tkvBr���V�h�9p�E�y�<�k������p��;�v���"CT�� f����)�
І��)� V	�6���!��qFF ��1q���=�����O�@?�$"���$��je����TCP Aut��r�<520 H5n�J53E193��9��96�!8��9���	 �B574��5�2�Je�(�� Se%!Y�����u��ma>�Pqtool�ԕ������conr�el�Ftrol �Reliable��RmvCU!��H51������ a55�1e"�CNRE ¹I�c�&��it��l\sfutst "UTա��"X�\u��g@�i�6Q]V�0�B,Eѝ6A�  �Q�)C���X��Yf�hI�1|6s@6i��T6IU��vR�d�
$ae%1��2�C58�E6��8�Pv�iV4OFH�58SOeJ� mvBM6E~O58�I�0�E �#+@�&�F�0���F �P6a���)/++�</>N)0\tr1������P ,K�ɶ�rmwaski�msk�a$A���ky'd�h	A	��P�sDispla�yIm�`v����J887 ("A��+Hyeůצprds�ҨIϩǅ�h�0pl�2"�R2��:�Gt�@��PRD�TɈ�r�C�@�Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@��^Sp��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@�P�firmQ����P@p�2�=bk�6�r�3��6��tppl��PAL���O�p<b�ac�q 	��g1J�U�d�J��gait_9e��Y��&��Q���	�Sha�p��eratio�n�0��R674�51j9(`sGen@�ms�42-f��r�p`�5����2�rsgl��E��p�G���qF�20�5p�5S���Ձ�re�tsap�BP�O�\}s� "GCR��z�? �qngda�AG��V��st2ax�U��Aa]��bad��_�btputl�/�&�e���tpli1bB_��=�2.����5���cird�v�sqlp��x�hex���v�re?�Ɵx�key�v�pm��x�sus$�6�gcr���F������[�q27j9�2�v�ollis�mqSk�9O�ݝ� �(pl.���t��p!o��29$Fo8��cg�7no@�tptcls` CLS�o�b�F\�km�ai_
�s>�v�o	�t�b���ӿ�E�H��6�1e_nu501�[m���utia|$cal�maUR��CalMwateT;R51%�i=1]@-��/V� ���Z�� �fq1�9 "�K9E�L����2m�CLMTq�S#��3et �LM3!}t �F�c�nspQ�<c���c_moq��� ��c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 �̆�N�ve��C�cl�m�&Ao# �|$fi�nde�0S�TD ter FiLANG���R��
��n3���z0Cen���r, ������J����� � ��K��Ú�=���_�����r� "FNCDR�� 3��f��tguid�䙃N�."��J�tq�� ��� ����������J����_������c��	m��Z��\fndrA.��n#>
B2p��>Z�CP Ma������38A��� c��6� (���N�B���@���� 2�$�81�B�m_���"ex� z5�.Ӛ��c��0bSа�efQ���	��RBT;�OPTN �+#Q� *$�r*$��*$r*$%/ s#C�d/.,P�/0*ʲDPN��$����$*�Gr�$k E�xc�'IF�$MA�SK�%93 H5��%H558�$548 H�$4-1�$�d�#1(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9j0�"M�49�4  ���4�4tpsh���4�P�4- DQ�� �3�Q�4�R�4�pR@%0�2�r�4.b
E\���5�A�4��3adq}\�5K979":E��ajO l "DQ ^E^�3i�Dq ��4�ҲO ?R�? ��q@�5��T��3rAq�OF�Lst�5~��7p�5`��REJ#�2�@av^E�ͱ�F���4��.�5y� N� �2il(iqn�4��31 JH1��2Q4�251ݠ�4r'mal� �3)�RE o�Z_�æOx����4��8^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4$�REM���4yݱ"u<@�RER5932fO��47Z��5lity�,�U��e"Dil�\�5��o ��79�87�?�25 �3hk910�3��FE�0�=0P_�Hl\mhm �5��qe�=$�^��
E��u�IAympt�m�U��BU��vst e�y\�3��me�b�Dv I�[�Qu�:F�Ub�*_0�
E,�su��_	 Er��ox���4huse�E-�?�sn�������FE��,�Gbox�����c݌ ,"�������z���M��g��pdspw )�	��9���b���(��1���c�� Y�R�� �>�P���W�@�������'�0ɵ��[��͂��� � � ,K@�� �A�bu�mpšf��B*�BCox%��7Aǰ60�pBBw���MC� (6��,f�t I�s� ST��*��}B������w��"BBF�
�>�`���)��\�bbk968 "��4�ω�bb�9�va69����etb�Š��X�����ed�	�F��u�f� �s�ea"������'�\���,���b�ѽ�oH6�H�
�x�$�f����!y���Q[�! toperr�fd� �TPl0o� Rec�ov,��3D��R/642 � 0��C@�}s� N@��(U�rro���yu2r���  �
 � ����$$CL~e� ������������$z�_�DIGIT��������.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�o$j��+c:PR�ODUCTM�0\�PGSTKD��V�&ohozf99��D����$FEAT_INDEX���xd�� � 
�`ILEC�OMP ;����#��`�cSET�UP2 <�e��b�  N ��a�c_AP2BC�K 1=�i G �)wh0?{%&c����Q�xe% �I�m���8� �\�n����!���ȏ W��{��"���F�Տ j���w���/�ğS�� �������B�T��x� �����=�үa����� �,���P�߯t���� ��9�ο�o�ϓ�(� :�ɿ^���Ϗϸ� G���k� �ߡ�6��� Z�l��ϐ�ߴ���U� ��y����D���h� �ߌ��-���Q����� �����@�R���v�� ��)�����_����� *��N��r�� 7��m�&��3\�i
pP }2#p*.VRc�*��� /��PC/1/�FR6:/].��/+T�`�/�/F%��/�,�`r/?�*#.F�8?	H#&?�e<�/�?;STM� �2�?�.K �?�=�iPenda�nt Panel�?;H�?@O�7.O�?8y?�O:GIF�O�O��5�OoO�O_:JPG _J_�56_�O_�_��	PANEL1'.DT�_�0�_�_�?O�_2�_So�W Ao�_o�o�Z3qo�o@�W�o�o�o)�Z4�o�[�WI��
�TPEINS.XSML��0\����qCustom� Toolbar�	��PASSW�ORDyFR�S:\L�� %�Password Config�� �֏e�Ϗ�B0��� T�f����������O� �s������>�͟b� �[���'���K��� �����:�L�ۯp��� ��#�5�ʿY��}�� $ϳ�H�׿l�~�Ϣ� 1�����g��ϋ� ߯� ��V���z�	�s߰�?� ��c���
��.��R� d��߈���;�M��� q������<���`��� ����%���I������ ��8����n��� !��W�{" �F�j|�/ �Se��/�/ T/�x//�/�/=/�/ a/�/?�/,?�/P?�/ �/�??�?9?�?�?o? O�?(O:O�?^O�?�O �O#O�OGO�OkO}O_ �O6_�O/_l_�O�__ �_�_U_�_y_o o�_ Do�_ho�_	o�o-o�o Qo�o�o�o�o@R �ov��;�_ ���*��N��G� �����7�̏ޏm�� ��&�8�Ǐ\�돀�� !���E�ڟi�ӟ��� 4�ßX�j�������� įS��w������B��#��$FILE_�DGBCK 1=���/���� ( �)�
SUMMARY�.DGL���MD�:�����Di�ag Summa�ry��Ϊ
CONSLOG��������D�ӱConso?le logE�ͫ���MEMCHECCK:�!ϯ���X��Memory D�ata��ѧ�{�)��HADOW�ϣϵ�J���Sh�adow Cha�ngesM�'�-��)	FTP7�Ф�3ߨ���Z�mment TBD���ѧ0=4)ET?HERNET��������T�ӱEth�ernet \�f�iguratio�nU�ؠ��DCSV�RF�߽߫������%�� veri?fy all��'��1PY���DIF�F�����[���%=��diff]�������1R�9�K���c ���X��CHGD������cB��r����2Z8AS� ��GD���k��qz��FY3b8I[� �/"GD���s/�����/*&UPDATES.� �/��?FRS:\�/�-�ԱUpdate?s List�/���PSRBWLD.CM(?���"<?�/�Y�PS_ROBOWEL��̯�?�?� �?&�O-O�?QO�?uO OnO�O:O�O^O�O_ �O)_�OM___�O�__ �_�_H_�_l_o�_�_ 7o�_[o�_lo�o o�o Do�o�ozo�o3E �oi�o���R �v���A��e� w����*���я`��� ������O�ޏs�� ����8�͟\����� '���K�]�쟁���� 4���ۯj������5� įY��}������B� ׿�x�Ϝ�1���*� g�����Ϝ���P��� t�	�ߪ�?���c�u� ߙ�(߽�L߶��߂� ��(�M���q� �� ��6���Z������%� ��I���B�����2�����h����$FoILE_� PR� ���������MDO?NLY 1=.��? 
 ���q ����������~ %�I�m �2��h��!/ �./W/�{/
/�/�/ @/�/d/�/?�//?�/ S?e?�/�??�?<?�? �?r?O�?+O=O�?aO �?�O�O&O�OJO�O�O �O_�O9_�OF_o_
?VISBCKL6>[*.VDv_�_>.PFR:\�_�^�.PVisio�n VD file�_�O4oFo\_joT_ �oo�o�oSo�owo �oB�of�o� +������� +�P��t������9� Ώ]�򏁏��(���L� ^�������5���ܟ k� ���$�6�şZ���~�����
MR_�GRP 1>.�L��C4  B���	 W������*u����RHB ���2 ��� ��� ���B����� Z�l���C���D��������Ŀ��J8��L�J�ZG�F�5U��Ra�O���ֿ G�n�E��.E8�8�-���:uϚ{@ ����@�A�A��'f�?h!A���r���E�� F@� ������ھ��N�Jk�H9��Hu��F!��/IP�s�?�����(�9�<9���896C'�6<,6\b=��B�Y%���AD��=�@�eߋ�NҞ�A��߲�v��� r������
�C�.�@� y�d��������������?�Z�lϖ�B�H�� ��R�?��VE�������
�0�PJ��P�Hp1�ۿ���B���</ ��@�33:��q.�gN�UUU��U��q	>u.�?!rX��	��-=[z�=��̽=V6<��=�=�=�$q�����@8��i7G��8��D�8@9!�7�:�����D�@ D��g Cϥ��C������'/0-��P/� ���/N��/r��/���/ �??;?&?_?J?\? �?�?�?�?�?�?O�? O7O"O[OFOOjO�O �O�O�OPгߵ��O$_ �OH_3_l_W_�_{_�_ �_�_�_�_o�_2oo VohoSo�owo�o�i�� �o�o�o��);�o _J�j���� ���%��5�[�F� �j�����Ǐ���֏ �!��E�0�i�{�B/ ��f/�/�/�/���/� �/A�\�e�P���t��� �����ί��+�� O�:�s�^�p�����Ϳ ���ܿ� ��OH�� o�
ϓ�~ϷϢ����� �����5� �Y�D�}� hߍ߳ߞ��������o �1�C�U�y��߉� ������������-� �Q�<�u�`������� ��������;& _J\������� ���ڟ�F�j 4�������� �!//1/W/B/{/f/ �/�/�/�/�/�/�/? ?A?,?e?,φ?P�q? �?�?�?�?O�?+OO OO:OLO�OpO�O�O�O �O�O�O_'__K_� o_�_�_�_l��_0_�_ �_�_#o
oGo.okoVo ho�o�o�o�o�o�o �oC.gR�v �����	��� <�`�*<��`�� ���ޏ��)��M� 8�q�\�������˟�� �ڟ���7�"�[�F� X���|���|?֯�?�� ���3��W�B�{�f� ����ÿ�������� �A�,�e�P�uϛ�b_ �����Ϫ_��߀�=� (�a�s�Zߗ�~߻ߦ� ������� �9�$�]� H��l�������� ����#��G�Y� �B� ������z�������
 ԏ:�C.gRd� �����	� ?*cN�r�� ���/̯&/�M/ �q/\/�/�/�/�/�/ �/�/?�/7?"?4?m? X?�?|?�?�?�?�?�� O!O3O��WOiO�?�O xO�O�O�O�O�O_�O /__S_>_P_�_t_�_ �_�_�_�_�_o+oo Oo:oso^o�o�op��o �� ��$�� o�o�~���� ���5� �Y�D�}� h�������׏��� �
�C�.�/v�<��� 8������П���� ?�*�c�N���r����� ���̯��)��?9� _�q���JO�����ݿ ȿ��%�7��[�F� �jϣώ��ϲ����� ��!��E�0�i�T�y� �ߊ��߮��߮o�o� �o>�t�>��b �����������+�� O�:�L���p������� ������'K6 oZ�Z�|�~��� ��5 YDi �z������ /
//U/@/y/@��/ �/�/�/���/^/?? ?Q?8?u?\?�?�?�? �?�?�?�?OO;O&O 8OqO\O�O�O�O�O�O��O�O_�O7_��$�FNO ����VQ��
F0fQ kP oFLAG8�(LR�RM_CHKTY/P  WP��^P��WP�{QOM��P_MIN�P�����P�  X�NPSSB_CFG� ?VU ��_���S o�oIUTP_DEF�_OW  �|�R&hIRCOM�P�8o�$GENOV�RD_DO�V��6�flTHR�V dz�edkd_ENBWo� k`RAVC_?GRP 1@�WCa X"_�o_1 U<y�r�� ���	��-��=� c�J���n�������� ȏ����;�"�_�F��X���ibROU�`F\VX�P�&�|<b&�8�?���埘������� � D?�јs���@@g�B�7�p�)�ԙ\���`SMT�cG�m�M���� �LQHO7STC�R1H���P���at�SM���f�\����	127.0��1��  e��ٿ� ����ǿ@�R�d�v����0�*�	anonymous�����������/[�� � �����r����� �ߺ�����-���&� 8�[�I�π���� ��1�C��W�y� ��`�r������ߺ��� ����%�c�u�J\ n�������� �M�"4FX��i ������7/ /0/B/T/���m/ ��/�/�/??,? �/P?b?t?�?�/�?� �?�?�?OOe/w/�/ �/�?�O�/�O�O�O�O �O=?_$_6_H_kOY_ �?�_�_�_�_�_'O9O KO]O__Do�Ohozo�o �o�o�O�o�o�o
 ?o}_Rdv���_ �_oo!�Uo*�<� N�`�r��o������̏ ޏ�?Q&�8�J�\����>�ENT 1I��� P!􏪟  ����՟ğ�� �����A��M�(�v� ��^�����㯦��ʯ +�� �a�$���H��� l�Ϳ�����ƿ'�� K��o�2�hϥϔ��� ���ϰ�������F� k�.ߏ�R߳�v��ߚ� �߾���1���U��y��<�QUICC0 ��b�t����1�����%���2&���u��!ROUTER�v�R�d���!PC�JOG����!�192.168.�0.10��w�NA�ME !��!�ROBOTp�S_CFG 1H��� �A�uto-star�ted�tFTP�������  2D��hz� ���U��
//./A�#����~/ ����/�/�/�/�  ?2?D?V?h?�/?�? �?�?�?�?�?��� @O?dO�/�O�O�O�O �?�O�O__*_MON_ �Or_�_�_�_�_	OO -O�_A_&ouOJo\ono �o�o=o�o�o�o�oo �o4FXj|�_ �_�_o�7o�� 0�B�T�#x������� ���e�����,�>� ����ŏ���Ο ������:�L�^� p�����'���ʯܯ�  �O�a�s�����l��� ������ƿؿ�����  �2�D�g��zόϞ� �����#�5�G�I�� }�R�d�v߈ߚ�iϾ� �������)߫�<�N��`�r��XST_ERR J5
����PDUSIZ  ���^J����>~��WRD ?t���  guest}��%��7�I�[�m�$SCD�MNGRP 2K�t�������V$�K�� 	�P01.14 �8��   y�����B  �  ;����� ����������
 ������������~��`��C.gR|����  i  _�  
��������� +��������
���lZ .r���"�!l��� m
d�������_GROU���L�� �	����07EQUPOD  	պ�JV�TYa �����TTP_AUTH� 1M�� <!�iPendan�y��6�Y!KAREL:*��
-KC///A/� VISION SETT�/v/�"�/�/�/#�/�/ 
??Q?(?:?�?^?p>��CTRL Nв���5�
�?FFF9E3�?��FRS:DEF�AULT�<F�ANUC Web Server�:
�����<kO}O�O�O�O�O��WR_C�ONFIG OΡ� �?��ID�L_CPU_PC�@�B��7P�;BHUMIN(\��~<TGNR_IO�������PNPT_�SIM_DOmV�w[TPMODNT�OLmV �]_PR�TY�X7RTOLN/K 1P����_�o!o3oEoWoio�RMASTElP��R��O_CFG�o�iU�O��o�bCYCL�E�o�d@_ASG� 1Q����
  ko,>Pbt�� �������sk.�bNUM����K@�`IPCH�o��`RTRY_CN@xoR��bSCRN����Q��� �b�`�b�R���Տ��$�J23_DSP_�EN	����OBPROC�U�i�JOGP1SY@~��8�?�!��T�!�?*�POSR�E�zVKANJI�_�`��o_�� ��T��L�6͕����CL�_LGP<�_���EY�LOGGIN�`���LANG?UAGE YF7R�D w���LG���U�?⧈�xR� �����=P��'0��$ N�MC:\RSCH�\00\��LN_DISP V��`
��������OC�Rv.RDzVT=#�K@�9�BOOK W�
{��i��ii��X�����ǿٿ���b��"��6	h������e�?�G_B�UFF 1X�]��2	աϸ���� �������!�N�E� W߄�{ߍߺ߱����߀�����J���D�CS Zr� =����^�+�ZE���������a�IO 1[
{ ُ!� �!�1�C�U�i�y��� ������������	 -AQcu�������EfPTM  �d�2/AS ew������ �//+/=/O/a/s/p�/�/��SEV�����TYP��/??y͒�RS�@"��×�FL 1\
������?�?��?�?�?�?�?/?TP�6��">�NG�NAM�ե�U`�UPS��GI}�𑪅}mA_LOAD��G %�%D?F_MOTN���O��@MAXUALRM<��J��@sA�Q�����WS ��@C �]�m�-_���MP2�7�^�
{ ر�	�!P�+ʠ�;_/��Rcr�W�_�WU�W �_��R	o�_o?o"o coNoso�o�o�o�o�o �o�o�o;&Kq \�x����� ��#�I�4�m�P��� |���Ǐ���֏��!� �E�(�i�T�f����� ß��ӟ���� �A� ,�>�w�Z�������ѯ ����د���O�2� s�^�������Ϳ����ܿ�'��BD_LDXDISAX@	��MEMO_APR@�E ?�+
 � *�~ϐϢϴ�����������@ISC ;1_�+ ��I� �T��Q�c�Ϝ߇��� ������w����>�)� b�t�[����{��� �������:���I�[� /������������o� ����6!ZlS� �s���� 2�AS'�w� ���g��.//�R/d/�_MSTR� `�-w%SCD 1am͠L/�/H/ �/�/?�/2??/?h? S?�?w?�?�?�?�?�? 
O�?.OORO=OvOaO �O�O�O�O�O�O�O_ _<_'_L_r_]_�_�_ �_�_�_�_o�_�_8o #o\oGo�oko�o�o�o �o�o�o�o"F1 jUg����� ����B�-�f�Q����u�����ҏh/MK�CFG b�-�㏕"LTARM_���cL��� σQ�N�<�ME�TPUI�ǂ����)NDSP_CM�NTh���|�  d�.��ς�ҟ|ܔ|�POSCF�����PSTOL �1e'�4@�<#�
5�́5�E�S�1� S�U�g�������߯�� ӯ���	�K�-�?����c�u�����|�SIN�G_CHK  ���;�ODAQ,�f���Ç��DEV �	L�	MC:>!�HSIZEh��-���TASK �%6�%$1234?56789 �Ϡ���TRIG 1g.�+ l6�%����ǃ�����8�p�YP�[� ��EM_IN�F 1h3�� `)AT?&FV0E0"ߙ��)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ������H�����A���AI�q�,��|���� ���ߵ����� J���n������W��� ��������"����X ��/����e�� ����0�T;x �=�as��/ �,/c=/b/�/A/ �/�/�/�/��?� ��^?p?#/�?�/�? s?}/�?�?O�?6OHO �/lO?1?C?U?�Oy? �O�O3O _�?D_�OU_�z_a_�_�ONIT�OR��G ?5� �  	EXESC1Ƀ�R2�X3�XE4�X5�X���V7�X8�X9Ƀ�RhBLd �RLd�RLd�RLd
bLd bLd"bLd.bLd:bLdTFbLc2Sh2_h2khU2wh2�h2�h2�hU2�h2�h2�h3Sh�3_h3�R�R_G�RP_SV 1i�n���(ͅ�
��Å��ۯ_MO�x�_D=R^��PL�_NAME !�6��p�!De�fault Pe�rsonalit�y (from �FD) �RR2�eq 1j)TUX�)TX��q��X dϏ8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������2'�П�����*� <�N�`�r��<���� ����ү�����,��>�P�b� �Rdr 1�o�y �\�, Ӗ3���� @oD�  ��?���➱?䰺��A'��6����;�	l�ʲ	 �xoJ������ �<; �"�� �(p�K�K ���K=*�J���J���JV��0�Z�����rτ���p@j�@T;f���f��ұ]�^l��I��p������������b��3��´  �
`��>����bϸ�z���꜐r�Jm��
� B�H�˱`]Ӂt�q�	� p��  P�pQ��p��p|  ���g���c�	'� �� ��I� �  �����:�È
�È=G���"�s��	����I  �n @B�cΤ�\��ۤ�!�tq�y߁rN���  '�����@2��@����¬��/�C��C�C��@ C�������
�A���   @<�*P�R�
h�B�b�A��j�����������Dz۩��߹������j��( ?�� -��C�`��'�7�����q��Y����� �?�ff ��gy �����q�:a��
>+�  PƱj�(����7	����|�?���xZ�p<
6b�<߈;܍��<�ê<� �<�&Jσ�A�I�ɳ+���?ff�f?I�?&�k�@��.��J<?�`�q�.�˴ fɺ�/��5/���� j/U/�/y/�/�/�/�/��/?�/0?q��F �?l??�?/�?+)��?�?�E�� E��I�G+� F� �?)O�?9O_OJO�OXnO�Of�BL޳B� ?_h�.��O�O��%_�O L_�?m_�?�__�_�_x�_�_�
�h�Îg>��_Co�_`goRodo�o�GA�ds�q�C�o�o�o|����$]Hq�m��D��pC����pCHmZZ7t����6q�q��ܶN'�3�A�A�AR1�AO�^?�$��?�K�0±
�=ç>�����3�W
=�#��W��e�צ�@�����{�����<��(��B�u��=�B0�������	L��H�F��G���G���H�U`E����C�+���I#��I��HD��F��E���RC�j=��
�I��@H��!H�( E<YD0q�$�� H�3�l�W���{����� ���՟���2��V� A�z���w�����ԯ�� ������R�=�v� a������������߿ ��<�'�`�Kτ�o� �Ϻϥ��������&� �J�\�G߀�kߤߏ� �߳�������"��F� 1�j�U��y����� �������0��T�?��Q����(�1���3/E�����5�������q3�8������q4Mgs8&IB+2D��a���{� ^^	������JuP2P7Q4_�A��M0bt��R������/   �/�b/P/ �/t/�/ *a)_3/�/�/�%1a?�/?p;?M?_?q?  �?��/�?�?�?�?O 2� F�$�vGb	�/�A��@�a�`�qC��C@�o�O2��~�OF� DzH@��� F�P DC���O�O�ys<O�!_3_E_W_i_s?̯��@@pZ.tR22!2~
 p_�_�_�_	o o-o?oQocouo�o�op�o�o��Q ��+���1��$MS�KCFMAP  ��5� ��6�Q�Q"~�cON�REL  
�q3�bEXCFENB?w
s1uXq�FNC_QtJOG_OVLIM?wdIp�Mrd�bKEY?w��u�bRUN�|��u�bSFSPD�TY�avJu3sSI�GN?QtT1MO�T�Nq�b_CE_GRP 1p�5s\r���j��� ��T��⏙������ <��`��U���M��� ̟��🧟�&�ݟJ� �C���7�������گ��������4�V�`T�COM_CFG 1q}�Vp�����}
P�_ARC_\r�
jyUAP_C�PL��ntNOCH�ECK ?{ 	r��1� C�U�g�yϋϝϯ����������	��({NO_WAIT_L�l	uM�NTX�r{z�[m�_ERRY�s2sy3� &�������r�c� �^�T_MO��t��, �D$�k�3�_PARAM��u{��V[��!�u?��� =9@345678901��&� ��E�W�3�c�����{�0������ �����=�UM_RSPACE �Vv���$ODRDSP����jxOFFSE?T_CARTܿ��DIS��PEN_FILE� �q���c֮�OPTION�_IO��PWO_RK v_�ms �P(�R�Q
�8j.j	 ��Hj�&6$� RG_D?SBL  �5Js��\��RIEN�TTO>p9!C�ܧPq=#�UT�_SIM_D�
r�b� V� LCT ww�bc��U)>+$_PEXE�d&RATp �vju�p���2X�j)TUX)�TX�##X d-�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?O�H2�/oO�O�O�O�O�O �O�O�O_]�<^O;_ M___q_�_�_�_�_�_��_�_o���X�OU�[�o(��(����$o�, ��IpB` @D7�  Ua?�[cAa1?��]a]�DWcUa<쪋l;�	lmb�`��xJƯ`�����a��< ��`� ���b, H(��H�3k7HSM5G��22G���G�p
��
�!��X'|, CR�>��>q�GsuaT�37���  �4spBp�yr  ]o�*SB_�����j]��gt�q� ���rna �,���6�  ��PQ*�|N�M�,�k�!�	'� �� ��I� ��  ��%�=�C�ͭ���ba	����I  �n @��~���p��1��� �N U�[��'!o�:q�pC\�C��@@sBq�|��� �m�
�A\��h@�ߐ�n����Z�B�\��A���p� �-�qbz�P���t�_������(� �� -���恊�n�ڥ[A]Ѻ��b4�'!��(p �?�ff� ��
��B��OZ�R��8��tz���>΁  Pia��(�ವ@���ک�ax�c�dF#?�����x����<
6b<�߈;܍�<��ê<� <G�&�o&�)�A��lcΐI�*�?fff�?�?&c���@��.uJ<?�`��Yђ^�nd�� ]e��[g��Gǡd<�� ��1��U�@�y�dߝ� �ߚ����߼�	���-��������&��"�E��� E��G+� Fþ�������� ���&��J�5��bB��AT�8�ђ��0� 6���>���J�n�7���[m�0��h���1��>� M�I
�@��#A�[��C-�x)��?���P� /�YĒ��Jp��vav`CH/������}!@I��Y�'�3A�A��AR1AO�^?�$�?�����±
=ç>�����3�W
�=�#����+e���ܒ�����{����<��.�(�B�u�����=B0�������	�*H��F�G���G���H�U`E���C�+�-�I#�I���HD�F���E��RC�j=�U>
I��@�H�!H�( E<YD0/ �?�?�?�?�?O�?3O OWOBOTO�OxO�O�O �O�O�O�O_/__S_ >_w_b_�_�_�_�_�_ �_�_oo=o(oaoLo �o�o�o�o�o�o�o �o'$]H�l �������#� �G�2�k�V���z��� ŏ���ԏ���1�� U�g�R���v�����ӟ@�������-��(��g�������a����Q�c�,!�3�8�}���,!4�Mgs����ɢIB�+կ篴a���{���A�/�e�PS���w��P!�P�������7��ӯ�ϑ�R9�Kτ�o�X�ϓϥ�  ���� �����)��M����@������{߉ߛ����ߒߤ�������  )�G�q�_�����2 F�$N�&Gb���n�[XZjM!C�s�@j�/�A�S���F� �Dz��� F�P D��W����)�����������~x?���@@
�9�E�E��:E��
 v ��������*<N`�*P ����˨�1���$PARAM_M�ENU ?-���  �DEFPUL�SEl	WAI�TTMOUT��RCV� S�HELL_WRK�.$CUR_ST�YL�,OP9T�/PTB./("�C�R_DECSN���,y/�/�/�/ �/�/�/?	??-?V?�Q?c?u?�?�USE�_PROG %�%�?�?�3CCR������7_HO�ST !�!�44O�:T̰�?PCO�)ARC�O�;_TI�ME�XB�  ~�GDEBUGV@���3GINP_FOLMSK�O�IT`�\�O�EPGAP �L���#[CH�O�HTWYPE����? �?�_�_�_�_�_oo 'o9obo]ooo�o�o�o �o�o�o�o�o:5 GY�}���� �����1�Z��EWORD ?	7]�	RS`�	�PNS�$��J9OE!>�TEs@WV�TRACECTL� 1x-��� ��e ⹰Ӱ��ɆDT �Qy-���D� � ��ӱ4�P :�L �:�GP:�D :�@ :��8�8�	8�
8��8�8�8�8��8�X@:�8�8��8�8�8��:�"8�8�x�:�8�P�(:�d :�8�8��Ш:�
�:�!8�"8�#�8���:�%8�&8�'*8�(8�)8�*8����:�,8�-8�.8�/
8�08�18�,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� (�p������������� �� $6HZl ~�������  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_d��_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�_���*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p�������� //$)�$PG�TRACELEN�  #!  �_�" �8&�_UP z����g!o S!�h 8!_CFG �{g%Q#"!x!��$J �#|"DEFS_PD |�,!!�J �8 IN T_RL }�-" �8�%�!PE_CO�NFI� ~g%'�g!�$�%�$WLID�#�-74?GRP 1�7Q!��#!A ����&ff"!A+3�3D�� D]� CÀ A@+6
�!�" d�$�9�9*1~*0� 	 +9p�(�&�"�? ´	C�?�;B@3AO�?O�IO3OmO"!>�T?�
5�O�O�N�O� =��=#�
�O_�O_J_5_n_ Y_�O}_�_y_�_�_�_�  Dzco" 
 oBo�_Roxoco�o�o �o�o�o�o�o>�)bM��;
V�7.10beta�1�$  A��E�rӻ�Ay " �p?!G��q/>���r��0�q��ͻqBQ��qA\�p�q�4�q�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏��� 4��1�j�U���y��� ��֟������0�� T�?�x�c�������ү ����!o�,�ۯP�;� M���q�����ο��� ݿ�(��L�7�p�+9<��sF@ �ɣ� �ϥ�g%������+� !6I�[߆������ߵ� ����������!��E� 0�B�{�f������ �������A�,�e� P���t���������� ��=(aL^ ������� '9$]�Ϛ��ϖ �������/<�5/ `�r߄ߖߏ/>�/�/ �/�/�/?�/1??U? @?R?�?v?�?�?�?�? �?�?O-OOQO<OuO `O�O�O�O�O���O_ �O)__M_8_q_\_n_ �_�_�_�_�_�_o�_ 7oIot���o�o� ��o�o�o(/!L/^/ p/�/{*o���� �����A�,�e� P�b����������Ώ ��+�=�(�a�L��� p������Oߟ񟠟�  �9�$�]�H���l�~� ����ۯƯ���#�No `oro�on��o�o�o�o Կ���8J\n g����vϯϚ����� ��	���-��Q�<�u� `�r߫ߖ��ߺ����� ��;�M�8�q�\�� ������z������%� �I�4�m�X���|��� ��������:�L�^� ��Z��������� ��$�6�H�S wb������ �//=/(/a/L/�/ p/�/�/�/�/�/?�/ '??K?]?H?�?��? �?f?�?�?�?O�?5O  OYODO}OhO�O�O�O �O�O�O&8J4_F_ ����_�_��_�_ "4-o�O*ocoNo �oro�o�o�o�o�o �o)M8q\� �������� 7�"�[�m��?����R� Ǐ���֏�!��E� 0�i�T���x������� �_$_V_ �2�l_~_�_�����R�$PL�ID_KNOW_�M  �T������SV ���U͠�U��
��.�ǟ�R�=�O�����mӣM_GRP 1�પ!`0u��T@ٰo�ҵ�
���Pз j��`���!�J�_� W�i�{ύϟϱ����ϰ����߱�MR���b��T��s�w� s� �ߠ޴߯߅��ߩ߻� ����A���'��� ������������ =���#���������`}������S��ST���1 1��U# �v��0�_ A . ��,>Pb��� �����3( iL^p������2*���<-/3/)/;/M/4f/x/�/�/A5�/�/�/�/6??(?:?7S?e?w?�?8�?�?�?�?�MAD  d�#`PARNU/M  w�%O�SCH?J ME
��G`A�Iͣ�EUPD�`OrE
a�OT_C�MP_��B@�P@'�˥TER_CHK'U��˪?R$_�6[RSl�¯��_M�OA@�_�U_�_RE__RES_G � �>�oo8o+o\oOo �oso�o�o�o�o�o�o �o�W �\�_% �Ue Baf�S� � ���S0����S R0��#��S�0>�]��b��S�0}������RV� 1�����rB@c�]��t�(@c�\����D@c�[�$���RTHR_INRl�DA��˥�d,�MASS9� �ZM�MN8�k�MO�N_QUEUE ����˦��x� *RDNPUbQN{�P[���END���_ڙEcXE�ڕ�@BE�|ʟ��OPTIOǗ��[��PROGRAoM %��%���ۏ�O��TASK_�IAD0�OCFG ����tO��ŠDA�TA���Ϋ@��27�>�P�b�t��� ,�����ɿۿ������#�5�G���INFO
Uӌ�������ϭ� ����������+�=� O�a�s߅ߗߩ߻��ߠ�����^�jč� �yġ?PDIT ��ίc���WER�FL
��
RGA�DJ �n�AЄ���?����@���I�ORITY{�QV�>��MPDSPH������Uz����OT�OEy�1�R� _(!AF4�E�P�]���!tcp|h���!ud�>�!icm��ݏn6�XY_ȡ�R�{�ۡ)� *+/ ۠�W: F�j����� �%7[Bz�*��PORT#��BC۠����_CARTREP
�|R� SKSTAz�^�ZSSAV���n��	2500H8�63���r�$!�*R����q�n��}/�/�'� URGE��B��rYWF� DO{�rUVWV��$�A��WRUP_DE?LAY �R��$�R_HOTk��%�O]?�$R_NOR�MALk�L?�?p6S�EMI?�?�?3AQ�SKIP!�n�l#x 	1/+O+  OROdOvO9Hn��O�G �O�O�O�O�O_�O_ D_V_h_._�_z_�_�_ �_�_�_
o�_.o@oRo ovodo�o�o�o�o�o �o�o*<Lr�`���n��$R�CVTM������pDCR!�L�ЈqC`N�C����C�Q?���>r��<|��{4M�g�&���/��Z���t����l4��{�4Oi��O �<
6b<߈�;܍�>u.��?!<�& {�b�ˏݏ��8���� �,�>�P�b�t����� ����Ο���ݟ�� :�%�7�p�S������ ʯܯ� ��$�6�H� Z�l�~�������ƿ�� �տ���2�D�'�h� zϽ��ϰ��������� 
��.�@�R�d�Oψ� �߅߾ߩ������� ��<�N��r���� ����������&�8� #�\�G�����}����� ������S�4FX j|������ ���0T?x �u����'/ /,/>/P/b/t/�/�/ �/�/�/�/�?�/(? ?L?7?p?�?e?�?�? ��?�? OO$O6OHO ZOlO~O�O�O�?�?�O �O�O�O __D_V_9_ z_�_�?�_�_�_�_�_ 
oo.o@oRodovo�X��qGN_ATC �1�� �AT&FV0E0��kATDP/6/9/2/9�h�ATA�n,�AT%G1%B�960�i++U+�o,�aH,�q�IO_TYPE � �u�sn_�oR�EFPOS1 1}�P{ x�o�Xh_�d_��� ��K�6�o�
���.�ාR����{{2 1�P{���؏V�ԏxz����q3 1���$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����<�>��S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB��-�f��S8 1� ����Y�������y��SMASK 1��P  
9�G��XNOM���a~߈�~�qMOTE  h��~t��_CFG ᢥ����рrPL_�RANG�ћQ��POWER ��e���SM_DRYPRG %i��%��J��TART� �
�X�UME_PRO'�9��~t�_EXEC_EN�B  �e��GS�PD������c��T3DB���RM���MT_!�T����`OBOT_NA_ME i�����iOB_ORD_�NUM ?
��\qH863�  �T���������bPC_TIMoEOUT�� x�`oS232��1��k� LTEA�CH PENDA1N �ǅ�}����`Mainte�nance Co#ns�R}�m
"{�d?KCL/Cg��Z� ��n� ?No Use}�8	��*NPO��Ѯ����(C7H_L��������	�mMAVA#IL��{��ՙ��SPACE1 2��| d��(>��&���p��M,?8�?�ep/ eT/�/�/�/�/�W/ /,/>/�/b/�/v?�? Z?�/�?�9�e�a�=? ?,?>?�?b?�?vO�O�ZO�?�O�O�Os�2�/O*O<O�O`O �O�_�_u_�_�_�_�_[3_#_5_G_Y_o }_�_�o�o�o�o�o[4.o@oRodovo $�o�o����"�	�7�[5K]o� �A����	�̏�?�&�T�[6h�z��� ����^�ԏ���&�� ;�\�C�q�[7���� ����͟{���"�C�@�X�y�`���[8�� ��Ưدꯘ��0�?π`�#�uϖ�}ϫ�[Gw �i� ��:�
G� ���� $�6�H�Z�l�~ߐ��8  ǳ�����߈��d(���M�_�q�� ����������?� ��2�%�7�e�w����� ��������������� !�RE�W����� �����?�Q `�� @ 0��ߖrz	�V_�����
/ L/^/|/2/d/�/�/�/ �/�/�/?�/�/�/*? l?~?�?R?�?�?�?�?@�?�?�?2O�?
���O[_MODE � �˝IS �"��vO,*ϲ��O-_��	M_v_#dCWORK_AD�M�D�$bR  ���ϰ�P{_�P_I�NTVAL�@�����JR_OPTIO�N�V �EBpV�AT_GRP 2ݭ���(y_Ho �e_vo�o �oYo�o�o�o�o�o *<�bOoNDpw ������	�� �?�Q�c�u�����/� ��ϏᏣ����)�;� ��_�q���������O� ɟ���՟7�I�[� m�/�������ǯٯ� ���!�3���C�i�{� ��O���ÿտ���� ��/�A�S�e�'ωϛ� ��oρ�������+� =���a�s߅�Gߕ߻� ���ߡ���'�9�K� ]��߁����y��� �������5�G�Y��E��$SCAN_T�IM�AYuew�R� �(�#((��<0.a�aPaP
Tq >��Q��o������OO2�/���d;2BaR��WY��^��p�^R^	r  P���� � � 8�P�	�D��GYk} ��������Qp/@/R/x/)P;�o\T���Qpg-�t�_DiKT��[  � lv%��� ���/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OWW �#�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o lO~Od+No`oro�o�o �o�o�o�o�o& 8J\n����8��u�  0�"0g �/�-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q�����$o ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E��� ��Do��������ҿ� ����,�>�P�b�t� �ϘϪϼ���������w
�  58�J�\� n߀ߒߜկ������� ��	��-�?�Q�c�u�p����� �� -����� �2�D�V�@h�z�������������������& ���%	123�45678�" +	��/� ` r������� �(:L^p ������� / /$/6/H/Z/l/~/� �/�/�/�/�/�/? ? 2?D?V?h?�/�?�?�? �?�?�?�?
OO.O@O o?dOvO�O�O�O�O�O �O�O__*_YON_`_ r_�_�_�_�_�_�_�_ ooC_8oJo\ono�o �o�o�o�o�o�oo "4FXj|���������	���s3�E�W�{�C�z  Bp��  � ��2���z��$SCR_GRP� 1�(�U8(�\x^ �@  �	!�	 ׃�� �"�$� ��-��+���R�w����D!~�����#����O����M-10i�A 890990�5 Ŗ5 M61CA >4��Jׁ
� ���0�����#�1�	"�z���О���¯Ҭ � ��c���O�8�J� ������!�����\ֿ��B�y����������A��$�  !@��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ �϶�������%��I� 4�m��<�l߃ߕ��߹�B���\���� 1��U�@�R��v�� ����������;���*<=�
F���?�<d�<�>HE����s@�:��� B����ЗЙ���EL�_DEFAULT�  �����B�MIP�OWERFL  ��$1 WFD�O $��ER�VENT 1������"�pL!�DUM_EIP���8��j!AF�_INE �=�!'FT���9!��4 ��[�!RPC_MAIN\>�J�n'VISw=���o!TP�PU��	d�?/!
PM�ON_PROXY@/�e./�/"Y/��fz/�/!RDMO_SRV�/�	g�/�#?!R C?�h,?o?!
pM�/��i^?�?!RLSgYNC�?8�8�?>O!ROS�.L�4�?SO"wO�#DO VO�O�O�O�O�O_�O 1_�OU__._@_�_d_ v_�_�_�_�_o�_?o�ocoiICE_K�L ?%y (�%SVCPRG�1ho8��e���o�m3��o�o�`4 �`5�(-�`6PU�`7@x}�`���l9��{�d:?��a�o� �a�oE��a�om��a ���aB���aj叟a ���a�5��a�]� �a����a3����a[� ՟�a�����a��%��a ӏM��a��u��a#��� �aK�ů�as���a�� mob�`�o�`8�}�w� ������ɿ���ؿ� ��5�G�2�k�VϏ�z� �Ϟ����������1� �U�@�y�dߝ߯ߚ� �߾�������?�*� Q�u�`������� �����;�&�_�J� ��n������������sj_DEV ~y	�MC:�L!`OUT�",REC� 1�Z� d =  	 	�������

 �Z�{0H6 lZ�~���� �� //D/2/h/z/ \/�/�/�/�/�/�/�/ ?�/,?R?@?v?d?�? �?�?�?�?�?�?OO (ONO<OrOTOfO�O�O �O�O�O�O_&__J_ 8_Z_\_n_�_�_�_�_ �_�_�_"ooFo4oVo |o^o�o�o�o�o�o�o �o0TBxf ����(��� ,��P�>�`���h��� ������Ώ��(�:� �^�L���p������� ܟ���� �6�$�Z� H�~���r�����دƯ ����2��&�h�V� ��z�����Կ�ȿ
� ����.�d�RψϚ� |ϾϬ��������� <��`�N�pߖ߄ߺ� ����������8�&��\�J�l��jV 1-�w Pl�	�� � �F<��
TYPEV�FZN_CFG ;�x�d�7�GRP 1y�A�c ,B� �A� D;� B}���  B4�RB21H�ELL:�(
� X����%RSR����E0 iT�x���� ��/Sew��  ��%@w�����#�1����A��2#�d����HK7 1��� ��� m/h/z/�/�/�/�/�/ �/�/
??E?@?R?d?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he�s_ (_:_L_^_��_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}.xcopy �fr:\*.* �virt:\tm�pback�Q=>�inspiron?:1228 �R�_x�_�_	o  }/�Ua�_�_�P�_aoso�o�d3�Ts:ord�erfil.dat.l�]�o�o�o	`=*�Rmdb:+o�] �o\n�i�_2o�_ ���
�o�Ao��d�v����
xyz�rate 61 �+�=�O������|���x4064 �� ̏]�o�������+�=��O������)�2076��˟\�n����o �o./�ӯ���	� ��/�˯\�n����� ��4�O������� ��7�пa�sυϘ��� 3�N�������(�:� ��]�o߁ߔ���9�ʿ �������$ϵ�H�Y� k�}�Ϣϴ������� ��� ߻�D�U�g�y���}6���emp��`192.168�.4��46:38�92������}.��*.d������`r���1 +=O���� ��2� ��cu��4~ �:prgst��.dg���U���
/��conslog�� �e/w/�/)io�</N/�/��/?�2�err?all.ls�/��p�/f?x?�? }9�����=?S�?�?O}0  ��?�:�?bOtO�O����?9?R@8736  WO�O�O�O�O�I�O `_r_�_��;_M_�_ �_o'�T�_�_co uo�o�?�?5O�G�o�o �oO"O�o�H�obt`����3�=6 U8��
� }5 � ��g�y����o�o9 T���	���@ҏ�c�u������$SN�PX_ASG 1ߺ������� P 0 �'%R[1�]@1.1����?���%֟��&�	� �\�?�f���u����� ���ϯ��"��F�)� ;�|�_�������ֿ�� ˿���B�%�f�I� [Ϝ�Ϧ��ϵ����� ��,��6�b�E߆�i� {߼ߟ���������� �L�/�V��e��� ����������6�� +�l�O�v��������� ������2V9 K�o����� ��&R5vY k�����/� �<//F/r/U/�/y/ �/�/�/�/?�/&?	? ?\???f?�?u?�?�? �?�?�?�?"OOFO)O ;O|O_O�O�O�O�O�O �O_�O_B_%_f_I_ [_�__�_�_�_�_�_ �_,oo6oboEo�oio {o�o�o�o�o�o�o L/V�e�� ������6���+�l�O�v�������PARAM ������ �	���P����O�FT_KB_CF�G  ヱ���P�IN_SIM  ���C�U�g������RVQSTP_DSB,�򂣟�����SR �/��� & MULT�IROBOTTA�SK�����T�OP_ON_ER/R  ����PTN /��@�A	�RI�NG_PRM� ���VDT_GR�P 1�ˉ�  	������������ Я�����*�Q�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߣ� �߲����������� 0�B�i�f�x���� ���������/�,�>� P�b�t����������� ����(:L^ p�������  $6HZ�~ �������/  /G/D/V/h/z/�/�/ �/�/�/�/?
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8___\_���VPRG_COUNT��@���R'ENBU��UM�S���__UPD 1�>/�8  
s_� oo*oSoNo`oro�o �o�o�o�o�o�o+ &8Jsn��� ������"�K� F�X�j���������ۏ ֏���#��0�B�k� f�x���������ҟ�� ����C�>�P�b��� ������ӯί������UYSDEBU)G�P�P�)�d�YH�SP_PASS�U�B?Z�LOG [��U�S)�9#�0�  ��Q)�?
MC:\��6���_MPC���U�$��Qñ8� �Q趿SAV ���ج�ǲ&�ηSV�;�TEM_TIM�E 1��[ (�m��&����}YT1SVGUNS�P֕U'�U���AS�K_OPTIONДP�U�Q�Q��BC?CFG ��[u�� n�A�a�` a�gZo��߃ߕ��߹� ������:�%�^�p� [��������� � ����6�!�Z�E�~�i� ��������&����� ��&8��nY� }�?��ԫ � �(L:p^� ������/ / 6/$/F/l/Z/�/~/�/ �/�/�/�/�/�/2?8  F?X?v?�?�??�? �?�?�?�?O*O<O
O `ONO�OrO�O�O�O�O �O_�O&__J_8_n_ \_~_�_�_�_�_�_�_ o�_ o"o4ojoXo�o D?�o�o�o�o�oxo .TBx��j �������� ,�b�P���t�����Ώ ��ޏ��(��L�:� p�^�������ʟ��� �o��6�H�Z�؟~� l�������د���ʯ  ��D�2�h�V�x�z� ��¿���Կ
���.� �>�d�Rψ�vϬϚ� �Ͼ�������*��N� �f�xߖߨߺ�8��� ������8�J�\�*� ��n���������� ��"��F�4�j�X��� |������������� 0@BT�x� d�����> ,Ntb���� ��/�(//8/:/ L/�/p/�/�/�/�/�/ �/�/$??H?6?l?Z? �?~?�?�?�?�?�?O �&O8OVOhOzO�?�O �O�O�O�O�O
__�O @_._d_R_�_v_�_�_ �_�_�_o�_*ooNo <o^o�oro�o�o�o�o �o�o J8n $O�����X����4�"�X�B�v���$TBCSG_G�RP 2�B��  �v�� 
 ?�   ������׏�������@1��U�g�z���ƈ��d, ���?~v�	 HC��d��>����e�CL  B���Пܘ��w���\)���Y  A�ܟ$�B�g�B�Bl�i�X��ɼ���X��  DA	J���r�����C�����үܬ���D�@ v�=�W�j�}�H�Z����ſ���������v�	V3.0�0��	m61c�	*X�P�u�g�&p�>���v�(:��� ��p͟�  O����p�����z�JCFG �B���� �����������=��=�c�q�K�qߗ߂� �ߦ��������'�� $�]�H��l����� ��������#��G�2� k�V���z��������� �����p*<N ���l����� ��#5GY} h����v�b�� >�// /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?d?R?t?v?�? �?�?�?�?O�?*OO :O`ONO�OrO�O�O� �O�O�O_&__J_8_ n_\_�_�_�_�_�_�_ �_�_�_oFo4ojo|o �o�oZo�o�o�o�o�o �oB0fT�x �������,� �P�>�`�b�t����� Ώ�������&�L� �Od�v���2�����ȟ ʟܟ� �6�$�Z�l� ~���N�����دƯ� � �2��B�h�V��� z�����Կ¿���� .��R�@�v�dϚψ� ���Ͼ�������<� *�L�N�`ߖ߄ߺߨ� ���ߚ�������\� J��n������� ���"���2�X�F�|� j��������������� .TBxf� ������ >,bP�t�� ���/�(//8/ :/L/�/�ߚ/�/�/h/ �/�/�/$??H?6?l? Z?�?�?�?�?�?�?�? O�?ODOVOhO"O4O �O�O�O�O�O�O
_�O _@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<oro`o�o�o�o�o �o�o�o&�/>P �/������ ���4�F�X��(� ��|�����֏���� Ə0��@�B�T���x� ����ҟ������,� �P�>�t�b������� ��������:�(� ^�L�n�������2d �����̿�$�Z�H� ~�lϢϐ��������� �� ��0�2�D�zߌ� �߰�j���������� 
�,�.�@�v�d��� �����������<� *�`�N���r������� ������&J\ �t��B��� ���F4j| ��^����/��  2 6# �6&J/6"�$TB�JOP_GRP �2���?  ?�X,i#��p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�x�'�!�!>���
5�59>�0+1�33=�CL� �fff?+0?�ffB� J1�%Y?d7�.���/>��2�\)?0�5����;��hCY� ��  @� �!B� � A�P?�?�3EC�  D�!�,�0�*BOߦ?�3JB���
:���Bl�0��0�$�1�?O6!?Aə�AДC�1sD�G6�=q�E�6O0�p��B�Q�;�A�� �ٙ�@L3D	��@�@__�O�O>BÏ\JU�OHH�1ts}�A@33@?1� C�� �@�_�_&_8_>��D�UV_0��LP�Q30<{�zR� @�0�V�P!o3o �_<oRifoPo^o�o�o �oRo�o�o�o�oM (�ol�p~���p4�6&�q5	�V3.00�#m761c�$*(��$�1!6�A� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,IR�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^S@;Q��|8�E`rz@/&�8�6&�<��1�w�^$ES�TPARS  �*({ _#HR��AB_LE 1�p+Z�6#|�Q� � 1�|��|�|�5'=!|�	�|�
|�|�˕6!�|�|�|���RDI��z!ʟܟ� ��$���O������ ¯ԯ�����S��x# V���˿ݿ��� %�7�I�[�m�ϑϣ� �����������U-�� ��ĜP�9�K�]�o���-�?�Q�c�u���6�N�UM  �*z!� >  Ȑ�����_CFG ������!@b IMEBF_TT����x#��a�VER��b�w�a�R 1�p+
' (3�6"1 ��  6!����������  �9�$�:�H�Z�l�~� ���������������^$��_��@x�
�b MI_CHAN�m� x� kDBGLV;0o�x�a!n �ETHERAD �?�� �y��$"�\&n ROUmT��!p*!�*�SNMASK��x#�255.�h�fx^$OOL�OFS_DI���[ՠ	ORQCTRL �p+;/�� �/+/=/O/a/s/�/ �/�/�/�/��/�/�/�!?��PE_DET�AI��PON_�SVOFF�33P_MON �H��v�2-9STRTC_HK ����42VTCOMPA�Ta8�24:0FPR�OG %�%�MULTIROB�OTTO!O06�P�LAY��L:_IN�ST_MP GL�7YDUS���?�2L�CK�LPKQUIC�KMEt �O�2SC�RE�@�
tps��2�A�@�I���@_Y���9�	S�R_GRP 1Ҿ� ��� \�l_zZg_�_�_�_�_�_�^�^�oj�Q'O Do/ohoSe��oo�o �o�o�o�o�o! WE{i�������	1234�567��!���X��E1�V[
 �}�ipnl/a�g?en.htmno���������ȏ~�P�anel setup̌}�?��0�B�T�f� ��񏞟 ��ԟ���o���� @�R�d�v������#� Я�����*���ϯ ůr���������̿C� �g��&�8�J�\�n� ����϶��������� uϣϙ�F�X�j�|ߎ� �����;��������0�B��*NUALR�Mb@G ?�� [���������� �� ��%�C�I�z�m�������v�SEV � ����t�E?CFG Ձ=]�/BaA$   B�/D
 ��/C� Wi{�����@�� PRց;C �To\o�I�6?K0(%����0 �����//;/ &/L/q/\/�/�/�/lƇD �Q�/I_��@HIST 1׾�9  (�0� ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1 Ec0p?0�?�?�?/C�'=?O>71n?�?	OO-O�1y3�?O5edit[2?MULTIRf?O��O�O2O� FOP=962vO __$_6_�O�O�A36�O�_�_�_ �_IR�_�_�_oo+o =o�_aoso�o�o�o�o Jo�o�o'9I|��a81�ou��� ���o���)�;� M��q���������ˏ Z�l���%�7�I�[� ��������ǟٟh� ���!�3�E�W���� ������ïկ�v�� �/�A�S�e�Pb�� ����ѿ������+� =�O�a�s�ϗϩϻ� ������ߒ�'�9�K� ]�o߁�ߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y��� v�����������	 �?Qcu��( ����)� M_q���6� ��//%/�I/[/ m//�/�/�/D/�/�/ �/?!?3?�/W?i?{? �?�?�?�����?�?O O/OAOD?eOwO�O�O �O�ONO`O�O__+_ =_O_�Os_�_�_�_�_ �_\_�_oo'o9oKo �_�_�o�o�o�o�o�o jo�o#5GY�o�}������?���$UI_PAN�EDATA 1������  	�}��0�B�T�f�x��� ) �����4�ۏ���� #�5���Y�@�}���v� ����ן�������1���U�g�N������ �1��Ïȯگ� ���"�u�F���X�|� ������Ŀֿ=���� ��0�T�;�x�_Ϝ� �ϕ��Ϲ������,���M��j�o߁ߓ� �߷������`��#� 5�G�Y�k��ߏ��� �����������C� *�g�y�`��������� F�X�	-?Qc ����߫���� ~;"_F� �|�����/ �7/I/0/m/�����/ �/�/�/�/�/P/!?3? �W?i?{?�?�?�?? �?�?�?O�?/OOSO eOLO�OpO�O�O�O�O �O_z/�/J?O_a_s_ �_�_�_�O�_@?�_o o'o9oKo�_oo�oho �o�o�o�o�o�o�o# 
GY@}d�� &_8_����1�C� �g��_��������ӏ ���^���?�&�c� u�\�������ϟ��� ڟ�)��M����� ������˯ݯ0��� ��7�I�[�m������ ����ٿ�ҿ���3� E�,�i�Pύϟφ���0����Z�l�}���1� C�U�g�yߋ�)߰� #������� ��$�6� ��Z�A�~�e�w��� ��������2��V��h�O����v�p��$�UI_PANEL�INK 1�v��  ��  ��}12�34567890 ����	-?G� ��o�����a ��#5G�	�����p&���   R�����Z� �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?.O@O ROdOvO�O O�O�O�O �O�O_�O�O<_N_`_0r_�_�_�0,���_ ��_�_�_ o2ooVo hoKo�ooo�o�o�o�o �o�o��,>r} ��������� ���/�A�S�e�w� �������я���t v�z����=�O�a� s�������0S��ӟ� ��	��-���Q�c�u� ������:�ϯ��� �)���M�_�q����� ����H�ݿ���%� 7�ƿ[�m�ϑϣϵ� D��������!�3�E� �_i�{�
�߂����� �������/��S�e� H���~��R~'�'� a��:�L�^�p��� ������������  ��6HZl~�� �#�5��� 2 D��hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?�/ �?�?�?�?�?�?m?O O&O8OJO\O�?�O�O �O�O�O�O�O[�_�� 4_F_)_j_|___�_�_ �_�_�_�_o�_0oo Tofo��o��o��o �o�o,>1b t����K�� ��(�:����{O ������ʏ܏�uO� $�6�H�Z�l������� ��Ɵ؟����� �2� D�V�h�z�	�����¯ ԯ������.�@�R� d�v��������п� ��ϕ�*�<�N�`�r� ���O�Ϻ�Io������ ���8�J�-�n߀�c� �߇����߽����o 1�oX��o|���� ���������0�B� T�f������������ ��S�e�w�,>Pb t��'���� �:L^p� �#���� // $/�H/Z/l/~/�/�/ 1/�/�/�/�/? ?�/ D?V?h?z?�?�?�??? �?�?�?
OO.O��RO dO�߈OkO�O�O�O�O �O�O_�O<_N_1_r_ �_g_�_7OM�m��$UI_QUI�CKMEN  >��_Ao�bRESTORE� 1�?  �|��Rto�o�im�o�o�o�o �o:L^p� %������o� ���Z�l�~����� E�Ə؏���� �Ï D�V�h�z���7����� ��/���
��.�@�� d�v�������O�Я� ����ßͯ7�I��� m�������̿޿��� �&�8�J��nπϒ� �϶�a�������Y�"� 4�F�X�j�ߎߠ߲� �����ߋ���0�B�T�gSCRE`?�#mu1s]co`u2��3��U4��5��6��7��y8��bUSERq�dv��Tp���ks����4��5��6��7���8��`NDO_�CFG �#k � n` `PDA�TE ����NonebSE�UFRAME  ��TA�n�RTO?L_ABRTy�l�Α�ENB����GR�P 1�ci/aCz  A�����Q@�� $6HR�d��`U�����MSK  �����MNv�%�U�%����bVISCAN�D_MAX�I���FAIL_�IMG� �PݗP#���IMREGN�UM�
,[SI�Z�n`�A�,~VONTMOU��@���2���a��a��~��FR:\� � MC{:\�\LOG�7B@F� !�'/�!+/O/�Uz �MCV�8#U�D1r&EX{+�S|�PPO64_���0'fn6PO��LIb�*�#9V���,f@�'�/�� =	�(SZV��.����'WAI��/STAT 	����P@/�?�?�:�$�?�?��2DW�P  ��P yG@+b=��� H��O_JMPE�RR 1�#k
 � �2345678901dF�ψO{O �O�O�O�O�O_�O*_�_N_A_S_�_
� M�LOWc>
 �_�TI�=�'M�PHASE  ���F��PSHI[FT�1 9�]@<�\�Do�U#oIo �oYoko�o�o�o�o�o �o�o6lCU �y����� �@�	�V�-�e2����	VSFT1�2�	VM�� ��5�1G� ���%A_�  B8̀̀E�@ pكӁ˂�у���z�ME@�?��{��!c>&%�aM�1��k�0�{ �$�`0TDINEND��\�O� �z���S��w��P��=�ϜRELE�Q���Y���\�_ACT�IV��:�R�A ���e���e�:�R�D� ���YBOX� �9�د�6���02���1�90.0.�83v��254�:�QF�	 �X��j��1�ro�bot���  � p�૿�5pc��̿������7�����-�f�ZABC�����,]@U��2 ʿ�eϢωϛϭϿ� ���� ���V�=�zߐa�s߰�E�Z��1� Ѧ