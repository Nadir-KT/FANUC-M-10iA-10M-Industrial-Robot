��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  �(��ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1����|UREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|�R�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"�SBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5� UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8�W�+0�$Y $DB\� 6COMW!2�MO� H.	 �\rVE�1$F8�RA{$O�UD�cB]CTMP1_FtE2}G1_�3�B�2��XD�#
� d $CARD_EXIST4�$FSSB_T�YP!AHKBD�_SNB�1AGN G�n $SLO�T_NUM�AP�REV4DEBU�� g1� ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�U0LEToE_OK�BUS�oP_CR�A$;4xAV� 0LACIw�1�R�@k �1$@M{EN�@$D�V��Q`PvVA{QLv� OU&R ,AЧ0�!� B� LM�_O�
eR�"CAsM_;1 xr~$ATTR4��@� ANNN@5I�MG_HEIGH|�AXcWIDTH4�VT� �UU0F_�ASPEC�A$�M�0EXP�.@A�X�f�CF�D ?X $GR� � �S�!.@B�PNFL�I�`�d� UIREx 3T!GITCH+Cj�`N� S�d_LZ`2AC�"�`EDp�dL� J�4S�0� <z�a�!p;G0 �� 
$WARNM�0f�!�@� -s�p�NST� CORN��"a1FLTR{uT�RAT� T}p ? $ACCa1�pp��|{�rORI�Pl�C�kRT0_S~B�\qHG,I1 E[ T�`�"3I�pCTYD�@*2 3`�#@� �!�B*HD�DcJ* Cd�2_�3�_�4_�5_�6_�7�_�8_�94�ACO�$ <� �o�o�h8K3 1#`O_Mc@AC_ t � E#f6NGPvABA�  �c1�Q8��`,��@n!r1�� d�P�0e�,��axnpUP&P�b26���p�"J�p_)R�rPBC��J�rĘߜJV�@U� B��s}��g1�"YtP_*0O�FS&R @� RcO_K8T��aIT�3�T�NOM_�0�1�p�34 >��D Ԑ� Ќ@��hPV��mE!X�p� �0g0ۤ�p��r
$TF�2C$7MD3i�TO�3�0yU� F� ��)Hw2tC1(�Ez�g0#E{"F�"F�40�CP@�a2 �@�$�PPU�3Nc)ύRևAX�!�DU��AI�3B�UF�F=�@1 �|pp���pPITV� PP�M�M��y��F�SIMQ�SI�"ܢVAڤT��=�w T�`(zM��P�B�qFACTb�@EW�P1��BTv?�MC�5 �$*1JB`p�*1DEC��F��ŏ��� �H0CH�NS_EMP1�#$G��8��@_4�3d�p|@P��3�TCc� (r/�0-sx��ܐ� `MBi��!����JR� �i�SEGFR��ITv �aR�TpN�C���PVF�?�bx &��f{uJc !�Ja��� !28�ץ�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb���q@�۽�н����L�83�B���CRC�e�3CCp����c��m cҞb�1J�cѿ�.���*�D$ICb�Cq�5r��ե��@v�'���EVT���zF��_��F,p)N��ܫ�?�4�0A�! �r���h �Ϩ��p�2�͕a��� �د�R�Dx Ϗ��o"27��!ARV�O`C�$L	G�pV�B�1�P��@��t�aA�0'�|�+0Ro�� MEp`"1 �CRA 3 AZ�V�g6p�O �FCCb�`�`F�`K������ADI��a�A �bA'�.p��p�`�c¢`S4PƑ�a�AMP���-`Y�3P�M���CUR��QUA1 � $@TITO1�/S@S�!����"0�D�BPXWO��B0!5�$SK���2ѓDBq�!"�"�PR�� 
� =���΁!# S q1$�2�$z���L�)$��/���� %�/�$Cr�!&?�$ENE�q�.'*?PA�!R�E�p2(H z��O�0#$L|3$$�#�B[�;���F�O_D��RO�Sr�#������3R�IGGER�6PA�pS����ETURN��2�cMR_8�TUrw��0EWM�ҍM�GN�P���BL�AH�<E���P��'&$P� �'P@�Q"3�CkD{��DQ���4�11��FGO_A7WAY�BMO�ѱQ�#!�DCS_޾)  �PIS � I gb {s�C��A��[ �B$�S��A�bP�@�EW-�TNT	Vճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_�SV�bEXCLUt��nONL2�b�SY�*a&�OT�a'�HI_V�4��B<���_ *P0� r9�_z��p �"v�@SG�� +nr r�@6Acc*b��G�#@�E�V.iHb?fANNcUN$0.$fdID�	U�2�SC@�`�i�a���j�f�(�@�pO�GI$2,O�$F�ibW$}�OT9@�1� $DUMMY T��da��dn�� � ��E- ` ͑HE4(sg�*b�SAB���SUFFIW�V�@CA=�c5�g�6r�!MSW�E.{ 8Q�KEYI5���TM�10s�qA�v�IN����D��/{ D��HOST_P!�rT��ta��tn��tsp�pEMӰV������pLc ULI�0  8	=ȳ��� Tk0�!1 � �$S��ESAMPL��j�۰f璱f����I�0��[ $SUB�k�#0�C��T�r#a�SAVʅ��c��`�C��P�fP$n0yE�w YN_B#72 0Q�DI{dlp�O(��9#$�R�_I�� �EN�C2_S� 3 ! 5�C߰�f�-  �SpU����!4�"g��޲�1T���5@X�j`ȷg��0�0K�4x�AaŔAVER�q8ĕ9g�DSP�v��PC��r"��(����ƓVALUߗHE4�ԕM+�IPճ���OPP ��TH��֤��P�S� �۰	F��df�J� �u�C1+6 H�bLL_DUs�~a3@{�0�3:���OTX"����s� ��0NO�AUTO�!7�p!$)�$�*��c4�(��C� 8�C, �"��!&�L�� 8H *8�LH <6� ���c"�`, `Ĭ�k� ��q��q��sq��~q���7��8��9��0T����1��1̺1ٺU1�1�1 �1ʕ1�2(�2����2�̺2ٺ2�2�2� �2�2�3(�3R��3��̺3ٺ3�U3�3 �3�3ʅ4(®�`��?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?g �@P?9��5�9�E�@A�!��A� ;p$T�P�$VARI�:�Z���UP2�P< ���TDe����K`Q�����BAC�"= T�p��e$�)_,�bn�kp+ IF�IG�kp�H  ��Pİ�"F@`�!>Gt ;E��sC�ST�D� D���c�<� 	C��{�� _���l���R  ���FORCEUP?b^��FLUS�`H��N>�F ���RD_CM�@E������ ��@vMP��REMr F �Q��1k@���7Q
�K4	NJ�5EFF�ۓ:�@IN2Q��O�VO�OVA�	TgROV���DTՀ�DTMX� � �@�
ے_PH"p��CL��_TpE�@d�pK	_(�Y_T��Tv(��@A;QD� ������!0tܑ&0RQ���_�a��2��M�7�CL�dρ�RIV'�{��EAmRۑIOHPC�@d����B�B��CM9@����R �GCLF�e!DYk(M�a6p#5TuDG��t� �%��`FSSD �s? P�a�!�1��E�P_�!�(�!1���E�3�!3�+5�&��GRA��7�@��4;�PW��ONn��EBUG_SD2H�P|{�_E A`��A��TERM�`5Bi5���O�RI#e0C�9SM�_�P��e0Di5=���TA�9Ei5�p�U}P\�F� -�A�{�AdPw3S@B$gSEG�:� EL{UwUSE�@NFIJ�B$�;1젎4�4C�$UFlP=�$,�|QR@��_G90qTk�D�~SNST��PAT����APTHJ3Q�E�p%B�`�'EC���@Rx$P�I�aSHFTy��A�A�H_SHOR(Р꣦6 �0$�7P9E��E�OVR=��aRPI�@�U�b �Q�AYLOW���I�E"��A��?���ERV��XQ�Y��mG>@@�BN��U\��R2!=P.uASYMH�.uFAWJ0G�ѡEq��A�Y�R�Ud>@��EC���EP;�uP;��6WOR>@M`� �0SMT6�G3�G1R��13�aPAL@����p�q�uH � :���TOCA�`yP	P�`$OP����p�ѡ�`0O,��RE�`R4C�A�O�p낎Be�`R��Eu�h�A��e$P�WR�IMu�RR�_�cN��q=B I�&2H���p_ADD�R��H_LENG��B�q�q�q$�R��S��JڢSS��SK�N��u\��u̳�uٳS�E�A�jrS��MN�!K�����b����OLX��p�<���`ACRO3pJ� �@��X�+��Q��6�OUP3�b_�IX��a�a1��}򚃳� ��(��H��D��ٰ���氋�IO2S��D�����	�7��L $l��`Y!_O�FFr��PRM_������HTTPu_+�H:�M (|p�OBJ]"�p��$���LE~Cd���N� � ��֑AB%_�TqᶔS�`6H�LVh�KR"u�HITCOU��B-G�LO�q����h�����`��`SS� ���HW�#A:��Oڠ<`INCP}U2VISIOW� ͑��n��to��to�ٲ�H�IOLN��P� 8��R��r�$�SLob PUTM_n�$p��P& �¢ ��Y F_AS:�"Q��$L�������Q  U�0	P4A0��^���ZPHY��-���x��UOI �#R `�K����$�u�"pPpk����$�����Y�UJ5�S�-���NE6WJOG�KG̲DIS���K�p���#T (�uAV8F�+`�CTR�C
��FLAG2�LG�dU ���؜�13?LG_SIZ����`b�4�a��a�FDl�I`�w� m�_�{0a� ^��cg���4�����������{0��� SCH�_���a7�N�d�V
W���E�"����4�"�UM�Aљ`LJ�@�7DAUf�EAU�p�X�d|�r�GH�b6��OGBOO��WgL ?�6 IT㸰�y0�REC��S#CR ܓ�D
�\���MARGm�!��@զ ��d%�����S�����W���U� �JG=M[�MNCHJ���_FNKEY\�K��7PRG��UF��7Pn��FWD��HL��STP��V��=@��,�А�RS��HO`����C9T��b ��7�[�UL���6�(RD� �d���Gt��@PO���������MD�FOC�U��RGEX��TKUI��I��4� @�L�����P� ���`��P��NE��C�ANA��Bj�VA�ILI�CL !�UDCS_HII4��s"�O�(!�S����S�瞴 ��BWUFF�!X�?PTH$m���v`��ěԃ�AtrY��?P��j�3��`OS1
Z2Z3ZD��� >� Z � ��[apEȤ��ȤIDX�d	PSRrO���zA�+STL�R}�Y&��� Y$E�C ���K�&&8�п![ LQ��+00�	P����`#qdt
�U�dt�$;��_ \ ��`4Г�\��Ѩ#w�MC4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#�1D���'B�LD�%�$�%ORGڰ5�2�P@VŇVY8�s�T�r �#}d^ ���$6��$
�%S�`T� �B0�4}�6RCLMC�4`]?o?�9세�MI�p�}d_ d=њRQz��DSTB�pƽ ;F�HHAX��R JHdLEXC#ESrD�BM!p�a`4�/B�T8B�j�`a�p=F_A7J�i��KbOtH�0K�db� \Q���v$MB�C�LI|�)SREQUIR�R�a.\o�AXODEBUZ�ALt M��c�b�{P����2ANDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��X�� N&��aZ�� ܺ �QPST� �ezrLOC�RI,rp�EX<fA�p��9AAODAQ��f� XY�OND��"MF,Łf�s"��}%��e/� �8FX3@I�GG�� g ���t"��ܓs#N�s$R�a%��iL��hL�xv�@�DATA#�?pE�%�tR��Y�N�h t $MD`qI}�)nv� ytq�ytHP`�Pxu��(�zsANSW)�yt@��yuD+�)\b���0no�i �@CUw�qV�p 0XeRR2���j Du�{Q��7Bd�$CALIA@��Gt��2��RIN���"�< �INT	E��Ck�r^�آXb,]���_N�qlk����9�D���Bm��DI�VFDH�@���qn�I$V,��S�$��$Z�X�o�*����oH �$BELTʾu!ACCEL�8.�~�=�IRC�� �䰠D�T�8�$P)S�@�"L���r���#^�S�Eы T�PACTH3���I���3x�p�A_W��ڐ���2rnC��4�_MG�$DD��T���$FW�Rp9��I��4��DE7�PPA�BN��ROTSPCEE�[g�� J���[�C@4���$U'SE_+�VPi�ƣSYY���1 �aY�N!@A�ǦOFFܐqǡMOU��NG����OL����INC�tMa6��HB��0HBENCS+�8q9B�p�4�FDm�IN�I`Ԓ]��B��VE��|#�y�23_UP�^��LOWL����p� B���Du�9B#P�`�x ���BCv�r�MgOSI��BMOU���@�7PERCH  ȳOV��â
ǝ ����D�ScF�@MP����� Vݡ�@y��j�LUk��Gj�p�U�P=ó���ĶTRK|��AYLOA�Q e��A��Ԓ����N`��F�RTI�A$��MOUІ�HB�BS0�p7D�5���ë�Z�D�UM2ԓS_BC?KLSH_CԒk� ���ϣ���=���xޡ �	ACLAL"�q��1м@��CHKt� �S�RTY�� ^�%E1Qq_�޴'_UM�@�C#���SCL0�r�LMT�_J1_L��9@H�qU�EO�p�b�_�8e�k�e�SPC�㡘u���N�PC�N�H�z \P��C�0~"X�T��CN_:�N�9��I�SF!�?�V ���U�/���ԒT���CB!�SH�:�� E�E1T�T����y����T��PA ��_P��_� =������!(����J6 L�@��晰OG�G�TORQU��ONֹ��E�`R��H�E�g_W2���_郅���UI�I�I��Ff`�xJ�1�~1�VC"3�0BD:B�1�@8SBJRKF�9�0DBL_SMt��2M�P_DL��2GRV����fH_��d����COS���LN H������� �!*,�aZ����fMY�_(�TH|��)THET0��NK23���"��[CB�&CB�CAA��B�"��!��!�&SqB� 2�%GTS�Ar�CIMa�����,4x#97#$DU�� �H\1� �:Bk62�:A9Q(rSf$NE�D�`AI��B+5��$̀�!A�%�5�7����LPH�E�2���2S C%C%�2-&FC(0JM&̀V�8V�8߀�LVJV!KV/KV�=KVKKVYKVgIH��8FRM��#X!KH�/KH=KHKKHYKH*gIO�<O�8O�YNUOJO!KO/KO=KUOKKOYKOM&F�2��!+i%0d�7SPBALANCE_o!�[cLE0H_�%S�Pc� &�b&�b&PFULC�h�b�g�b�%p�1k%�UTOy_��T1T2�i/�2N��"�{�t#�@Ѱ`�0�*�.�T���OÀ<�v INSE9G"�ͱREV4vͰ�l�DIF�ŕ�1llzw��1m�0OBpq�я?�MI{���n?LCHWARY����AB��!�$ME�CH�!o ��q�AX��P����7Ђ�`�n 
�d(�U�ROB��CRr�H�����(�MSK_|f`�p P �`_��R/�k�z�����1S�~�|�z�{���z���qINUq�MT�COM_C� �q�  ���pO��$NOREn�����pЂr 8p G�Re�uSD�0AB��$XYZ_D�A�1a���DEBU�Uq������s z`$COD�� �L���p�$B�UFINDX|��  <�MORm�t $فUA��֐�H��y��rG���u � $SIMUL  S�*�Y�̑�a�OBJE�`̖A�DJUS�ݐAY_IS�D�3���n�_FI�=��Tu 7�~�6�'��p} �=�C�}p�@b�D��F�RIr��T��RO�@ \�E}'���OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1�0e��M��ED}�*�p ��N�PMֲ���rc�w�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B�P2�G�B�_�M����q�E� x Hxw��p��ATUSWЅ��C�0o�s���BSTM�ǌ�I�k��4��x�԰q�y DBw�E&���@E�r���7��жЗ�EXE ��ἱ�����f q�gz @w���UP'�f�$�pQ�XN����������� �P�G΅{ h $GSUB����0_��|�!�MPWAIv�P7ã�LOR�٠F�\p˕$RCVF�AIL_C��٠B�WD΁�v�DEF�SP!p | L�w���Я�\���UCNI+�����H�R�,p}_L\pP��t�	P��p�}H�> �*��j�(�s`~�N�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��G���PLI��p� � $ˀP_S�WI�pq�J_PL~��AL_ ���J��A��B��� C���D�$E���.�C_�U�� � � ���*��J3K0����TIA�4��5��6��MOM��������ˀB��AD��������6��PU� NR�������G��m��?� A$PI�6q� �	�����K4��)6�U��w`��SPEEDgPG���� ����Ի�4T�� �� @��SAM�r`��\�]��MOV_�_$�npt5��5$���1���2���� ����'�S�Hp�IN�'�@�+�����4($4+T+GA�MMWf�1'�$G#ET`�p���Da���=

pLIBR>�I]I2�$HI=�_g�Ht��2�&E;��(A�.� �&LW�-6<�)@56�&]��v�p��V���$PDCK����q��_?���� �q�&���7��4����9+� �$I/M_SR�pD�s�r�F��r�rLE���O0m0H]��0�-�p�q��PJqUR_�SCRN�FA���S_SAVE_D��,dE@�NOa�CAA� b�d@�$q�Z�Iǡs	 �I� �J�K� ����H �L��>�"hq�� ����ɢ�� bWP^US�A�p��M4���a��)q`��3�W@W�I@v�_�=���MUA�o�� � $P9Y+�$W�P�vNG�{��P:��RA�0�RH��RO�PL������q� ��s'�X;�O�I�&�Zxe ���m��# p��ˀ�3s�O@�O�O�O�O�aa�_т� |��q�d@��.v ��.v��d@��[wFv���E���%w�.r;B��w�|�tP���P�MA�QUa ���Q8��1٠QTH��HOLG�QHY�S��ES��qUE��pZB��Oτ�  ـPܐ(�A����v�J!�t�O`�q��u��"���FA��IROG�����Q2���o�"�x�p��INFOҁ��׃V����R�H�O�I��� (�0SLEQ������Y�3�H���Á��P0Ow0Ԟ��!E0NU���AUT�A�COPY�=�/�'��@Mg�N��=�}1������� ��RG��Á�f��X_�P�$;�(���`��W��P��@������EXT_CYC bHᝡRprÁ�r��_NAec!А���ROv`~	�� � ���POR_�1�E2��SRV �)_�I�DI��T_�k�}�'����dЇ�����5��6J��7��8i�H�SdBZ���2�$��F�p���GPLeAdA
�TAR�Б@���Pp�2�裔d� ,�0cFL`�o@YN���K�M��Ck��PW�R+�9ᘐ��DE�LA}�dY�pAD��a"�QSKIPN4� �A�$�OB`�NT����P_ $�M�ƷF@\bIpݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q����TQ������ ���`�#�RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�d"�REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"�������2�Қ�߼���P������3�қ'�@9�K�]�o���4���������������5�ҝ!�3�E�W�i�{��6�Ҟ������P�������7�ҟ@-?Qcu�8����������SMSKÁ�l��a��EkA��MOT-E6�����@��݂TQ�IO}5�I�S�tR�W@���� �pJ���n Ȝ�����E�"$DSB_SIGN�1�UQ�x�C\��S2�32���R�iDE?VICEUS�XR>SRPARIT��4!_OPBIT�QI�OWCONTR+��TQ��?SRCU� M~pSUXTASK�3�N�p�0p$TATUF�PE#�0������p_XPC)�$F�REEFROMS8	pna�GET�0���UPD�A�2��S�P� :��� !>$USAN�na8&����ERI�0_�&RpRYq5*"_j@_�qPm1�!�6WRK9�KD���6��QFR�IEND�Q�RUFxg�҃�0TOOL�6�MY�t$LEN�GTH_VT\�FCIR�pC�@ˀE> �+IUFIN-RM�ΕRGI�1ÐAITI�$GXñ3IvFG2v7G1���p3��B�GPR�p�1F�Oa_n 0��!RE��0p�53҅U�TC��3A�A�F �G(��":���e1n!��J�8 �%���%]��%�� 74��X O0�L
��T�3H&��8���%�b453GE�W�0�WsR�TD����T��M�����Q�T]�$V �2����1�а91T�8�02�;2k3�;3�:ifa�9-i�aQ0��NS��ZR$V��2B%VwEV�2ALQ�B
;�����&�S�`���F�"�k�@�2a�PS�E��$r1C���_$Aܠ6wPR��7vMU�cS�t '�/89�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx_�����BSOC����N��DUMMY�14�p�0SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU""ƐS�P �M�)0NS��cM�"r�$HW_C��U��S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}��#!�_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�S�AC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EG� �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G + AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC  o�ER|f�5� � $�@�_ A��!�PO���à�0#�
�_M�RAt�� d r� T��ٔERR��L��;TY&���I��qV�0�cz�TOQ�d�PL[ �d�"�� ?�|w�! � pp`qT)0���_V1VrP�aӔ����2ٛ2薈E����@�H�E����$W�����V!��$�P��o�cI���aΣ	 HELL�_CFG!�� 5��B_BAS�q�SR3��� Ea#Sb���1�U%��2��3��4��U5��6��7��8����RO����I0�0NL�\CAB+�����ACK4�����,��p2@�&�?�_PUﳳCO. U�OUG�P�~ ����m�������T=Pհ_KAR�l�&_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h��]�l0SEM�4�(��M4�6�TYN�SO���DIZ�~�A������m_TM�MA'NRQ��k0E�����$KEYSWI�TCH���m���H=E��BEAT���E- LE~�����U±�F!Ĳ���B�O_�HOM=OGREFUPPR&��y!� �[�C��O��-EC�OC��Ԯ0_IOC�MWD
�a�B(8k��� � Dh1���UX���M�βgPgCFORC������OM.  � @��5(�U�#P, 1���, 3��45~	�NPX_ASt�w� 0��ADD�о�$SIZ���$VAR���TI�P/�.��A�ҹ�M�ǐ��/�1�+ U"S��U!Cz���FRI	F��J�S���5Ԓ��NF�Ѝ� � mxp`SI��TE�C\���CSGL��TQ2��@&����� ��S'TMT��,�P �&�BWuP��SHOW�4���SV�$��� �Q�A00 �@Ma}���� ��ਅ�&���5��6��7*��8��9��A��O ����Ѕ�Ӂ���0��F ��� G��0G���0 G���@G��PG��U1	1	1	1+	U18	1E	2��2��U2��2��2��2��U2��2��2��2��U2	2	2	2+	U28	2E	3��3��U3��3��3��3��U3��3��3��3��U3	3	3	3+	U38	3E	4�4��U4��4��4��4��U4��4��4��4��U4	4	4	4+	U48	4E	5�5��U5��5��5��5��U5��5��5��5��U5	5	5	5+	U58	5E	6�6��U6��6��6��6��U6��6��6��6��U6	6	6	6+	U68	6E	7�7��U7��7��7��7��U7��7��7��7��U7	7	7	7+	e78	7E��VP���UPDs�  ��`NЦ�5�YSL}Ot�� � L�`��d���A�aTA�80d��|�ALU:ed��~�CUѰjgF!aIgD_L�ÑeHI�j�I��$FILE_����d��$2�fS�A>�� hO��`E_BLCK��b$�>�hD_CPUyM�@yA��c�o�d��Y��ޅ�R �Đ
P�W��!� oqLA®�S=�ts�q~tRUN�qst�q~t���p�qst�q~t �T���ACCs��Xw -$�qLEN;� �tH��ph�_�I��ǀLOW_AXI�SF1�q�d2*�MZ���ă��W�Im�ւ�a�R�TOR��pg�Dx�Y���LACEk��ւ�pV�ւ~�_MA�2�v�������TCV��؁��T��ي���@��t�V����V�Jj�R�MA�i�J��m�u�)b����q2j�#аU�{�t�K�JK��V�K;���H���3��J�0����JJ��JJ��AAL��ڐ��ڐ�Ԗ4Օ5���N1����ʋƀW�LP�_�(�g�,��pr��{ `�`GROUw`���B��NFLI�C��f�REQUI;RE3�EBU��qB���w�2����p��x�q5�p�� \��/APPR��C}�Y��
ްEN٨CLO7��S_M��H����u�
�qu�� ���MC�����9�_MG��C�Co��`M��в�N�BRKL�N�OL|�N�[�R��_CLINђ�|�=�J����Pܔ�����������������6ɵ�̲�8k�+��q����# ��
��q)��7�PATH3�L�BàL��H�wࡠ�J�CN�CA�Ғ�ڢB�IN�rUCV�4a��-C!�UM��Y,����aE�p����ʴ�~��PAYLOA���J2L`R_AN�q�Lpp���$��M�R_F2LSHR��N�LOԡ�R����`ׯ�ACRL_@G�ŒЛ� ��Hj`�߂$HM���FL�EXܣ�qJ�u� :�����׀�������1�F1�V�j�@�R�d�v�������E����ȏڏ ����"�4�q���6� M���~��U�g�y����T��o�X��H��� ���藕?�����ǟ ِݕ�ԕ����%��7��P��J�� � �V�h�z���`AT؃採@�EL�� �S��J|�Ŝ�JE�y�CTR��~�TN��FQ��HAND_VB-���v`�7� $��F2M�����ebSW�r�'��?� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)F�QAW�Z`i�Aw�A��PX X�'pi�Dw�D��ePf�G�p�)STk�h�!x��!N��DY�p נM�9$`%Ц�H�� H�c�׎���0� ��Pѵڵ�������t��J��� ����1��R�6��QAS�YMvř���v��pJ���cі�_SH>� �ǺĤ�ED����������J�İ%��C�I\Dِ�_VI�!X|�2PV_UNIX�FThP�J��_R�5_R c�cTz�pT�V��@��� İ�߷��U ��������Hqpˢ���aEN,P3�DI�����O4d�`J�S� x g"IJAA�a z�aabp�coc�`a�p�dq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a�i�T�@<� $D�UMMY9Q�$7PS_��RFC��;$v � ���Pa� XƠ����STE���SBR�Y�M21_VF�8�$SV_ERF�O���LsdsCLRJtA���Odb`O�p �� D $GgLOBj�_LO����u�q�cAp�r�@aS;YS�qADR``�`TCH  �� ,��ɩb�W_N�A���7����TSR���l ���
*?�&Q� 0"?�;'?�I)?�Y)�� X���h���x������) ��Ռ�Ӷ�;��Ív��?��O�O�O�D�XS�CRE栘p��f��ST��s}y`�����/_HAΗq� TơgpTYP�b���G�aG�j��Od0IS_�䓀e�UEMd�# ����ppS�qa�RSM_�q*eUNEXCEP)fW�`S_}pM�x���g�z�8����ӑCOU��S��Ԕ 1�!�UE�&��Ubwr��PRO�GM�FL@$CUgpPO�Q��5��I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp��OUS�� �� @6p�v$BU�TTp�RpR�CO�LUMq�e��SE�RV5�PANE|H�q� � �@'GEU���Fy��?)$HELPõ)B/ETERv�)ෆ� ��A � ��0`��0��0ҰIN簊�c�@N��IH�1��_� �v��LN�r� �qprձ_ò=�$H���TEXl����F�LA@��RELVB��D`��������M��?,�ű�m�����"�USRVwIEW�q� <6p�`U�`�NFI<@;�FOCU��;�7PRI@m�`�Q�Y�TRIP�qm��UN<`Md� x#@p�*eWARN)e�6�SRTOL%���g��ᴰONCOR�N��RAU����T����w�VIN�Le�� $גPA�TH9�גCACH���LOG�!�LI�MKR����v���HwOST�!�bz�R��OBOT��d�IM>� �� ����Zq�Zq;�V�CPU_AVAIYL�!�EX	�!AN���q��1r��1r���1 �ѡ�p� � #`C����@$�TOOL�$��_wJMP� ���e$SS�����VSHIF��Nc߃P�`ג�E�ȐR�����OSUR��Wk`RADILѮ��_�a��:�9a��`a�r���LULQ$OUTPUT_BM����IM�AB �@�r�TILSCO��C7����� ��&��3��A��@�q���m�I�2G��ϑV�pLe�}��yD�JU��N�WA�IT֖�}��{�%�! NE�u�YBO��� �� �$`�t�SB@T;PE��NECp�Jp^FY�nB_T��R�І�a$�[Yĭc	B��dM���F� `�p�$�pb�OP?�wMAS�_DO�!QT�pD��ˑ#�%��p!"DELAY�:`7"JOY�@(� nCE$��3@ �xm��d�pY_[�!"�`�"��[���P? �ϑZABC%�� � $�"R��
�ϐ�$$CLAS>������!pxϐ� � VIRT]ќ�/ 0ABS����1� 5� < �! F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $�6HZi{0-�AX�L�p2��!�63  ��{tIN��qztP#RE�����v�p�u�LARMRECO�V 9�rwtN�G�� .;	 �A   �.�0PoPLIC��?5��p�Ha�ndlingTo�ol o� 
V�7.50P/23~-�  �Pf���
��_SWt� �UP�!� x�F�0��t���Aϐv�� 864�� �it�y� r��" 7D�A5�� �� �Qf@��o�Ngoneisͅ˰ ��T���!�LAex>�_�l�V�uT��s9�U�TO�"�Њt�y��HGAPON
0g�1z��Uh�D 1581����̟ޟxry����Q 1���p�,�蘦����;�@��q_��"=�" �c�.��H���D�HTTHKYX��"�-� ?�Q���ɯۯ5���� #�A�G�Y�k�}����� ��ſ׿1�����=� C�U�g�yϋϝϯ��� ��-���	��9�?�Q� c�u߇ߙ߽߫���)� ����5�;�M�_�q� �������%���� �1�7�I�[�m���� ������!����- 3EWi{��� ���)/A Sew����/ ��/%/+/=/O/a/ s/�/�/�/�/?�/�/ ?!?'?9?K?]?o?�? �?�?�?O�?�?�?O#O]���TO�E�W��DO_CLEAN������CNM  � �__/_�A_S_�DSPDR3YR�O��HIc��M@�O�_�_�_�_oo +o=oOoaoso�o�o���pB��v �u���a�X�t������9�PL�UGG���G��U�P�RCvPB�@���_�orOr_��SEGF}�K[mwxq �O�O�����?rqLAP�_�~q�[� m��������Ǐُ�����!�3�x�TOT�AL�f yx�USE+NU�p�� �H����B��RG_STR�ING 1u�
_�Mn�S5��
ȑ_ITEM1Җ  n5�� � �$�6�H�Z�l�~��� ����Ưد���� ��2�D�I/O �SIGNAL̕�Tryout �ModeӕIn�p��Simula�tedבOut���OVERR~�P = 100֒�In cycl���בProg OAbor��ב���StatusՓ	�Heartbea�tїMH Fa�ul��Aler '�W�E�W�i�{ύϟ�p�������� �C Λ�A����8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|���WOR{pΛ��(ߎ� ���� ��$�6�H�Z� l�~�������������p�� 2PƠ �X ��A{��� ����/A Sew�����SDEV[�o� #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1?�C?U?g?y?PALTݠ1��z?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_�?GRI�`ΛDQ�? _l_~_�_�_�_�_�_ �_�_o o2oDoVoho@zo�o�o�o2_l�R� �a\_�o"4FX j|����������0�B�T��oPREG�>�� f��� Ə؏���� �2�D� V�h�z�������ԟ����Z��$ARG�_��D ?	����;��  	$Z�W	[O�]O��Z��p�.�SBN_CONFIG ;�ꎱ����CII�_SAVE  �Z�����.�TCE�LLSETUP �;�%HOM�E_IOZ�Z�%�MOV_��
�R�EP�lU�(�UTOoBACKܠ���FRA:\�z� \�z�Ǡ'�`�z���ǡi�I�NI�0z���~n�MESSAG����ǡC���ODE_!D������%�O�4��n�PAUSX!�~;� ((O>� �ϞˈϾϬ������ ����*�`�N߄�r��߶�g�l TSK � wͥ�_�q�UP3DT+��d!�AſWSM_CF���;���'�-�GRgP 2:�?� N��BŰA��%�XSC�RD1�1
7� 	�ĥĢ�������� ��*�������r��� ��������7���[� &8J\n��*�>t�GROUN�UϾ�UP_NA��:�	t��_ED��17�
 �%�-BCKEDT�-�2�'K�`�ܵu�z�q�,q�z���2t1�����q�k�(/��ED3/��/��.a/�/;/M/ED4�/t/)?�/.?p?�/�/ED5`??�?�<?.�?O�?�?ED6O�?qO�?.MO�O'O9OED7�O`O_��O.�O\_�O�OEDa8L_,�_�^-p�_ oo_�_ED9�_�_]o�_	-9o�oo%oCR_ 9]��oF�o�k� � NO�_DEL��GE?_UNUSE���LAL_OUT �����WD_ABORﰨ~��pITR_RTN�=��|NONSk����˥CAM_PARAM 1;��!�
 8
SO�NY XC-56� 2345678�90 ਡ@����?��( �А\�
���{��:��^�HR5q�̹���ŏR57ڏ�A�ff��KOW�A SC310M�
�x�̆�d @<�
���e�^ ��П\����*�<���`�r�g�CE_R�IA_I�!��=�F��}�z� ]��_LIU�]�V����<��FB��GP 1���Ǯ�M�_�q�0�Cg*  ����C1���9��@��G���CVR�C]��d��l��Es��R�����[ԴUm��v�������_�� C����(������=�HE�`O�NFIǰ�B�G_�PRI 1�{ V���ߖϨϺ�����������CHKPA�US�� 1K� ,!uD�V�@�z�d� �߈ߚ��߾������.��R�<�b���OƯ�������_MkOR�� �6��� 	 �����*��N�<�����H��?��q?;�;����R��K��9�P���>ça�-:���	�

��M���p U�ð��<��,~���DB���튒)
�mc:cpmidcbg�f�:����s��p�/� ' �Q�	� �,s>܋�3Q��?􋐒�Yg �/�مXf�M/�w�O/�
DEF �l��s)�< b?uf.txts/��t/��ާ�)�	`z�����=L���*[MC��1����X?43��1��t�~īCz  BHH�ދ�B�$�y6��y��.�4D��Y�D���/�4E�CeYF��Y��,�'w�1���s�U��.�p�����1�BDw�M@x8�K�cCҨ��0fADȷ0��0E�?EX��EQ�EJP �F�E�F� �G��=F^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE ���F 
Q��;��(P  B_<_��Rb����	op6C4P)�Y
s@ ]AQ�2Js@C�0B3�MaC{@�@*cw��UT�pFPROG %�z�o�oigI�q���v���ldKEY_TBL�  �&S�#� �	�
�� !�"#$%&'()�*+,-./01�i�:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇���������������������9��p`LCK�l4�<p`�`STAT ��S�_AUTO_DO��5�INDTO_ENB!���R�Q�?�1�T2}�^�STsOPb���TRLr`�LETE��Ċ_�SCREEN ��Zkcsc���U��MMENU� 1 �Y  <�l�oR�Y1�[� ��v�m���̟����� ٟ�8��!�G���W� i��������ïկ�� 4���j�A�S���w� ����迿�ѿ���� T�+�=�cϜ�sυ��� �ϻ�������P�'� 9߆�]�o߼ߓߥ��� �����:��#�p�G� Y����������� $����3�l�C�U��� y����������� ���	VY)�_MAN�UAL��t�DBC�O[�RIG�DOBNUM� ��B1� e
�PXWOR/K 1!�[�_�U/4FX�_A�WAY�i�GC�P  b=�Pj_A!L� #�j�Y��܅t `�_�  1"�[_ , 
�o�d�&/~&lMZ�I�dPx@P@#ONT�IMه� d��`&�
�e�MOT�NEND�o�RECORD 1(�[qg2�/{�O��! �/ky"?4?F?X?�( `?�?�/�??�?�?�? �?�?)O�?MO�?qO�O �O�OBO�O:O�O^O_ %_7_I_�Om_�O�_ _ �_�_�_�_Z_o~_3o �_Woio{o�o�_�o o �oDo�o/�oS �oL�o����@ ���+�yV,�c� u��������Ϗ>�P� ����;�&���q��� 򏧟��P�ȟ�^�� ����I�[����� � ��$�6�������j�TOLERENC�wB���L���� CS_CFG �)�/'dM�C:\U�L%04�d.CSV�� cl��/#A ��CH��z� //.ɿ��(�S�RC_OUT �*���SG�N +��"���#�28-JAN�-20 15:1�9015l�0:5�1+ P/V�t�ɞ�/.��f�p�a�m��PJ�PѲ��VERS�ION Y�V2.0.84,�EFLOGIC {1,� 	:�ޠ=�ޠL��PR?OG_ENB��".p�ULSk' �����_WRSTJN�K ��"fEMO_�OPT_SL ?�	�#
 	R575/#=������0�B����TO � �ݵϗ��V_VF EX�d�%��PATH AYʇA\�����5+IkCT�Fu-��j�#eg�S�,�STBF_TTS�(�	d���l#!:w�� MAU��z�.^"MSWX�.��Q4,#�Y�/�
!J �6%ZI~m���$SBL_FA�UL(�0�9'TD�IA[�1<�� ����1234?567890
��P��HZl~� ������/ /@2/D/V/h/�� P� ѩ�yƽ/�� 6�/�/�/??/?A? S?e?w?�?�?�?�?�?p�?�?�,/�UMP��f�� �ATR��8��1OC@PMEl�OO�Y_TEMP?�Ç��3F���G�|DU�NI��.�YN_B�RK 2_�/�E�MGDI_STA���]��ENC2_S_CR 3�K7 (_:_L_^_l&_�_�_`�_�_)��C�A14_ �/oo/oAoԢ�B�T5�K�ϋo~o l�{_�o�o�o' 9K]o���� �����#�5��/ V�h�z��л`~����� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T��� x���������ү��� ��,�>�P�b�t��� ������ο���� (�f�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������:� �2�D�V� h�z���������� ��
��.�@�R�d�v� ������������� *<N`r�� �����& 8J\n����� �����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?��?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__�NoETMODE �16�5�Q �d�X
X_j_|Q��PRROR_PR�OG %GZ%��@��_  �UTAB_LE  G[�?�oo)oRjRRSE�V_NUM  <�`WP�QQY`��Q_AUTO_ENB  �eOS�Tw_NOna 7G[��QXb  *�*�`��`��`��`d`�+�`�o�o�o�dHI�SUc�QOP�k_AL�M 18G[ �2A��l�P+�ok@}�����o_Nb.�`  G[�a�R�
�:PTCP_VE/R !GZ!�_��$EXTLOG_7REQv�i\��SIZe�W�TOL�  �QDzr��A W�_BWD��p��xf́t�_DIn�� 9�5�d��T�QsRֆSTEP���:P�OP_D�Ov�f�PFAC�TORY_TUN�wdM�EATUROE :�5̀rQ�Handl�ingTool ��� \sfm�English �Dictiona�ry��roduAA Vis�� Master��ީ�
EN̐nalog I/O��ީ�g.fd̐ut�o Softwa�re Update  F OR��matic Ba�ckup��H59�6,�ground Editޒ�  1 H5�Camera�F���OPLGX�elyl𜩐II) X�7ommՐshw���7com��co����\tp���pan}e��  opl���tyle sel�ect��al C�nJ�Ցonit;or��RDE���tr��Relia�b𠧒6U�Dia�gnos(�푥�5�528�u��he�ck Safet�y UIF��En�hanced Rob Serv%��q ) "S�r�U?ser Fr[������a��xt. D�IO �fiG� �sŢ��endx�Ekrr�LF� pȐ�ĳr됮� ���� � !��FCTN /Menu`�v-�ݡ|���TP Inې�fac�  ER_ JGC�pב_k Exct�g���H558��igh�-Spex�Ski~1�  2
P���?���mmunic�'�ons��&�l�uqr�ې��ST Ǡ���conn��2ި�TXPL��nc=r�stru�����"FATKA�REL Cmd.� LE�uaG�54�5\��Run-T�i��Env��d�
!���ؠ++�s�)�S/W��[�LicenseZ��� 4T�0�ogB�ook(Syڐm�)��H54O�MA�CROs,\�/O�ffse��Loa��MH������r,� k�MechStop Prot����� lic/�MiвShif����ɒ�Mixx��)���x�StS�Mode �Switch�� �R5W�Mo�:�.�� 74 ����g��K�2h�ult�i-T=�M���LN (Pos�Regiڑ������|d�ݐt Fun��⩐.�����Numx~����� lne�|�ᝰ Adjup������  - W���tatuw᧒T��RDMz�o}t��scove U�9���3Ѓ�uest 492�b*�o�����62;�?SNPX b ����8 J7`���Li3br��J�48����"�� �Ԅ�
�6O��� Parts i�n VCCMt�3�2���	�{Ѥ�J9�90��/I� 2� P��TMILI�B��H���P�A�ccD�L�
TE�$TX�ۨ�ap1�S�Te����pke�y��wգ�d���Unexcep=tx�motnZ���������є�� qO���� 90J��єSP CSXC`<�f��Ҟ� Py�sWe}���PRI��>vr�t�menz�� ��iPɰ�a�����vGri=d�play��v���0�)�H1�M-�10iA(B20�1 �2\� 0\}k/�Ascii��l�Т�ɐ/�Col���ԑGuar� �
�� /P-�ޠ"Kv��st{Pat �:�!S�Cyc��΂�orie��IFn8�ata- quҐ��� ƶ��mH57m4��RL��am����Pb�HMI D�e3�(b����PC�Ϻ�Passwo�+!��"PE? Sp�$�[���tp��� vKen��Tw�N�p��YELLOW B�OE	k$Arc��v�is��3*�n0W�eldW�cialh�7�V#t�Op�����1y� 2F�a�portN�(�p�T1�T� �� �ѳxy]�&TX��t�w�igj�1� b� �ct\�JPN �ARCPSU P�R��oݲOL� S;up�2fil� &�PAɰאcro�� �"PM(����O$SuS� eвtex�ԣ r���=�t�s'sagT��P���P@�Ȱ�锱�rt�W��H'>r�dpn��n1
t�!�� z ��ascbi?n4psyn��+A}j�M HEL��NCL VIS �PKGS PLOA`�MB �,�4�VW�RIPE �GET_VAR {FIE 3\t���FL[�OOL: �ADD R729.FD \j8'�iCsQ�QE��DVvQ��sQNO WTW�TE��}PD  ��^��biRFOR ���ECTn�`��ALSE ALAfP�CPMO-130�  M" #h�D�: HANG F�ROMmP�AQfr���R709 DR�AM AVAIL?CHECKSO!���sQVPCS SU��@LIMCHK �Q +P~dFF PO�S��F�Q R59�38-12 �CHARY�0�PR�OGRA W�SwAVEN`AME�P�.SV��7��$E�n*��p?FU�{�TR}C|� SHADV0�UPDAT KC|JўRSTATI�`~�P MUCH y��1��IMQ MO?TN-003��}��ROBOGUIDE DAUGH�a8���*�tou�����I� Šhd�ATH|�PepMOVET��ǔVMXPACK� MAY ASS�ERT�D��YCL�fqTA�rBE C�OR vr*Q3rA�N�pRC OPToIONSJ1vr̐PSH-171Z@-x�tcǠSU1�1`Hp^9R!�Q�`_T�P���'�j�d{tb�y app wac 5I�~d�PHI����p�aTEL�MX?SPD TB5bLu� 1��UB6@�qEN�J`CE2�61��p���s	�may n��0� R6{�R� >�Rtraff)��� 40*�p��fr���sysvar ?scr J7��cNj`DJU��bH �V��Q/�PSET �ERR`J` 68���PNDANT �SCREEN U�NREA��'�J`D��pPA���pR`IgO 1���PFI�p}B�pGROUN�P�D��G��R�P�QnRS�VIP !p�a�PD�IGIT VER�S�r}BLo�UEW~ϕ P06  �!��MAGp�abZV��DI�`� SS�UE�ܰ�EPL�AN JOT` D�EL�pݡ#Z�@D�͐CALLOb�Q �ph��R�QIPN�D��IMG�R7{19��MNT/�PWES �pVL�c���Hol�0Cq���tP�G:�`C�M�caynΠ��pg.v�S�: 3D mK�v_iew d�` �p���ea7У�b� o�f �Py���ANN�OT ACCESGS M��Ɓ*�t47s a��lok��Flex/:�Rw�!mo?�PA?�-�����`n�pa S�NBPJ AUTO-�06f����TB���PIABLE1q �636��PLN:Y RG$�pl;pNW7FMDB�VI���t�WIT 9x�0@o���Qui#0�ҺPN� RRS?pUSB��� t & remov�@ )�_��&�AxEPFT_=� �7<`�pP:�OS�-144 ��h qs�g��@OST� �� CRASH �DU 9��$�P�pW� .$��L/OGIN��8&�J���6b046 issue 6 Jg���: Slow ��st��c (HCos`�c���`IL`�IMPRWtSPO�T:Wh:0�T�S�TYW ./�VMGqR�h�T0CAT��hos��E�q���� �O�S:+pRSTU' k�-S� ����E:��pv@�2�N� t\hߐ��m ���all��0�  �$�H� WA͐��3 CNT0 T��� WroU�alacrm���0s�d � @�0SE1���r R{�OMEBp���K� �55��REàSEs�t��g    } �KANJI��no���INIS?ITALIZ-p�d�n1weρ<��dr�� lx`�SCI�I L�fail�s w�� ��`�YSTEa���o��PvЧ IIH���1W�G�ro>Pm ol\�wpSh@�P��Ϡn� cflxL@АW{RI �OF Lq���p?�F�up��d�e-rela�d� "APo SY�c}h�Abetwe:0IND t0$gb#DO���r� `��GigE�#ope�rabilf  P�AbHi�H`��c�le{ad�\etf�P8s�r�OS 030��&: fig��GL�A )P ��i��7�Np tpswx�B��If�g�������5aE�a EXC�E#dU�_�tPCLO�S��"rob�NTdpFaU�c�!����PNIO V750�Q1��Qa��'DB ��P M�+Pv�QED�DET���-� \rk��ON�LINEhSBUG�IQ ߔĠi`Z�IB�S apABC �JARKYFq� ����0MIL�`� R��pNД �p0GAR��D*pR��P�"'! jK�0cT�P��Hl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P��`WIBPK05��!FȐB/��BUSY RUNN��C "�򁐈��R-p��LO�N�DIV�Y�CUL��fsfoaBW�p����30	V��ˠIT�`�a505.�@O=F�UNEX�P1bҬaf�@�E��SVwEMG� NMLq�� D0pCC_SA�FEX 0c�08"qD. �PET�`N@�#'J87����RsP�TA'�M�K�`K��H GUNCHG^۔MECH�pMcz� T�  y, g@��$ ORY LE�AKA�;�ޢSP�Em�Ja��V�tGR�Iܱ�@�CTLN�TRk�FpepR��j50�EN-`IN�����p �`�Ǒ�k!��T3/dqo�SKTO�0A�#�L�pA �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`D	U��aO�supk�t4� � P�F� Bnf��Q�PSVGN-18��V�SRSR)J�UP�a2�Q�#D�q� l O��QBRKCTR5Ұ�|"-��r�<pc�j!INVP�D ZO� ��T`�h#�Q�cHset,x|D��"DUAL� �w�2*BRVO117 A]�TNѫt�+bTa2473��q.?���sAUz�i�B�complete���604.� -^�`hanc�U�� F��e8��  ��npJtPd!q��`��w� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP��R�R(}\xPe� aʰ�I���E��1��p�� j  �� xSt�^t �A�AxP�q �5 sig��a��"AC;a��
�bCe�xPb_p��.pc�]l<bHbcb_cicrc~h<n�`tl1� ~`xP`o�dxP�b]o2�� �cb�c�ixP�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`�cptlibxzxP�l�cr�xrxP\�blpsazEdxP_fm�} gcxP�x���o|sp�or�mc(��ob_jzo"p�u6�wf��t���wms�1q��sld�)��jmc�o\�n�b�nuhЕ��|st�e���>�pl�qp�iwc1k���uvf0uߒ<��lvisn�CgoaculwQ
E �F  ! Fc.f9d�Qv�� qw����Data Acq/uisi��nF�|1��RR631`��TR��QDMCM �2֝P75H�1�P58�3xP1��71��559`�5�P57<PxP�Q����(���Q���o pxP!daq�\�oA��@�� �ge/�etdms�"�DMER"؟,�p#gdD���.�m���-��qaq.<᡾xP#mo��h���f{�u��`13��MACRO�s, SksaffP�@z����03�SR�QT(��Q6��1�Q9ӡ��R�ZSh��PxPJ6+43�@7ؠ6�P�@�PRS�@���e �Q��UС PIK�Q5?2 PTLC�W���xP3 (��p/O ��!�Pn �xP5���03\sfmn�mc "MNMCPq�<��Q��\$AcX�FM���ci,Ҥ�X�����cdpq+�
�sk��SK�xP�SH5�60,P��,�y�r�efp "REF�p�d�A�jxP	�of��OFc�<gy�to��TO_����ٺ����+je�u��caxis2�xPE�\�}e�q"ISDTc�|�]�prax ���MN��u�b�is�de܃h�\�w�xP!� isbasic���B� P]��QA7xes�R6�������.�(Ba�Q�ess��xP���2�pD�@�z�atis�� ��(�{�����~��m��FMc�u�{�
���MNIS��ݝ�� ��x����ٺ��x�� j75��Dev�ic�� Inte�rfac�RȔQJ�754��� xP�Ne`��xP�ϐ2��б����dn� "�DNE���
tpodnui5UI��ݝ	bd�bP�q_rsofOb
?dv_aro��u�����stchkc��z	 �(}�onl��G!ff L+H�J(��"l"/��n�b��z�haSmp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!2���xpc_2pcch=m��CHMP_�|8бpevws��2�ΌpcsF��#C �SenxPacro0�U·�-�R6�Pd�@xPk�����p��gT�L��1d M�2`��8��1c4ԡ�3 qem��GEM,\i(��Dgesnd�5���H0{�}Ha�@sy���c��Isu�xD��Fmd ��I��7�4���u���AccuCal�P��4� ��ɢ7ޠB0���6+6f�6��9!9\aFF q�S(�U��2�
X�p�!Bd�ѳcb_�SaUL�� � �� ?�ܖto���otplus\tsrnغ�qb�W�p��t���1��To�ol (N. A�.)�[K�7�Z�(P��m����bfclls� k94�"K4p���qtpap� �"PS9H�stpswo��p�L7��t\�q����D�yt5� 4�q��w�q��� �Mz�uk��rkey�����s��}t�sfe7atu6�EA��� cf)t\Xq�����df�h5���LRC0�md�!�587���a�R�(����2V��8lc?u3l\�pa3}@H�&r-�Xu���t,�� �q "�q�Ot��~ ,���{�/��1c�}����y�p�r��5����S�XAg�-�y���Wj�874�- iR�Vis���Queu�� Ƒ�-�6�1$���(����u����tӑ����
�tpv�tsn "VTS�N�3C�+�� v\pR�DV����*�prd�q\�Q�&�vst�k=P������nmx&_�դ�clrqν���get�TX��Bd���aoQϿ�0q�str�D[� ��t0�p'Z����npv��@�enlIP0��D!0x�'�|���sc ߸��tvo/��2�q���vb����q����!���h]��(� Control�PRAX�P5��5�56�A@59�P5-6.@56@5A��J69$@982 �J552 IDVR7�hqA���16�Hx���La�� ���Xe�frlparwm.f�FRL��am��C9�@(F �����w6{���A���QJ643�� 5}0�0LSE
_p�VAR $SGS�YSC��RS_UNITS �P�2�4�tA�TX.$VN�UM_OLD 5`�1�xP{�50+��"�` Funct ���5tA� }��`#@�`E3�a0�cڂ��9����@H5נ� �P���(�A����۶}�����ֻ}��bPR�b�߶~ppr4�TP�SPI�3�}�r�10�#;A� t�
`���1���96�����%C�� Aف��J�bIncr�	����\�`��1o5qni4�MNINp	xP�`����!��Hour_  � 2�21 �A�AVM���0 ���TUP ��?J545 ���6162�VC�AM  (��CLIO ���R6�N2�MSC� "P ��STYL�C�28�~ 13\�NRE� "FHRM S�CH^�DCS}U%ORSR {b��04 �E�IOC�1 j 5742 � os| �? egist��Ի��7�1�oMASK�934"�7 ��OCO ���"3�8��2���� 0 HB��ڢ 4�"39N� R�e�� �LCHK�
%OPLG%��3�"%MHCR.%MCd  ; 4? ��6 d�PI�54�s� D[SW%MD� pQ�K!637�0�0p"�Y1�Р"4 �6<2?7 CTN K � +5 ���"7��<2�5�%/�T�%FRD�M� �Sg!��9�30 FB( NBA��P� ( HLB  7Men�SM$@jB�( PVC ��290v��2HTC�C?TMIL��\@?PAC 16U�hA�J`SAI \@ELN���<29s�UE�CK �b�@FRM� �b�OR���I�PL��Rk0CSXsC ���VVFna}Tg@HTTP �N!26 ��G�@~obIGUI"%�IPGS�r� H863 qb�!�07r�!�34 �r�84 �\so`! Qx`CC3� Fb�21�!969 rb!51 ���!S53R% 1!s3!���~�.p"9js V{ATFUJ775"���pLR6^RP�WS�MjUCTO�@xT5�8 F!80���1X�Y ta3!770 ���885�UOL�  GTSo
�{` L�CM �r| TSS��EfP6 W�\@CPgE `��0VR� �l�QNL"��@00�1 imrb�c3� =�b�0���0�`6� w�b-P- R-��b8n@5EW�b9 �Ґa� ���b�`ׁ~�b2 2000���`3��`4*5�`5 !�c�#$�`7.%�`�8 h605? U�0�@B6E"aRp76� !Pr8 t�a�@�tr2 iB/d�1vp3�vp5 ȂRtr9Σ�a4@-pN�r3 F��r5&0�re`u��r7 ��r�8�U�p9 \h7�38�a�R2D7�"�1f��2&�7<� �3 7iC���4>w5Ip�Or60� C�L�1bEN�4 I�pyL�uP��@N�&-PJ8�N�8NeN�C9 H�r`�E�b7]�|���8�ВࠂG9 2��a`0�q�Ђ5�%U097 �0��@1�0���1� (�q�3 5R ���0���mpU���0�0�7*�H@(q��\P"RB6�q124�b;��@���@�06� x�3 pB�/x�u ��x�6 H606�a1� ��7 6 ���p��b155 ����7>jUU162 ��3 g��4*�65 2e "_��P�4#U1`���B1���`=0'�174 �q���P�E186 R L��P�7 ��P�8&��3 (�90 B�/�s191����@2s02��6 3���A�RU2� d��O2 b2h`��4��b��2�4���19v RQ�2��u2d�Tpt)2� ��H�a2hP�$2�5���!U2�p�p"
�2�p��@5�0-�@��8 @�9��T�X@�� �e5�`rb	26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0@�gqGA���a�52ѐ�Ḳ6�6�0ہ5� ׁ2��84�E��9�EU5@ٰE\�q5hQ`S�2ޖ5�p\w�۲�pJ �4-P��5�p1\t�H�-4��PCH�7j��phiw�@��P�x��?559 ldu� P �D���Q�@�������A �`.��P>��8�g581�"�q58�!�AM۲T�A iC�a589��@�x���F�5 �a��12׀ 0.�1���,�2�����,�!P\h8��Lp ���,�7��6�084�0\� ANRS 0C}A��p��{��sran��FRA�� �Д�е���A%�� �ѹ�Ҍ�����(�� ��Ќ���З���������ь����$�G��1��ը��������� xS�`�q�  �����`6�4��M��iC/50T-H������*��)p46��� C��xN����m75s֐�� Sp��b46���v����ГM-7�1?�7�З����4A2������C��-��F��70�r�E��/h����O$��rlD���c7c7C� q��Ѕ���L��/���2\imm7c7�g������`���(��e�����"� �������a r��&c�T,�Ѿ�"��,��� ��x�Ex�m7�7t����k���5������)�iC��-HS-� B
_� >���+�Т�7U�]P���Mh7�s��a7������-9?�?/260L_������Q�������]�9pA/@���q�S�х��^�h621��c��92������.�)92c0�g$�@������)$��5$���pcylH"O"
�21�8��t?�350� ���p��$�
�� F�350!���0�x�9�U/0\m9��M9A3��4%�� s��3M$��X%u<���"him98J3����� i d�"m4~��103p�� ����h�794̂�&R���H �0����\���g�5A U��՜��0���*2� �00��#06�а�Ճ�է!07{r  ��������kЙ@�����EP�#�������?��#!�;&0s7\;!�B1P��@�A��/ЁCBׂ2�!��:/��?�ҽCD25�L����0�"l�2BL
#��B��\20�2_�r�re� ��X��1��N����A@��z��`C�pU��`��04��Dy	A�\�`fQ��s�U���\�5  ��� p�^t��<$85���+P=�ab1l��1LT��lA8�!uDnE(�.20T��J�1 e�bH85���b�Ռ�5[�16Bs��������d2��x��m6t!`Q����b�ˀ���b#�(�6iB ;S�p�!��3� ���b�s��-`�_�W80�_����6I	$�X5�1�U85��R�p6S����/�/+q�!@�q��`�6o��5m[o)�m6sW��Q�|�?��set06p h��3%H�5��10p$@����g/�JrH��?  ��A��856����F�� ���p/2��h�܅�✐)�5��̑v�𘜐(��m6��Y�H�ѝ̑m�6�Ҝ��ae6�DM����-S�+��H2�����Ҽ� � �r̑��✐��l���p1���F����2�\t6h T6H����Ҝ�'Vl ���ᜐ�V7ᜐ/�(���;3A7��p ~S��������4�`堜��V���!3��2��PM[��%ܖO�chn��vel5���8�Vq���_arp#���̑�.���2l_h�emq$�.�'�6415���5���?����F�����5g�L�ј�[���1��𙋹1<����M7NU�Р���eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h������ u���㜐��ZS0�!ܑ4���M-����S�$̑�ք �� 0���<�����07shJ�H�v�À�sF� �S*󜐳���̑���vl�3�A�T�#��Q�0��Te��q�pr����T@75j�5�dd�̑ 1�(UL�&�(�,���0��\�?���̑�a�� xSt���a�eD�w�2��(�	�2�C��A/���\�+p�<����21 (ܱ�CL S����B̺@��7F���?�<�lơ1L����c� ���u19�0����e/q���O���9�K��r9 (��,�Rs�ז�5�<G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O���M1!41w���2T@� _std��G�y�� �ң�H� jdgm����w0\� �1L� ��	�P�~�W*�b���t 5������3�,���E{���d���L��5\L��3�L�|#~���~!���4�#��O����h�L6A�������a2璥���44������[6\j4s ��·���#��ol�E"w�8Pk�����?0x j�H1�1Rr�>��]�2a�2Aw�P ��	2��|41�8��ˡ��@{� �%�A<��� +� ?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R�� ˑb�W���Fs���) �ѐ�!���a�1�����5��16�16C���C����0\imBQ��d����b��\Be5�-���DiL����O�_�<ѠPEtL �E�RH�ZǠPgω�am1l��u���̑�b@�<����<�$�T� ̑�F����Ȋ�DpbĜ�X"�ᒢ��pĻ ���^t��9��0\� j971\�kckrcfJ�F�s�����c��e "CTME�r�����!|�a�`main.[�8�g�`run}�_vc�#0�w�1Oܕ�_u����bctme���Ӧ�`ܑ�j73�5�- KARE�L Use {�U���J��1���p� Ȗ�9�B@���L�9��7j[�atk208 "K��(Kя��\��9��a���̹����cKRC4�a�o ��kc�qJ� &s�����Grſ�fs�D��:y��s��A1X\�j|хrdtB�, L��`.v�q�� �spǑIf�Wfj52��TKQuto Seut��J� H5K7536(�932���-91�58(�9�BA��1(�74O,A$�(TCP Ak���/�)Y� �\tpqtool.v���v���! con�re;a#�Cont�rol Re�b{le��CNRE(� T�<�4�2���D�)���NS�552��q(g�� (򭂯4X�cOux~�\sfuts�UTS`�i�栜���At�棂��? 6�T�!�SA OO+D6���������,!��6c+� igt�t6i��I0�T�W8 ���la��vo58�o�bFå򬡯i��Xh��!Xk�0Y!8�\m6e�!6EC���v��6���������<16�A���A�6s����U�g�T|�,����r1�qR����Z4�T�����,#�eZp)g����<ONO0���uJ��tCR;��F<�a� xSt�f���prdsuchk� �1��2&&?���t��*D%$�r(�✑ �娟:r��'�s�qO��<scrc�C�\At�trldJ"o��\�V����Pay�lo�nfirm�l�!�87��7��A�3ad�! �?@ވI�?plQ��3���3"�q��x pl��`���d7��l�calC�uDu���;���mov�����initX�:s8O��a8�r4 ��r67A4|��e Genera#tiڲ���7g2q$g R� (S�h��c ,|�bE��$Ԓ\�:�"���4��4�4�. sg��5�F$d6"�e�!p "SHA�P�TQ ngcr pGC�a(�&"� ���"GDA¶��r�6�"aW�/�$d�ataX:s�"tp�ad��[q�%tput;a__O7;a�o8�1�yl+s�r�?�:�#$�?�5x�?�:c O�:Ay O�:�IO�s`O%g�qǒ�?�@0\ۜ�"o�j92;!�Pp�l.Collis�QSkip#��@5� �@J��D��@\ވ�C(@X�7��7�|s}2��ptcls�#LS�DU�k?�\_� ets�`�< �\�Q��@���`dcKLqQ�FC;��J,όn��` (��4eN����T�{���' j(�c�q���/IӸaȁ<��̠H������зa�e\mcc�lmt "CLM��/��� mate\v��lmpALM�?>p7qmc?�����2vm�q��%�3s��_�sv90�_x_msu�2L^v_� K�o��{in�8(3r<�c_logr��r�trcW� �v_3�~yc��d�<�ste��der$c;Ce� Fiρ��R��Q�?�l�enter߄|��(�Sd��1�TX�+fZK�r�a99sQ9+��5�r\tq\� _"FNDR����STDn$�LANG�Pgui��D⠓�S������csp�!ğ֙uf䟀ҝ�s����$�����e +�=����������������w�H�r\fn�_�ϣ��$`x�tcp�ma��- TCP������R638 aR�Ҡ��38��M7p,���Ӡ�$Ӡ��8p0Р�VS,�>�tk��99�a��B3���P�զԠ��D�2�����UI��t���hqB���8���������p���re8�ȿ��exe@4π��B���e38�ԡG�r�mpWXφ�var @�φ�3N�����v�x�!ҡ��q�R�BT $cOP�TN ask E�0��1�R MAS�0�H593/�96g H50�i�480ԅ5�H0��m�Q�K(��7�0�g�Pl�h�0ԧ�2�ORDP���@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`am��b��7�.f���u�d��r��splayD�E���1wПUPDT Ub��8o87 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60�q��B����qs�can��B���aAd@�������q`� �䗣�#��К�`2�� vlv��Ù�$�0>�b���! S���Easy/К�Ut�il��룙�511# J�����R7 ���Nor֠��inc�),<6Q�� �`c��"4�[���986(FVRx So����q�nd6����P��4� a\ (��
  ������"�d��K�bdZ����men7���- Me`tyFњ�Fb��0�TUa�577?i3R��\�5�au?��!� n����f������l\m�h�Ц�űE|h#mn�	��<\O�$��e�1�� l!���y��Ù�\|p�����B���Ћmh �@��:.aG!�� �/�t�55�6�!X��l�.us��Y/k)eOnsubL���eK�h�� �B\1;5g?�y?�?�?D��?*rmx�p�?Ktbox O�2K|?�G��C?A%das���?1ӛ#� � TR��/��P�4B�`�U@�P�V�P"�Q�P0�U �PO��P�"�T3�U�P �f�Pk"�2}�4�T�P �f�P2�"�Q5�S�Q@���R?Ă�Q3t.�PF׀al��P+O�n�P517��IN0a���Q(}g��PES	Tf3ua�PB�l�i�g�h�6�aq��P �� xS��` � n�0mbump�P�Q969g�69�Qq��P0�baAp�@>Q� BOX��,�>vche�s�>ve�tu㒣=wffse�3���]�;u`aW��:zol�sm<u�b�a-��]D�K�ib�Q�c����Q<twaǂ �tp�Q҄Taror Recov�br�O�P�642�����a�q��a⁠QErǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>��pjot��PXc��C��1�adb -�ail���nag���b�QR629�a�Q��b�P�  �
 � �P��$$CL~[q ����������$�PS?_DIGIT���"�!�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��������*璬1:P�RODUCT�Q0�\PGSTK�bV�,n�99�\����$FEAT_INDEX���~�� �搠ILECOM�P ;��)���"��SETUPo2 <��?�  N !��_AP2BCK �1=�  �)}6/E+%,/i/��W/�/~+/�/O/ �/s/�/?�/>?�/b? t??�?'?�?�?]?�? �?O(O�?LO�?pO�? }O�O5O�OYO�O _�O $_�OH_Z_�O~__�_ �_C_�_g_�_�_	o2o �_Vo�_zo�oo�o?o �o�ouo
�o.@�o d�o���M� q���<��`�r� ���%���̏[���� ���!�J�ُn����� ��3�ȟW������"� ��F�X��|����/� ��֯e������0��� T��x������=�ҿ �s�ϗ�,ϻ�9�b�t� P/ 2) *.VRiϳ�!�*���������Ɲ�PC�7�!�F'R6:"�c��χ��T��߽�Lը����x���*.F���>� �	N�,�k�x�ߏ��STM �⠸���Qа���!��iPendant? Panel���H��F���4������GIF�������pu����JPG&�P��<����	�PANEL1.D	T��������2�Y�G��
3w�����//�
4�a/��O///�/�
TP�EINS.XML�/���\�/�/�!�Custom T?oolbar?��PASSWOR�D/�FRS:�\R?? %Pa�ssword Config�?��? k?�?OH�6O�?ZOlO �?�OO�O�OUO�OyO _�O�OD_�Oh_�Oa_ �_-_�_Q_�_�_�_o �_@oRo�_voo�o)o ;o�o_o�o�o�o*�o N�or��7� �m��&���\� ����y���E�ڏi� �����4�ÏX�j��� �����A�S��w�� ���B�џf������� +���O��������� >�ͯ߯t����'��� ο]�򿁿�(Ϸ�L� ۿpς�Ϧ�5���Y� k� ߏ�$߳��Z��� ~�ߢߴ�C���g��� ��2���V����ߌ� ��?����u�
��� .�@���d������)� ��M���q�����< ��5r�%�� [�&�J� n��3�W� ��"/�F/X/�|/ /�/�/A/�/e/�/�/ �/0?�/T?�/M?�?? �?=?�?�?s?O�?,O >O�?bO�?�OO'O�O KO�OoO�O_�O:_�O ^_p_�O�_#_�_�_Y_��_}_o�_�_Ho)f��$FILE_DG�BCK 1=���5`��� ( �)
S�UMMARY.DyGRo�\MD:�o��o
`Diag� Summary��o�Z
CONSLOG�o�o�a
J�a�ConsoleO logK�[�`�MEMCHECK�@'�o�^qMe�mory Dat�a��W�)>�qHADOW����P��sShad�ow Chang�esS�-c-��)	FTP=��9�����w`qmmen�t TBD׏�W0�<�)ETHERNET̏�^�q��Z��aEther�net bpfiguration[���P��DCSVRF�ˏ��Ïܟ�q%��� verify� allߟ-c1P{Y���DIFFԟp��̟a��p%��diffc���q���1X�?�Q�� �����X��CH�GD��¯ԯi��px��� ���2`�G�Y��� ��� �GAD��ʿܿq��p���Ϥ�FY3h�O�aώ�� ��(�GAD������y��p�����0�UPDAT�ES.�Ц��[FORS:\�����a�Updates �List���kPS�RBWLD.CM�.��\��B��_pP�S_ROBOWEL���_����o��,o !�3���W���{�
�t� ��@���d�����/ ��Se����� N�r� =� a�r�&�J� ��/�9/K/�o/ ��/"/�/�/X/�/|/ �/#?�/G?�/k?}?? �?0?�?�?f?�?�?O �?OUO�?yOO�O�O >O�ObO�O	_�O-_�O Q_c_�O�__�_:_�_ �_p_o�_o;o�__o �_�o�o$o�oHo�o�o ~o�o7�o0m�o � ��V�z� !��E��i�{�
��� .�ÏR���������� .�S��w������<� џ`������+���O� ޟH������8���߯�n����$FIL�E_��PR����������� �MDONL�Y 1=4�� 
 ���w�į�� 诨�ѿ�������+� ��O�޿sυ�ϩ�8� ����n�ߒ�'߶�4� ]��ρ�ߥ߷�F��� j�����5���Y�k� �ߏ���B�����x� ���1�C���g���� ��,���P����������?��Lu�VI�SBCKR�<�a��*.VD|�4 OFR:\��4 �Vision VD file�  :LbpZ�# ��Y�}/$/� H/�l/�/�/1/�/ �/�/�/�/ ?�/1?V? �/z?	?�?�???�?c? �?�?�?.O�?ROdOO �OO�O;O�O�OqO_ �O*_<_�O`_�O�__�%_�_�MR_GR�P 1>4�L~�UC4  B�P�	 ]�ol`��*u����RHB ��2 ���� ��� ���He�Y�Q`ork bIh�oJd�o�Sc�o��oE�� L��K-�F�{5U�aS&.��o��osB���A��b �Q6����;o{0  >�>@�lqhr:ގ�xq�o� F@ �r�d�aX}J��N�Jk�H9��Hu��F!��/IP�sX}?�`��.9�<9���896C'�6<,6\b�X1�,.�g�R���v�A�PA�����|� ݏx���%��I�4� F��j�����ǟ��� ֟��!��E�`r�UBH�P�c�������ů�R
6�P;�kP<z�˯R��e�Q� cB��P5���@'�33@���4�m�^,�@UUU��U�~�w�>u.�?!x�^��ֿ���3���=[z�=����=V6<�=��=�=$q���~��@8�i�7G��8�D��8@9!��7ϥ�@Ϣ���cD��@ D�� CYώ���C��P��P'�6��_V� m�o�� To��xo�ߜo����� �A�,�e�P�b��� �����������=� (�a�L���p������� ����������*��N 9r]����� ���8#\n Y�}������ �/ԭ//A/�e/P/ �/p/�/�/�/�/�/? �/+??;?a?L?�?p? �?�?�?�?�?�?�?'O OKO6OoO�OHߢOl� �ߐߢ��O�� _��G_ bOk_V_�_z_�_�_�_ �_�_o�_1ooUo@o yodovo�o�o�o�o�o �oNu �������� �;�&�_�J���n��� ����ݏȏ��%�7� I�[�"/�描����� ٟ�������3��W� B�{�f�������կ�� �����A�,�e�P� b��������O�O�O ��O�OL�_p�:_�� ���Ϧ��������'� �7�]�H߁�lߥߐ� �ߴ�������#��G� 2�k�2��Vw���� �������1��U�@� R���v����������� ��-Q�u� ��r��6�� )M4q\n� �����/�#/ I/4/m/X/�/|/�/�/ �/�/�/?ֿ�B?� f?0�BϜ?f��?���/ �?�?�?/OOSO>OwO bO�O�O�O�O�O�O�O __=_(_a_L_^_�_ �_�_���_��o�_o 9o$o]oHo�olo�o�o �o�o�o�o�o#G 2kV{�h�� �����C�.�g� y�`����������Џ ���?�*�c�N��� r��������̟�� )��M�_�&?H?���? ���?�?�?����?@� I�4�m�X�j�����ǿ ���ֿ����E�0� i�Tύ�xϱϜ����� ����_,��_S���w� b߇߭ߘ��߼����� ��=�(�:�s�^�� ���������'� 9� �]�o����~��� ����������5  YDV�z��� ���1U@ yd��v����� /Я*/��
/�u/� �/�/�/�/�/�/�/? ?;?&?_?J?�?n?�? �?�?�?�?O�?%OO IO4O"�|OBO�O>O�O �O�O�O�O!__E_0_ i_T_�_x_�_�_�_�_ �_o�_/o��?oeowo �oP��oo�o�o�o �o+=$aL�p �������'� �K�6�o�Z������ ɏ��폴� ��D� / /z�D/��h/ş�� �ԟ���1��U�@� R���v�����ӯ���� ��-��Q�<�u�`� ��`O�O�O���޿� �;�&�_�J�oϕπ� �Ϥ��������%�� "�[�F��Fo�ߵ��� �ߠo��d�!���W� >�{�b�������� ������A�,�>�w� b����������������=��$FN�O ����\�
�F0l q  FL�AG>�(RRM�_CHKTYP � ] ��d ��] ��OM� _�MIN� 	����� �  XT S�SB_CFG �?\ ����O�TP_DEF_O/W  	��,�IRCOM� >��$GENOVRD7_DO��<�l�THR� d�d�q_ENB] �qRAVC_GR�P 1@�I X(/ %/7//[/ B//�/x/�/�/�/�/ �/?�/3??C?i?P? �?t?�?�?�?�?�?O OOAO(OeOLO^O�O.oROU�F\� �,�B,�8�?���O�O��O	__���  DaE_�Hy_�\@@m_B�=�vR/��I�O�WSMT�G�SU�oo&oRHOST�C�1H�I� Ĺ�zMSM��l[bo�	1�27.0�`1�o  e�o�o�o #z�oFXj|�l6�0s	anonymous�����F��)ao�&�&��o�x��o������ ҏ�3��,�>�a� O����������Ο�U %�7�I��]����f� x��������ү��� �+�i�{�P�b�t��� ���������S� (�:�L�^ϭ�oϔϦ� �������=��$�6� H�Zߩ���Ϳs����� ������ �2���V� h�z��߰������� ��
��k�}ߏߡߣ� ���߬���������C� *<Nq�_�� ����-�?�Q�c� eJ��n���� ���/"/E� X/j/|/�/�/� %'/?[0?B?T?f? x?��?�?�?�?�?? E/W/,O>OPObO�KDa�ENT 1I�K� P!�?�O  �P�O�O�O�O�O#_ �OG_
_S_._|_�_d_ �_�_�_�_o�_1o�_ ogo*o�oNo�oro�o �o�o	�o-�oQ u8n����� ���#��L�q�4� ��X���|�ݏ���ď�֏7���[���B�?QUICC0��h�z�۟��1ܟ��ʟ+��2,���{�!?ROUTER|�X��j�˯!PCJO�G̯��!19�2.168.0.�10��}GNAME� !�J!RO�BOT�vNS_C�FG 1H�I ��Aut�o-starte�d�$FTP�/ ���/�?޿#?��&� 8�JϏ?nπϒϤ�ǿ ��[������"�4ߵ& ����������濜��� �������'�9�K�]� o����������� ��/�/�/G���k��� �������������� 1T���Py�� ���"�4�	H- |�Qcu�VD� ���/�;/M/ _/q/�/����/
/ �/>?%?7?I?[?*/ ?�?�?�?�/�?l?�? O!O3OEO�/�/�/�/ �?�O ?�O�O�O__ �?A_S_e_w_�O4_._ �_�_�_�_oVOhOzO �O�_so�O�o�o�o�o �o�_'9Kno �o�����o*o <oNoP5��oY�k�}� ����pŏ׏���� 0���C�U�g�y���_��T_ERR J�;�����PDUSI�Z  ��^P�����>ٕWRD �?z���  �guest ���+�=�O�a�s�*��SCDMNGRPw 2Kz�Ð���۠\��K��� 	P01.�14 8�q  � y��B    ;�����{ �����������������������~ �ǟI�4�m�X��|��  i�  �  
����� ����+��������
����l�.x��
��"�l�ڲ۰s��d�������_G�ROU��L�� e��	��۠07K�QUPD  ����PČ�TYg������TTP_A�UTH 1M��� <!iPen'dan���<�_��!KAREL�:*�����KC�%�5�G��VISION SETZ���|��Ҽߪ��� ������
�W�.�@����d�v���CTRL� N�������
��FFF9E�3���FRS:DEFAULT��FANUC �Web Server�
������q�������������W�R_CONFIGw O�� ����IDL_CPU�_PC"��B���= �BH#MI�N.�BGNR_�IO��� ���% N�PT_SIM_D�Os}TPMO_DNTOLs �_PRTY�=!OLNK 1P���'9K]|o�MASTEr ������O_CFG���UO����C�YCLE���_?ASG 1Q���
 q2/D/V/h/ z/�/�/�/�/�/�/�/p
??y"NUM����Q�IPCH���£RTRY_�CN"�u���SC�RN������ ���R����?���$J23_D_SP_EN������0OBPROC��3��JOGV�1�S_�@��8��?�';ZO'??0CP�OSREO�KANJI_�Ϡu�A$#��3T ���E�O�ECL_LM B2e?��@EYLOGGI�N�������L�ANGUAGE Y_�=� }Q���LG�2U������ �x�����PZC � �'0������MC:\RSCH\00\˝�LN_DISP V�������T�OC�4Dz\A��SOGBOOK W+��o���o�o���Xi�o�o�o�o��o~}	x(y��	�ne�i�ekElG�_BUFF 1X���}2���� Ӣ������'� T�K�]����������� ɏۏ���#�P���~�qDCS Zxm =���%|d1h�`���ʟܟ�g�IOw 1[+ �?'����'�7�I�[�o� �������ǯٯ��� �!�3�G�W�i�{��������ÿ׿�El TM  ��d��#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U��g�yߋߝ߈t�SE�V�0m�TYP�� ��$�}�A�RS"�(_�s�2FLg 1\��0��� �����������5�STP<P���DmNGNAM�4�U�nf�UPS`GI�5��A�5s�_LOA�D@G %j%wDF��GI6����MAXUALRMB7�P8��y���3��0]&q��Ca]�s�3�~�� 8@=@^�+ طv	��V0+�P�A5d�cr���U� �����E( iTy����� ��/ /A/,/Q/w/ b/�/~/�/�/�/�/�/ ??)?O?:?s?V?�? �?�?�?�?�?�?O'O OKO.OoOZOlO�O�O �O�O�O�O�O#__G_ 2_D_}_`_�_�_�_�_ �_�_�_o
ooUo8o yodo�o�o�o�o�o�o��o�o-��D_LDXDISA^�� �MEMO_APX��E ?��
 �0y�����������ISC ;1_�� �O� ���W�i�����Ə �����}��ߏD�/� h�z�a��������� �����@���O�a� 5������������u� �ׯ<�'�`�r�Y��� ���y�޿�ۿ��� 8Ϲ�G�Y�-ϒ�}϶� ������m�����4���X�j�#�_MSTR� `��}�SCD 1as}�R���N� �������8�#�5�n� Y��}��������� ���4��X�C�|�g� �������������� 	B-Rxc�� �����> )bM�q��� ��/�(//L/7/ p/[/m/�/�/�/�/�/ �/?�/"?H?3?l?W?��?{?�?�?�?n�MK�CFG b����?��LTARM_��2cRuB� �3WpTNBpME�TPUOp�2�����NDSP_CM�NTnE@F�E�� d���N�2A�O|�D�EPOSCF�G��NPSTOL �1e-�4@�<#�
;Q�1;UK_YW7_ Y_[_m_�_�_�_�_�_ �_o�_oQo3oEo�o�io{o�o�a�ASIN�G_CHK  ��MAqODAQ2Cf�O�7J�eDEV �	Rz	MC:>'|HSIZEn@�����eTASK �%<z%$1234?56789 ��u��gTRIG 1g.�� l<u%����3���>svvYP�aq��kEM_IN�F 1h9G� `)AT?&FV0E0(����)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏ P��t�������]�ί �����(�۟�^� �#�5�����k�ܿ�  ϻ�ů6��Z�A�~� ��C���g�y������ ��2�i�C�h�ό�G� ���ߩ��ߙϫ���� ����d�v�)ߚ��߾� y��������<�N� �r�%�7�I�[���� ��9�&��J[��g��>ONIT�OR�@G ?;{ �  	EXESC1�3�2�3�E4�5��p�7�8�9�3�n�R �R�RRR R(R4R@RTLR2Y2e2qU2}2�2�2�U2�2�2�3Y�3e3��aR_G�RP_SV 1i�t��q(�5�
���5��۵MO�~q_DCd~�1PL�_NAME !�<u� �!De�fault Pe�rsonalit�y (from �FD) �4RR2�k! 1j)TEX�)TH��!�AX d�?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�Ox2-?�O�O�O__0_ B_T_f_x_�b<�O�_ �_�_�_�_�_o o2o�DoVoho&xRj" 1�o�)&0\�b, Ӗ9��b�a @oD�  �a?��c�a?�`�a�aA'��6�ew;�	l��b	 �xoJp��`��`	p �<; �(p� �.r� �K�K ���K=*�J���J���JV��k0q`q�P�x�|�� @j�@T;f�r�f�q�ac^rs�I�� ��p����p�r�ph}�3��´  ���>��ph�`z���꜖"�Jm�q� H�N��a`c��$�dw��  ��  P� Q�� �� |  ��m�Əi}	'� �� �I� �  �����:�È�È=G���(��#�a	����I  �n @H�i~�ab�Ӌ�b!�$w���"N0���  'Ж�q�p@2��@����r��q5�C�pC0C��@ C�����`
�A1]w@�B�V~X�
nwBD0h�A��p�ӊ�p@����aDz���֏࿯�Я	�pv�(� �� -���I��-�=��A�a��we_q�`�p �??�ff ��m�|�� �����Ƽ�!@ݿ�>1�  P�apv(�`ţ�� �=�qst��?˙��`x`�� <
�6b<߈;����<�ê<�? <�&P�ς��AO��c1��ƍ�?offf?O�?&���qt@�.�J<?�`��wi4� ���dly�e߾g;ߪ� t��p�[ߔ�߸ߣ� ���� ����6�wh�F0%�r�!�����1ى����E��� E�O�G+� F�!���/���?�e�`P���t���lyBL�cB��Enw4������� +��R��s���������h�yÔ�>���I�mXj���A�y�weC��������#/*/c/�N/wi�����v/C�`� CHs/`
=$��p�<!�!��ܼ�'��3A�A�AR�1AO�^?��$�?������
=ç>�����3�W
=�s#�]�;e��?������{�����<�>(��B�u���=B0�������	R��zH�F��G���G���H�U`E����C�+��}I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*O ONO9OrO]O�O�O�O �O�O�O�O_�O8_#_ \_G_�_�_}_�_�_�_ �_�_�_"oooXoCo |ogo�o�o�o�o�o�o �o	B-fQ� u������� ,��P�b�M���q��� ��Ώ���ݏ�(�� L�7�p�[������ʟ ���ٟ���6�!�Z��E�W���#1( �ٙ9�K���ĥ ������Ư!3��8���!4Mgqs��,�IB+8��J��a���{�d�d�����ȿ��쿔ڼ%P8�P�= :GϚ�S�6�h�z���R�Ϯ����������  %�� ��h� Vߌ�z߰�&�g�/9�$�������7�����A�S�e�w�   ������������̿2 F�$�&Gb��������!C���@���8������F� Dz�N�� F�P �D�������)#�B�'9K]o#?_���@@v
4$�8�8��8�.
 v��� !3EWi{�����:� ���ۨ�1��$M�SKCFMAP � ���� ���(.�ONREL  ��!9��EXC/FENBE'
#7%�^!FNCe/W$JO�GOVLIME'dtO S"d�KEYE'u�%�RUN�,��%�SFSP�DTY0g&P%9#S�IGNE/W$T1M�OT�/T!�_C�E_GRP 1p��#\x��?p� �?�?�?�?�?O�? OBO�?fOO[O�OSO �O�O�O�O�O_,_�O P__I_�_=_�_�_�_ �_�_oo�_:o��TCOM_CFG 1q	-�vo�o��o
Va_ARC_�b"�p)UAP_�CPL�ot$NOCHECK ?	+ �x�% 7I[m���������!�.+N�O_WAIT_L� 7%S2NT^ar�	+�s�_ERR�_12s	)9��  ,ȍޏ��x����&��dT_MO��t>��, K�*oq��9�PARAM��u	+��a�ß'g�{�� =?�345?678901�� ,��K�]�9�i�����`��ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDS�P�c#6p(OFFSET_CART�oη�DISƿ��PE?N_FILE尨!��ai��`OPTIO�N_IO�/��PW�ORK ve7s# ��V�ؤ!!p�p�4�p�	 ����p��<���RG_DSBL  ���P#��ϸ�RIE�NTTOD ?�Cᴭ !l�UT__SIM_D$�"����V��LCT w}�h�iĜa[�1ԟ_PEXE�j�R�ATvШ&p%� ��2�^3j)TEX)T�H�)�X d 3�������%�7�I� [�m��������������!�3�E���2 ��u���������������c�<d�AS ew������`��Ǎ�^0OUa0�o(��(�����u2, ����O H @D��  [?�aG?��cc�D][�Z��;�	ls��xJ��������<� ��� ���2�H(��H3�k7HSM5G��22G���Gpc
͜�'f�/,-,2�CR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t3�!�/ �/�"�t32����/6 W ��P%�Q%��%�|T��S62�q?�'e	'� � ��2I� � � ��+==�̡ͳ?�;	�h	�0��I  �n �@�2�.��Ov;���ٟ?&gN�]O  �''�uD@!� C�C��@F#H!�/�O�O Nsb
���@�@E��@�e`0B��QA�0Yv: �13Uwz$oV_�/z_�e_�_�_	��( �� -�2@�1�1ta�Ua�c����:Ar���.  �?�ff���[o"o�_!U�`oXÜQ8���o:�j>�1  Po�V(���eF0�f�Y����L�?����x�b�P<
6b<�߈;܍�<��ê<� <�#&�,/aA�;r��@Ov0P?fff?��0?&ip�T@�.�{r�J<?�`�u#	�Bdqt�Yc �a�Mw�Bo�� 7�"�[�F��j����� ��ُ����3�����,���(�E��� E��3G+� F��a��ҟ������,��P�;���B�pAZ�>��B��6�<O ίD���P��t�=����a�s�����6j�h�y�7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�<%?��?������(���#	Ę��P �N�||CH���Ŀx������@I�_��'�3A�A�A�R1AO�^??�$�?��� ��±
=ç>�����3�W
=�#� U��e����B��@��{�����<����(�B�u���=B0�������	�b�H��F�G���G���H�U`E����C�+��I�#�I��H�D�F��E��RC�j=[��
I��@H��!H�( E?<YD0߻� �������� �9�$� ]�H�Z���~������� ������#5 YD }h������ �
C.gR� ������	/� -//*/c/N/�/r/�/ �/�/�/�/?�/)?? M?8?q?\?�?�?�?�? �?�?�?O�?7O"O[O mOXO�O|O�O�O�O�O��O�O�O3_Q(���3���b��gUU���W_i_2�3ǭ8��_�_2�4M�gs�_�_�RIB+��_�_�a���{�miGo5okoYo(�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�u�,��  �p���o ��/��S��z
uү ܠ�������ڱ������������  /�M�w�e�������~�l2 F�$��'Gb��t��a�`�,p�S�C�y�@p�5��G�Y�۠F� D�z�� F�P D��]����پ��ʯܯ� ��~ÿ?���@@�J?�K�K���K���
 �|��� ����Ŀֿ������0�B�T�fϽ�V� ����{��1��$�PARAM_ME�NU ?3���  �DEFPULS�Er�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L��	�OPT���PTB4�.�C��R_DECSN ���e��ߑߣ����� ������!�3�\�W��i�{���USE_PROG %��q%�����CCR����e����_HOSoT !��!��:���T�`�V��/��X����_TIMqE��^��  ��?GDEBUG\�����GINP_FL'MSK����Tfp�����PGA  ��̹�)CH����TY+PE������� ����� - ?hcu���� ���//@/;/M/ _/�/�/�/�/�/�/�/��/??%?7?`?��W�ORD ?	=�	RSfu	P�NSUԜ2JO�K�DRTEy�]T�RACECTL �1x3��� �`�`&�?�3�6_DT Qy3�%@~�0D � �c2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�o&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�Z�.O|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv��p���� �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲπ����������(���$PGTRACE�LEN  )� � ���(��>�_UP _z���m�u��Y�n�>�_CFoG {m�Wӊ(�n���PЬ� ���DEFSPD �|��'�P���>�IN��TRL �}��(�8��I�PE_CONFI���~m���mњ��Ԛ�>�LI�D����=�GR�P 1��W���)�A ���&�ff(�A+33D��� D]� C�À A@1��Ѭ�(�d�Ԭ��0�0�� 	 1��1��� ´�����B �9����O�9�s��(�>�T?�
�5�������� =?��=#�
�� ��P;t_�������  Dz (�
H� X~i����� �/�/D///h/S/��/��
V7.1�0beta1���  A�E>�"ӻ�A (�� �?!G��!>���"����!����!BQ��!A\�� �!���!2p����Ț/8?J?\?n?};!� ���/��/�? }/�?�?OO:O%O7O pO[O�OO�O�O�O�O �O_�O6_!_Z_E_~_ i_�_�_�_�_�_�_' o2o�_VoAoSo�owo �o�o�o�o�o�o.�R=v1�/�#F@ �y�}��{m� �y=��1�'�O�a� �?�?�?������ߏʏ ��'��K�6�H��� l�����ɟ���؟� #��G�2�k�V���z� �������o��ί C�.�g�R�d������� ���п	���-�?�*� cώ���Ϯ��� ���B�;�f�x��� ����DϹ��߶����� ���7�"�[�F�X�� |�����������!� 3��W�B�{�f����� ���� �����/ S>wbt��� ���=Oz� �Ͼψ����ϼ�  /.�'/R�d�v߈߁/ 0�/�/�/�/�/�/�/ #??G?2?k?V?h?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O ���O�O�O__?_*_ c_N_�_r_�_�_�_�_ �_o�_)oTfx� to���/�o/ >/P/b/t/mo� |������� 3��W�B�{�f�x��� ��Տ�������A� S�>�w�b����O��џ ������+��O�:� s�^�������ͯ��� ܯ�@oRodo�o`��o �o�o��ƿ�o���* <N�Y��}�hϡ� ���ϰ��������
� C�.�g�Rߋ�v߈��� ������	���-��Q� c�N�ﲟ���l��� �����;�&�_�J� ��n����������� ,�>�P�:L������ ������(�:� 3��0iT�x� ����/�/// S/>/w/b/�/�/�/�/ �/�/�/??=?(?a? s?��?�?X?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O* \&_8_r���_�_���$PLID_�KNOW_M  ���| Q�TSV ����P� �?o"o4o�OXoCoUo��o R�SM_GROP 1��Z'0{`��@�`uf�e�`
�5� �gpk 'Pe]o� ��������V�SMR�c��mT�EyQ}? yR������ ����폯���ӏ�G� !��-����������� 韫���ϟ�C��� )�����������寧����QST�a1 1Ն�)���P0� A 4��E2�D� V�h�������߿¿Կ ���9��.�o�R�dπvψ��ϬϾ����2r�0� Q�<3߂�3�/�A�S��4 l�~ߐߢ��5���������6
��.�@��7Y�k�}���8��������MAD  )���PARNUM  �!�}o+��SCHE� S�
��f���S��UPDf�x���_CMP_0�`H�� �'�U�ER_CHK-����ZE*<RS8r��_�Q_MOG���_�X�_RES_G��!���D� >1bU�y� ����/�	/����+/�k�H/ g/l/��Ї/�/�/� 	��/�/�/�X�?$? )?���D?c?h?�����?�?�?�V 1�x�U�ax�@c]�@}t@(@c\�@}�@D@c[�*@���THR_IN�Rr�J�b�Ud2FM�ASS?O ZSGM�N>OqCMON_QUEUE ��UX�V P~P X�N$ �UhN�FV�@ENqD�A��IEXE�O��E��BE�@�O�CO�PTIO�G��@P�ROGRAM %�J%�@�?���B?TASK_IG�6^OCFG ��Oxz��_�PDATA�c]��[@Ц2=� DoVohozo�j2o�o�o �o�o�o);M^ jINFO[��m��D����� ���1�C�U�g�y� ��������ӏ���	�4dwpt�l )�Q~E DIT ��_|i��^WERFLX�	C�RGADJ ��tZA�����?�נʕFA��IORI�TY�GW���MPGDSPNQ����U�GyD��OTOE@�1�X� (!�AF:@E� c�Ч�!tcpn����!ud����!�icm���?<�XYm_�Q�X���Q)� *�1�5��P��]�@�L���p� �������ʿ��+�@=�$�a�Hυϗ�*��OPORT)QH��P��E��_CAR�TREPPX��S�KSTA�H�
SS�AV�@�tZ	2500H863��P�_x�
�'��X�@�swPtS�ߕߧ�^��URGE�@B��6x	WF��DO�F"�[W\�������WR�UP_DELAY� �X���R_HOTqX	B%�c����R_NORMAL�q^R��v�SEMI������9�QSKI�P'��tUr�x 	7�1�1��X�j� |�?�tU���������� ����$J\n 4������� �4FX|j �������/ 0/B//R/x/f/�/�/��/tU�$RCVT�M$��D�� DC�R'���Ў!=��Bv�4C� V�>�.>�z�6:e�:��������6��:�o?��� <
6b<�߈;܍�>u�.�?!<�&�?h?�?�?�@>� �?O O2ODOVOhOzO �O�O�O�O�O�?�O�O __@_+_=_v_Y_�_ �_�?�_�_�_oo*o <oNo`oro�o�o�o�_ �o�o�o�o�o8J -n��_���� ���"�4�F�X�j� U������ď���ӏ ���B�T��x��� ������ҟ����� ,�>�)�b�M������� �����ïկ�Y�:� L�^�p���������ʿ ܿ� ����6�!�Z� E�~ϐ�{ϴϗ����� -�� �2�D�V�h�z� �ߞ߰���������
� ��.��R�=�v��k� ����������*� <�N�`�r��������� ��������&J \?������ ��"4FXj�|��!GN_AT�C 1�	; �AT&FV0�E0�ATD�P/6/9/2/�9�ATA��,AT%G1�%B960�W+++�,�H/�,�!IO_TYPOE  �%�#t��REFPOS1� 1�V+ x	�u/�n�/j�/ 
=�/�/�/Q?<?u??��?4?�?X?�?�?�+2 1�V+�/�?�?�\O�?�O�?�!3 1�O*O<OvO�O�O_>�OS4 1��O�O��O_�_t_�_+_S5 1�B_T_f_�_o�	oBo�_S6 1� �_�_�_5o�o�o�oUoS7 1�lo~o�o��oH3l�oS8 1�%_����SMASK ;1�V/  
?�M�N�XNOS/�r�������!MOTE � n��$��_CFG� ����q���"P?L_RANG������POWER 壧���SM_�DRYPRG �%o�%�P��TA�RT ��^�U?ME_PRO-�?�����$_EXEC_?ENB  ���GSPD��Րݘ���TDB��
�RM\�
�MT_'�T�����OBOT_NAME o�����OB_OR�D_NUM ?��b!H863  �կ����PC_T�IMEOUT�� �x�S232Ă1��� LT�EACH PEN�DAN��w���-��Main�tenance �Cons���s�"����KCL/C�m��

���t�ҿ �No Use�-��Ϝ�0�NPO��򁋁���.�CH_L���̫��q	��s�MA�VAIL�����������SPACE1w 2��, j�@߂�D��s�߂� ��{S�8�?� k�v�k�Z߬��ߤ��� �� �2�D���hߊ� |��`������� ��� �2�D��h�� |���`���������y�
��2����0�B� ��f�����{���3);M _������/� /44FX j|*/���/�/�/ ?(??=?5Q/c/ u/�/�/G?�/�/�?O@�?$OEO,OZO6n? �?�?�?�?dO�?�?_�,_�OA_b_I_w_7 �O�O�O�O�O�_�O_ (oIoo^oofo�o8�_�_�_�_�_�oo 6oEf){����G �o�� ���
M�  ���*�<�N�`�r��� ����w���o�収���d.��%�S�e� w�����������Ǐَ ���Θ8�+�=�k�}� ������ůׯ͟��� �%�'�X�K�]����� ����ӿ�������#�E�W� `� @�������x�����\�e�������� ���R�d߂�8�j߬� �߈ߒߤ�������� ��0�r���X���� ��������8�����
�ύ�_MOD�E  �{��S ���{|�2�0� ����3�	S|�)CWORK_A�D����+R  �{�`� ��� _INTVAL����d���R_OPoTION� ���H VAT_GR�P 2��u�p(N� k|��_��� ��/0/B/��h�u/ T� }/�/�/�/�/�/ �/?!?�/E?W?i?{? �?�?5?�?�?�?�?�? O/OAOOeOwO�O�O �O�OUO�O�O__�O =_O_a_s_5_�_�_�_ �_�_�_�_o'o9o�_ Iooo�o�oUo�o�o�o �o�o�o5GYk -���u��� ��1�C��g�y��� M�����ӏ叧�	�� -�?�Q�c��������� ������ǟ�;��M�_����$SCAN_TIM��_%�}�R �(ӿ#((�<04�d d 
!D�ʣ��u�a/�����U�E�25���@�d5�"P�g��]	����������dd�x�  �P���� ��  8� ҿ�!���D��$�M�_� qσϕϧϹ�������p�ƿv���F�X��/� ;��ob��pm��?t�_DiQ̡>  � l�|� ̡ĥ�������!�3� E�W�i�{������ ��������/�A�S� e�]�Ӈ��������� ����);M_ q������� r���j�Tfx �������/ /,/>/P/b/t/�/�/�/�/�/�%�/  0 ��6��!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O*�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko�O�OJ�o�o�o�o �o�o�o 2DV hz������0�
�7?  ;�>� P�b�t���������Ǐ ُ����!�3�E�W��i�{�������ß �ş3�ܟ��&�8� J�\�n�����������a�ɯ����,�� �+�	12345678�ү 	� =5����f�x��������� ����
��.�@�R� d�vψϚ�៾����� ����*�<�N�`�r� �߳Ϩߺ�������� �&�8�J�\�n�ߒ� ������������"� 4�F�u�j�|������� ��������0_� Tfx����� ��I>Pb t������� !/(/:/L/^/p/�/@�/�/�/�/�/�2 �/?�#/9?K?]?�iCz  Bp˚_   ��h2���*�$SCR_G�RP 1�(�U�8(�\x}d�@ �� �'�	 �3 �1�2�4(1*�&�I3��F1OOXO}m���D�@�0ʛ)����HUK�LM-10iA 890?��90;��F;�M61C D�:�CP��1
\&V�1	�6F@��CW�9)A7Y	(R@�_�_�_�_�_�\���0i^�oOUO >oPo#G�/���o'op�o�o�o�oB�0!�rtAA�0*�  @�Bu&Xw?��ju�bH0{UzAF@ F�`�r ��o�����+� �O�:�s��mBqrr��0��������B�͏b� ���7�"�[�F�X��� |�����ٟğ���N��@�AO�0�B�CU
L����E�jqBq=���̔�$G@�@pϯ B���G�I
E�0�EL_DEFAU�LT  �T���E��M�IPOWERFL�  
E*��7�W7FDO� *��1�ERVENT 1O���`(�� �L!DUM_E�IP��>��j!?AF_INE�¿�C�!FT���丿�!o:� ���a�!RPC_OMAINb�DȺPϜ��t�VIS}�Cɻ�����!TP��P�U�ϫ�d��E�!
�PMON_PROXYF߮�e4ߑ���_ߧ�f����!R?DM_SRV�߫�9g��)�!R�Iﲰ�h�u�!
v�M�ߨ�id���!R�LSYNC��>��8���!ROS��4��4��Y�(�}� ��J�\����������� ��7��["4F �j|����!��Eio�ICE�_KL ?%�� (%SVCPRG1n>���3�"�3���4//"�5./3/�6V/[/�7~/�/��D�/�	9�/�+�@��/� �#?��K?��s? � /�?�H/�?�p/ �?��/O��/;O� �/cO�?�O�9?�O �a?�O��?_��? +_��?S_�O{_� )O�_�QO�_�yO�_ ��Os����>o �o}1�o�o�o�o�o�o �o;M8q\ �������� �7�"�[�F��j��� ����ُď���!�� E�0�W�{�f�����ß ���ҟ���A�,� e�P���t���������ί�y_DEV ���MC�:��_!�O�UT��2��REC 1�`e�j�w �	 � ����˿���ڿ��
 �`e���6�N� <�r�`ϖτϦ��Ϯ� ������&��J�8�n� ��bߤߒ��߶����� ��"��2�X�F�|�j� ������������� �.�T�B�x�Z�l��� ����������, P>`bt��� ���(L: \�d�����  /�$/6//Z/H/~/ l/�/�/�/�/.��/? �/2? ?V?D?f?�?n? �?�?�?�?�?
O�?.O @O"OdORO�OvO�O�O �O�O�O�O__<_*_ `_N_�_�_x_�_�_�_ �_�_oo8oo,ono \o�o�o�o�o�o�o�o �o "4jX� �������� �B�$�f�T�v����� �������؏��>��,�b�P�r���p�V 1�}� P
�ܟ�� A��TYPE�\��HELL_CFG �.�F�͟�  	�����RSR������ӯ�� �����?�*�<�u� `�����������ο�  �%@�3�E��Q�\���1M�o�p��d���2��d]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&��1�OW_REG�_UI���IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he�#�� ������������) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������n���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( �}��>Pbt�� ,���� �;M_q��( ����//�7/ I/[/m//�/$/�/�/ �/�/�/?�/3?E?W?�i?{?�? :&cop�y mc:dio�cfgsv.io� md:=>in�spiron:2260�?�?�?	O>�0�2frs:or�derfil.d�at virt:?\temp\�?`O�rO�O�O)1(.F*.dBOTHWO�O�O_;�
xyzrate 61 �O�O�On_�_�_%5.WOMH_Z_��_�_o"83.O@HmpbackNOboto܆o�o }*�3db�@*CoUjYo�o�o6!9.x.d:\�o8p@Rm�on��%5/.ua6HZq_��� '_���n������_>�Y3400 H�Z� ����"o4o�o��a� s������oE���Y�������z.�@OUe99�2 ޟo�����&4' �OH�Z�V�������0_¯ԯe�w���> ��W�G�Y�����!92.�@�O�`�rτϖ�)1)��I�سX������ :-.A�T���m� ߑ�$�G�۰]���  ��%�7�����l�~� ��ϵ���Y������ !�3���W�h�z����� ��B�������
�/� A�S�dv���H ����+���O� `r����:��_ �//'����n/��/�/���Y1844 ǏY/�/�/?!�3� �(a?s?�?�?��E?�(�Y?�?�?O!8�$S�NPX_ASG �1����9A�� P 0� '%R[?1]@1.1O 9?�#3%dO�OsO�O �O�O�O�O�O __D_ '_9_z_]_�_�_�_�_ �_�_
o�_o@o#odo GoYo�o}o�o�o�o�o �o�o*4`C� gy������ �	�J�-�T���c��� ����ڏ�����4� �)�j�M�t�����ğ ������ݟ�0��T� 7�I���m�������� ǯٯ���$�P�3�t� W�i��������ÿ� ���:��D�p�Sϔ� wω��ϭ��� ���$� ��Z�=�dߐ�sߴ� �ߩ������� ��D� '�9�z�]������ ����
����@�#�d� G�Y���}��������� ����*4`C� gy����� �	J-T�c� �����/�4/ /)/j/M/t/�/�/�/ �/�/�/�/?0?4,D�PARAM ��9ECA �	U��:P�4�0$H�OFT_KB_CFG  p3?E�4�PIN_SIM  9K�6�?�?�?��0,@RVQSTP/_DSB�>�21O|n8J0SR ��;� & =O{Op0��6TOP_ON_ERR  p4��9�APTN ��5�@A��BRING_PR�M�O J0VDT_GRP 1�Y9�@  	�7n8_ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2Dk hz������ �
�1�.�@�R�d�v� ��������Џ���� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\����������� ȯگ����"�I�F� X�j�|�������Ŀֿ ����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�tߛ� �ߪ߼��������� (�:�a�^�p���� �������� �'�$�6� H�Z�l�~���������������3VPRG_�COUNT�6�8�A�5ENB�O�M=�4J_UPD� 1��;8  
p2����� � )$6Hql ~�����/� / /I/D/V/h/�/�/ �/�/�/�/�/�/!?? .?@?i?d?v?�?�?�? �?�?�?�?OOAO<O NO`O�O�O�O�O�O�O �O�O__&_8_a_\_�n_�_�_�_YSDOEBUG" � �P�dk	�PSP_PA�SS"B?�[L�OG ���m�P�X�_  ��g�Q
MC:�\d�_b_MPC m��o�o�Qa�o� �vfSAV žm:dUb�U�\gSV�\TEM_TIME 1�� (�PF�TNu]�qT1SVGUNYS} #'k�sp�ASK_OPTICON" �gosp�BCCFG ���| �b��z`����4��X�C� |�g�����ď֏���� ��	�B�-�f�Q�c� ���������ϟ�� ,�>�)�b��YR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz��rBr�|�|� ���z� �%��I� 4�m�X���|������� �֏���3��W�B� g���x�����՟���� ����S�>�w�b� ����'2A ��ʯܯ�� ����E�0�i�T��� x���ÿտ翢���� /��?�e�1�/���/ �ϜϮ��������,� �P�>�`߆�tߪߘ� �߼��������L� :�p�^������� ����� �6�H�>/`� r�������������� �� 0Vhz8 ������
 .�R@vd�� �����//</ */L/r/`/�/�/�/�/ �/�/�/�/?8?&?\? J?�?n?�?�?�?�?�� �?OO�?FO4OVOXO jO�O�O�O�O�O�O_ _�OB_0_f_T_v_�_ �_�_z_�_�_�_oo >o,oboPoroto�o�o �o�o�o�o(8 ^L�p���� ���$��H�6�l� ~�(O����f�d��؏ ���2� �B�D�V��� ����n����ԟ
��� .�@�R�d����v��� �����Я���*�� N�<�^�`�r�����̿ ���޿��$�J�8� n�\ϒπ϶Ϥ����� ��ߊ�(�:�L���|� jߌ߲ߠ��������� �0�B�T��x�f�� ������������,� �P�>�t�b������� ��������:( JL^����� � �6$ZH ~l��^���d� � //D/2/h/V/x/ �/�/�/�/�/�/�/? 
?@?.?d?v?�?�?T? �?�?�?�?�?OO<O *O`ONO�OrO�O�O�O �O�O_�O&__6_8_ J_�_n_�_�_�_�_�_ �_�_"ooFo��po �o,oZo�o�o�o�o �o0Tfx�H �������,� >��b�P���t����� ����Ώ��(��L� :�p�^�������ʟ�� �ܟ� �"�$�6�l� Z���~�����دꯔo ��&�ЯV�D�z�h� ������Կ¿��
�� .��R�@�v�dϚτ��  ���� ��������$TBJ�OP_GRP 2�ǌ�� � ?������������_xJBЌ���9� �< ��X���� @����	 �C��} t�b  C��<��>��͘Ր���>̚йѳ33�=�CLj�f�ff?��?�ff�BG��ь�����t��ކ�>�(�\�)�ߖ�E噙�;���hCYj�� � @h��B�  �A����f��C�  Dhъ�1���O�4�N����
:���Bl^���j�i�l�l����A�ə�A�"��D9��֊=qH����нp�h�Q�;�A�j��o��@L��D	2��������$�6�>B��\��T���Q�ts>x�@33@���C���y�1�����>��Dh�����x�����<{�h�@i� ��t ��	���K& �j�n|��� p�/�/:/k/������!��	V�3.00J�m61cI�*� IԿ���/�' Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I�!CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;��;Q�T,8�4`� *�ϴ?�2����3\�X/O��ESTPARS  ���	���HR@ABL/E 1����0�É
H�7 8��9
GB
H
H����
G	
HE

H
HYE��
H�
H
H6FRD	IAO�XOjO|O�O�O�ETO"_4[>_P_�b_t_�^:BS _�  �JGoYoko}o�o�o�o �o�o�o�o1C Ugy����`#o RL�y�_�_�_�_�O�O��O�O�OX:B�rNUoM  ���P��� V@P:B_CFG ˭��Z�h�@��IMEBF_TT%AU��2@��VERS�q���R 1���
 �(�/����b�  ����J�\���j�|��� ǟ��ȟ֟����� 0�B�T���x�������R2�_���@�
��MI_CHAN��� � ��DBGL�V���������E�THERAD ?U��O������h�����ROUT6�!��!����~��SNMASKD�|�U�255.���#�����OOLO_FS_DI%@�u�.�ORQCTRL �����}ϛ3r� �Ϲ���������%� 7�I�[�:���h�z߯��APE_DETA�I"�G�PON_S�VOFF=���P_?MON �֍��2��STRTCH/K �^������VTCOMPAT���O�����FPRO�G %^�%  BCKEDT-Q�<��9�PLAY&H��_INST_Mްe ������US��q��LCK���Q?UICKME�=�ރ�SCREZ�>G�tps� �� �u�z����_��@@�n�.�SR_GRP� 1�^� �O����
��+ O=sa�쀚 �
m������L/ C1gU�y �����	/�-/�/Q/?/a/�/	1?234567�0�/��/@Xt�1���
� �}ipnl�/� gen.htm�? ?2?D?V?`�Panel _setupZ<}P���?�?�?�?�?�?  �??,O>OPObOtO�O �?�O!O�O�O�O__ (_�O�O^_p_�_�_�_ �_/_]_S_ oo$o6o HoZo�_~o�_�o�o�o �o�o�oso�o2DV hz�1'�� �
��.��R��v����������ЏG���U�ALRM��G ?9� �1�#�5� f�Y���}�������џ�ן���,��P��S�EV  �����ECFG ���롽�A�� :��Ƚ�
 Q��� ^����	��-�?�Q��c�u�����������Ԇ� �����I2��?���(%D�6�  �$�]�Hρ�lϥϐ� �ϴ�������#��Gߌ��� �߿U�I�_Y�HIST 1}��  (��� ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1����(�:�� ����962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V