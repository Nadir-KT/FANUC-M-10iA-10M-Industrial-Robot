��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1�~FPCUREQ1� � $SO{FT; T_ID��TOTAL_EQf� $� � NO��PS_SPI_I�NDE��$�X��SCREEN_�NAME ^�SIGN���� PK_FIL~	$THKYM�PANE�  	$DUMMY )� u3|4|G�RG_STR1� � $TIT�P$I��1��{�����5��6�7�8�9�0��z���T��1�1�1 '�1
'2"GSBN�_CFG1  �8 $CNV_�JNT_* |$�DATA_CMN�T�!$FLAG�S�*CHECK��!�AT_CEL�LSETUP � P $HO_ME_IO,G�}%�#MACRO�"�REPR�(-DR�UN� D|3S�M5H UTOBA�CKU0 � ?$ENAB��!oEVIC�TI� � D� DX�!2ST� ?0B�#$�INTERVAL�!2DISP_UNsIT!20_DOn6�ERR�9FR_F�!2IN,GRE5S�!0Q_;3!4C_WA�471�8G�W+0�$Y $D�B� 6COMW�!2MO� H.	� \rVE�1$qF�RA{$O��UDcB]CTMP1_5FtE2}G1_�3�B\�2���AXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6*_�7_�8_�94� w�CO�$ <� ��o�o�hK3 1#`O_�Mc@AC t 2� E#6NGPvABA� �c1�Q8��`,��@nr1�� d��P�0e�]p� cvnpUP&Pb26���p��"J�p_R�rPBCb��J�rĘߜJV�@ U� B��s}�g1�"Yt�P_*0OFS&R; @� RO_K8T��aIT�3T�NOMI_�0�1p�30?��D �� Ќ@�2�hPV��mEX�p� Ĝ0g0ۤ�p�r
$�TF�2C$MD3&i�TO�3�0U� F�/ ��Hw2tC%1(�Ez�g0#E{`"F�"F�40CP@��a2 �@$�PPqU�3N)ύLRևAX�!DU�v�AI�3BUF�F8=�@1 |pp��ցpPIT� PP��M�M�y��F>�SIMQSI�"�ܢVAڤT��A@�w T�`(zM��P�B^�qFACTb�@EW�P1�BTv?��MC� �$�*1JB`p�*1DE�C��F���=��� �H0CHNS�_EMP1�$G��8��@_4�3�p|@P��4�TCc�(r/� 0-sx��ܐ� MBi���!����JR� i�S/EGFR��Iv �a�R�TpN�C��P�VF4>�bx &��f{uJc!�Ja ��� !28�ץ�AJ����SIZ�3S�c�B�T�M���g��JaRSINFȑb���q�۽��н����L�3�B����CRC�e�3CC p����c��mcҞb��1J�cѿ�.����D
$ICb�Cq�5r�ե�0�@v�'���EV���zUF��_��F,pN��
ܫ�?�4�0A�! �r���h�Ϩ� �p�2�͕a�� �د��R�Dx �Ϗ��o"27�!ARtV�O`C�$LG�pV�B�1�P��@�t�a!A�0'�|�+0Ro�� MEp`"1 C3RA 3 AZV�g46p�O �FCCb�`��`F�`K������ADI��a�A�bA�'�.p��p�`�c�`S04PƑ�a�AMP��-`IY�3P�M�]pUR���QUA1  $@TITO1/S@S�!�����"0�DBPXW�O��B0!5�$SiK���2@DBq��!"�"�PR��� 
� =����!# �S q1$2�$z���L�)$�/���R� %�/�$C�!&?��$ENE�q.'�*?�Ú RE�p2(�H ��O�07#$L|3$$�#�B�[�;���FO_D��ROSr�#�������3RIGGE�R�6PApS����E�TURN�2�cMR-_8�TUw��0�EWM��M�GN�P���BLAH�<E��y�P��&$P�" �'P@�Q��CkD{��DQ���4�1���FGO_AWAY�B�MO�ѱQ#!��DCS_�)  �PIS� I gb @{s�C��A��[ �B�$�S��AbP�@�EW�-�TNTVճ�BV �Q[C�(c`�UWr�P��J��P�$0��SAF�E���U_SV�bEOXCLU��n'ONL2��SY�*a�&�OT�a'�HI_�V�4��B���_ #*P0� 9�_z��pg p��ASG�� +nrr�@6Acc *b��G�#@E�V.iHb>?fANNUN$0.$�fdID�U�2�S�C@�`�i�a��j�f\�!�pOGI$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6�a�DM�SW�E. 8Q�KgEYI5���TM�100s�qA�vIN���Ѹ�!��/ D��H7OST_P!�rT���ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  �8	=ȳ�r�DT�k0�!1 � $|S��ESAMPL��@j�۰f璱f���I�0|��[ $SUB��k�#0�C��T�r#a�SAVʅ��c���CX��P�fP$n0E��w YN_B#2 M0Q�DI{dlpO(���9#$�R_I��� �ENC2s_S� 3  5�C߰�f�- �SpU����!4�"g�޲�19T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9�g�DSP�v��PC���r"��(���ƓV7ALUߗHE�ԕ�M+�IPճ��OP5P ��TH��֤D��P�S� �۰F���df�J� ���(�T�ET+6 }H�bLL_DUs��~a3@{��3:���O�TX"���s��0N_OAUTO�!7�pC$)�$�*��c4�*(�Cp�8�C, �"�p�&�L�� 8/H *8�LH < 6����c"�`, `Ĭ� kª�q��q��sq��T~q��7��8��9���0����1��1̺1�ٺ1�1�1 �1*�1�2(�2����U2̺2ٺ2�2�U2 �2�2�3(ʥ3��3��̺3ٺ3��3�3 �3�3��4(�ɢT�?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?�p�@P?9��5�9�E�@A�a�A�z� ;p$TP�?$VARI:�Z�n��UP2�P< ���TDe���K`Q�t�����BAC�"G= T�p��e$)_,p�bn�kp+ IFIG� kp�H  ��P�!��F@`�!>t �;E��sC�ST �D� D���c�<�� 	C��{��_����l���R  ���FO�RCEUP?b��FWLUS�`H�N>�xF ���RD_CM�@E������ ��@vMP.��REMr F�Q��@1k@���7Q
K4	9NJ�5EFFۓ:f�@IN2Q��OVO�OVA�	TRO�V���DTՀ�DTMX� ��@�
�ے_PH"p��CL��_TpE�@�pK	_(�Y_T��v(���@A;QD� �������!0tܑ0R�Q���_�a����M̝7�CL�dρRIqV'�{��EARۑIOHPC�@����B�B��CM9@���R{ �GCLF��e!DYk(M�ap#5TuDG��� �%��ʠFSSD �s?C P�a�!�1���PQ_�!�(�!1��E�3�!3�+5�&�GR)A��7�@��;�P�W��ONn��EBUG_SD2H�P{�__E A`����TERM�`5Bi5$Z �O�RI#e0C�9SMQ_�P��e0Di5r1�A�9E�9UP\�F�� -�A{�A�dPw3S@B$SEG��:� EL{UUSE.�@NFIJ�B$��;1젎4�4C$UFlP=�$,�|QR@"��_G90Tk�D��~SNST�PATx����APTHJ3Q�E�p%B`�'EC���AR$P�I�aSHFTy�A�A�H_SHORР꣦6% �0$�7PE��E�GOVR=��aPI�@��U�b �QAYLOW���IE"�r�A8��?���ERV��XQ �Y��mG>@�BN��U\��R2!P.uA�SYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC����EP;�uP;�6WOR�>@M`�0SM5T6�G3�GR��13�aPAL@���`�q�u_H � ���'TOCA�`P	P�`$OP����pѡ�`0O��R%E�`R4C�AO�p��Be�`R�Eu�h|�A��e$PWR�3IMu�RR_�cN�\�q=B I&2H���p_ADDR��H_LENG�B�q�qT�q$�R��S�JڢSS��SKN��u\�0�u̳�uٳSE�A�� R�HS��M-N�!K�����b����OLX��px����`ACRO3p J�@��X�+��Q��N6�OUP3�b_�IX��a�a1��}� ����(��H��D��`ٰ��氋�IO2S�D������`�7�L $d��`Y!�_OFFr�PR�M_���aTT�P_+�H:�M (�|pOBJ]"�p��-$��LE~Cd����N � ��֑AKB_�TqᶔS�`lH�LVh�KR"~uHITCOU��[BG�LO�q����h�����`��`S9S� ���HW�#A�:�Oڠ<`INC�PU2VISIO W�͑��n��to��to�~ٲ �IOLN��P 8��R��p�$SLob PU�T_n�$p��P�& ¢��Y F_AS:�"Q��$L�������Q  U�0	P4A0��^���ZPHY��-���x��UOI �#R `�K����$�u�"pPpk���h$��������UJ5��S-���NE6WJO9GKG̲DIS���1Kp���#T (�uAqVF�+`�CTR�C�
�FLAG2�LG�dU ���؜�~13LG_SIZ�����b�4�a��a�FDl�I`�w� m�_�{0 a�^��cg���4������Ǝ���{0��� SC#H_���a7�N�d�VW���E�"����D4��UM�Aљ`LJ�n@�DAUf�EAU�0p��d|�r�GH�ba����BOO��WL3 ?�6 IT���y0�REC��SCR ܓ�D
�\���MARGm�!��զ  ��d%�����S�����W���U� �JGM�[�MNCHJ���F�NKEY\�K��PRG��UF��7P��FWD��HL��STP��V��=@�����RS��HO`����C9T��b ��7�[�UL���6�(RD� ��2��Gt��@PO���������MD�FOCUޛ�RGEX��TU%I��I��4�@� L�����P�����`��P��NE��CA�NA��Bj�VAI�LI�CL !�UDCS_HII4��s�O�(!�S����S��Ǵ ��BU�FF�!X�?PTH$m���v`��TZ1��AtrY�?Pp��j�3��`OS1Z2Z3ZD��� � Z � ��[aE�Ȥ��ȤIDX�dP�SRrO���zA�S�TL�R}�Y&�� _Y$E�C���K�&&z�� [ LQ��+00�	P ���`#qdt
�U�dw<�~��_ \ ?��4Г�\��Ѩ#�M�C4�] ��CL�DPL��UTRQL�I��dڰ�)�$FLAG&�� 1�#�D����'B�LD�%�$�%ORGڰ5�2�PVŇV�Y8�s�T�r �#}d^� ���$6��$�%SB�`T� �B0�4�6RCLMC�4]?o?��9�9MI�p}d_� d=њRQ���DSTB�p� �;F�HHAX�R �JHdLEXCESHrpCM!p�a`��A/B�TF��`a�p=F_A7Ji��KbOttH�0K�db \Q����v$MBC�LI�|�)SREQUIR�R�a.\o�AXDEB}UZ�G2�MLt M��c�b�{P����2ANDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��X�� N&��aZ��W��SPST� �ezrLOC�RI,rp�EX<fA�p��9AAODAQ��f� XY�OND�rMF,Łf�s"��}%��e/� �8FX3@I�GG�� g ���t"��ܓs#N�s$R�a%��iL��hL�xv�@�DATA#�?pE�%�jq��Y�N�h t $MD`qI}�)nv� ytq�ytHP`�Pxu��(�zsANSW)�yt@4��yuD+�)]a��ܵ0o�i �@CU�w�V�p 0XeRR2��j Du�{Q��7B?d$CALIA@���G��2��RIN��"�<��NTE��Ck�r^�آXb]���_N�qlk���9��D���Bm��DIVFFDH�@���qnI�$V,��S�$��$Z�X�o��*����oH ?�$BELT�u!_ACCEL�.�~�=�IRC�� ����D�T�8�$PS�@�"Ly�r��#�^�S�Eы T�PAT!H3���I���3x�p�A_W��ڐ���2n�C��4�_MG��$DD��T���$FW�Rp9��I�4���DE7�PPAB�N��ROTSPE!E�[g�� J��[��C@4�y$US�E_+�VPi��S�YY���1 qYNr!@A�ǦOFF�qnǡMOU��NG����OL����INC �tMa6��HB��0HBENCS+�8q9Bp�X4�FDm�IN�Ix�0]��B��VE��#�>y�23_UP񕋳/LOWL���p� B���Du�9B#P`��x ���BCv�r�MO3SI��BMOU��@��7PERCH  ȳOV��â
ǝ� ���D�ScF�@MP����� Vݡ�@y�j��LUk��Gj�p�UPp=ó���ĶTRK�>�AYLOA�Qe� �A��x�����N`�F��RTI�A$��MO UІ�HB�BS0�p7D5����ë�Z�DU�M2ԓS_BCKLSH_Cx�k�� ��ϣ���=���ޡ< �	ACLAL"q�p�1м@��CHK� :�S�RTY���^�%E1Qq_�޴_�UM�@�C#��S�CL0�r�LMT_OJ1_L��9@H��qU�EO�p�b�_�e�k�e�SPC��u�L��N�PC�N�Hz �\P��C�0~"XT\��CN_:�N9�L�I�SF!�?�V����U�/���x�T���CB!�SH�:��E� E1T�T����y���T�f�PA ��_P��_� =������!����J6 L�@���OG�G�TORQU��ONֹ��E�R0��H�E�g_W2��ā_郅���I*�I�I��Ff`xaJ�1�~1�VC3�0BD:B�1�@SBJRKF9~�0DBL_SM�:�2M�P_DL2GRV�����fH_��d���CcOS���LNH ��������!*,�aZ���fcMY�_(�TH���)THET0��N�K23���"��C-B�&CB�CAA�B��"��!��!�&SB8� 2�%GTS�Ar�CIMa�����,4#<97#$DU���H�\1� �:Bk62�:AQ�(rSf$NE�D�`I ��B+5��$̀�!�A�%�5�7���LCPH�E�2���2S C%C%�2-&FC0JM&̀V�8V�8߀LUVJV!KV/KV=KUVKKVYKVgIH�8@FRM��#X!KH/KUH=KHKKHYKHgI�O�<O�8O�YNO�JO!KO/KO=KO*KKOYKOM&F�2�!�+i%0d�7SPBA?LANCE_o![c�LE0H_�%SP�c� &�b&�b&PFULC�h�b�g�b%�p�1k%�UTO_<��T1T2�i/�2N��"�{�t#�Ѡ�`�0�*�.�T��O�À<�v INSEG"�ͱREV4vͰl�gDIF�ŕ�1lzw6��1m��OBpq�ь�?�MI{���nL�CHWARY�_�A�B��!�$MEC�H�!o ��q�AX���P����7Ђ�`n� 
�d(�U�RO�B��CRr�H���(�MSK_f`��p P �`_���R/�k�z�����1 S�~�|�z�{���z��q�INUq�MTC�OM_C� �q � ���pO�$ONOREn����p�Ђr 8p GRle�uSD�0AB��$XYZ_DAx�1a���DEBUUqX������s z`$��wCOD�� L����p�$BU�FINDX|� � <�MORm�t $فUA��֐�Р�r�<��rG��u� � $SIMUL  S�*�Y�̑a��OBJE�`̖AD�JUS�ݐAY_	IS�D�3���_FI�=��T u 7�~�6�'��p} =��C�}p�@b�D��FRiIr��T��RO@ �\�E}'�y�OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1�0e��M��ED}�*�p ��N�PMֲ����c�w�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B��2�G�B�_�M�x� ��q�E� x �Hw��p��ATUS
W���C�0o�s��çBTM�ǌ�I��k�4��x�԰q�y �Dw�E&���@E��r��7��жЗ�EXE��ἱ�����f �q�z @w���UP�'��$�pQ�XN����������� ��PG΅{ h �$SUB����0_����!�MPWAI2v�P7ã�LOR����F\p˕$RCV?FAIL_C����BWD΁�v�DE�FSP!p | Lw���Я�\���UNI+�����H�RX�+�}_L\pP��t�P��p�}H�> *�j�(�s`~�N�`KSETB�%�J�PE �Ѓ~��J0SIZAE����X�'���S��OR��FORMA�T�`��c ��WrEeM�t��%�UX���G��PLI��p��  $ˀP_�SWI�pq�J_P�L��AL_ ������A��B��� C���D�$E���.�C_�U�� ?� � ����*�J3K0����TI�A4��5��6��MOM��������ˀB��AD������l����PU� NR�������m��� A$PI�6 q��	�����K4��)6�U��w`��S/PEEDgPG�� ������Ի�4T��� � @��SA�Mr`��\�]��MOV_�_$�npt5�H�5���1���2��@������'�S�Hp�IN�'�@�+�����4($4+T+G�AMMWf�1'�$GGET`�p���Da�z��

pLIBR>ѺII2�$HI=�_�g�t��2�&E;��(A�.� �&LW�-6<��)56�&]��v�p��V���$PDCK���q��_?�����q�&���7��4����9+� �$_IM_SR�pD�s0�rF��r�rLE���aOm0H]��0�-ܬpq��PJqUR_SCRN�FA����S_SAVE_DX��dE@�NOa�CA A�b�d@�$q�Z�Iǡ s	�I� �J�K� ��� �H�L��>�"hq� �����ɢ�� �bW^US�A�-M4���a��)q`��3��WW�I@v�_�q�.M�UAo�� � $sPY+�$W�P�vNG�{��P:��R`A��RH��RO�PL��@���q� ��s'�X;�	OI�&�Zxe ���m�G� p��ˀ�3s��O�O�O�O�O�aa�_т� |��q�d@�� .v��.v��d@��[wFv���E���%E�s;B��w�|�tP���P�MA�QUa ���Q8��1�QTH��HOLG�QHY�S��ES��qUE��pZB��Oτ�  ـPܐ(�A����v�J!�t�O`�q��u��"���FA��IROG�����Q2���o�"�x�p��INFOҁ��׃V����R�H�O�I��� (�0SLEQ������Y�3�H���Á��P0Ow0Ԟ��!E0NU���AUT�A�COPY�=�/�'��@Mg�N��=�}1������� ��RG��Á�f��X_�P�$;�(���`��W��P��@������EXT_CYC bHᝡRprÁ�r��_NAec!А���ROv`~	�� � ���POR_�1�E2��SRV �)_�I�DI��T_�k�}�'����dЇ�����5��6J��7��8i�H�SdBZ���2�$��F�p���GPLeAdA
�TAR�Б@���Pp�2�裔d� ,�0cFL`�o@YN���K�M��Ck��PW�R+�9ᘐ��DE�LA}�dY�pAD��a��QSKI�P4� �A�$�O�B`NT�} ��P_$�M�ƷF@\bIpݷ �ݷ�ݷd����� ���Š�Ҡ�ߠ�=9��J2R� ���� 4V�EX� TQQ����TQ�����p� ��`�#�RDC�V�� �`��X)�R��p�����r��m$R�GEAR_� IOBT�2FLG��fipER�DTC���Ԍ�>��2TH2NS}�O 1���G �T\0 ���u�M�\Ѫ`I�d"�REuF�1Á� l�h���ENAB��cTPE�04�]����Y� ]��ъQn#��*��"��(��|@��2�Қ�߼�@����������3���'�9�K�]�o���4�Ҝ����������� ��5�ҝ�!�3�E�W�i�{���6�Ҟ������������
��7�ҟ-?Q(cu��8�Ҡ��������SMS�KÁ�l��a��E�kA��MOTE6�����@�݂TQ�IO}5�IS�q���R�W@��� 8�pJ���TS���򘐤E�"$DSB_SIGN�1UQ��x�C\ЖtRS23�2���R�iDEVICEUS�XRSR�PARIT��4!O�PBIT�QI�O?WCONTR+�TQX��?SRCU� MpS�UXTASK�3Nx�p�0p$TATU�P!U1H �0�����p�_XPC)�$FREEFROMS	p�na�GET�0��UKPD�A�2E#P� �:��� !$USAN�na&�����ERI�0�RpRIYq5*"_j@�Pm1��!�6WRK9KD����6��QFRIE3ND�Q�RUFg�҃��0TOOL�6MY��t$LENGT�H_VT\�FIR��pC�@ˀE> +IU�FIN-RM��R�GI�1ÐAITI��$GXñ3IvFG2v7G1���p3�B�GcPR�p�1F�O_n 0��!RE��p�53҅U�TC��3A�A�FG �G(��":���e1n!��J�8�%����%]��%�� 74��X O0�L��T�3H&��8���%b453%GE�W�0�WsR�TD����T��M����Q��T]�$V 2!����1�а91�8�0U2�;2k3�;3�: ifa�9-i�aQ��NSL��ZR$V��2BVwE�V�	V�B;���� �&�S�`��F�"�k�@��2a�PS�E���$r1C��_$Aܠ6wPR��7vMU�c�S�t '�/89�� 0G�aV`��p�d`A���50�@��-�
25�S�� ��aRHW����B�&�N�SAX�!�A:@LA�h��rTHIC�1pI���X�d1TFEj�|�q�uIF_CH�3��qI܇7�Q�pG1@RxV���]��:�u�7_JF~�PRԀƱ��RVAT���� ��`���0RҦ�D9OfE��COUԱ���AXI���OFF{SE׆TRIGNS ���c����h������H�Y��IGMA�0PA�pJ�E�OR?G_UNEV�J�� �S�����d� �$CА�J�GgROU����TOށܒ!��DSP��JO1GӐ�#��_Pӱ�"�O�q����@�&KE�P�IR��ܔ�@ML}R��AP�Q^�Eh08��K�SYS�q"vK�PG2�BRK�B��߄�pY�=�d�����`AD_�����B�SOC���N��D?UMMY14�p@�SV�PDE_OP��#SFSPD_O+VR-���C��ˢ&ΓOR٧3N]0ڦ�F�ڦ��OV��S!F��p���F+�r!����CC��1q"LCH�DL��RECOV(ʤc0��Wq@M����F��RO�#��Ȑ_+���� @0�e@VE}R�$OFSe@3CV/ �2WD�}�`�Z2���TR�!����E_FDO>�MB_CM���B��BL�bܒ#��adtVQR�$0p���G$�7�AM5��� eŤ��_M;��"'�<���8$CA��'�|E�8�8$HBK(1,���IO<�����QPPA������
���Ŋ����DVC_DBhC;��#"<Ѝ�Dr!S�1[ڤ�S�3[�^��ATIOq 1q�� ʡU�3���CABŐ�2�CvP��9P^��B���_� �SUB'CPU""ƐS�P  �M�)0NS�cM�"~r�$HW_C���U��S@��SA�A�pl_$UNITm�l_��AT���e�ƐCY{CLq�NECA����FLTR_2_�FIO�7(��)&B�L�Pқ/�.�_SCT�CF_`�Fb�l����|�FS(!E�e�CH�A�1��4�D°"3�RSD��$"}��#!�;_Tb�PRO������ EMi_��a�8!�a !�a���DIR0�RAIL�ACI���Mr�LO��C���Qq��#q��դ�PR=�S�A��pC/�c 	��F�UNCq�0rRIN�P�Q�0��2�!RAC �B ��[����[WARn���BL�Aq�A�����DAk�\���L�D0���Q��qeq�TI"r��K��hPRIA�!r"AF��Pz!=�;��?,`(�RK���MǀI�!ÇDF_@B�%1n�L�M�FAq@HRDiY�4_�P@RS�A��0� �MULSE�@���a �h�ưt��m�$�1[$�1$1o�~���� x*��EG00����!AR���Ӧ�09�2,%� �7�AXE��ROB���WpA��_l-��S�Y[�W!‎&S�'W�RU�/-1��@�ST�R������Eb�C 	�%��J��AB� `���&9�����OTo0� 	$��ARY��s#2��Ԓ�	ёF�I@��$LINQK|�qC1�a_�#Ұ��%kqj2XY�Z��t;rq�3�C1�j2^8'0B��'`�4����+ �3FI����7�q����'��_J�ˑ���O3�QOP_d�$;5���ATBAd�QBC��&�DUβz�&6��TURN߁�"r�E11:�p��9GFL�`_���* �@�5�*y7��Ʊ 1�� %KŐM��&8���8"r��ORQ�� a�(@#p=�j�g�#q�XU�����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb� �T{�, ��@;�uQ�� �P\�i��UuQ�We��e�SERʑe	B��E� O���UdAa s��4S�/7����AX��B�'q��E1 �e��i��irp�jJ@ �j�@�j�@�jP�j@  �j�!�f��i��i� �i��i��i�y��y�'y�7yTqHyD7EBU8�$32����qͲf2G + A!B����رnSVS�7� 
#�d��L�#� L��1W��1W�JAW��A W��AW�QW�@!E@�?D2�3LAB�2�9U4�Aӏ��C � o�ERf�5� �� $�@_ A��!�PO��à�0�#�
�_MRAt��/ d � T��ٔ�ERR����;TY&���I��V�0�cz�'TOQ�d�PL[ �d��"�� ?�w�! � pp`T)0���_V1Vr�aӔ�����2ٛ2�E����@�8H�E���$W���j��V!��$�P@��o�cI��aΣ	 �HELL_CFG�!� 5��Bo_BASq�SR3�\�� a#Sb�T��1�%��2��U3��4��5��6��e7��8���RO�����I0�0NL�\CAqB+�����ACK4� ����,��2@�&�?�7_PU�CO. U�OUG�P~ ����m�ذ�����TPհ_KcAR�l�_�RE*��P���|�QUE����uP����CST?OPI_AL7�l��k0��h��]�l0SE�M�4�(�M4�6�T�YN�SO���DI�Z�~�A�����m_T}M�MANRQ���k0E����$KEYSWITCH��ص�m���HE��BE�AT��|�E- LE(~�����U��F!Ĳ�|��B�O_HOM=�OGREFUPPR�&��y!� [�C��O��-ECOC��Ԯ0_IOCMWD
�a��v(k��� �# Dh1���UX����M�βgPgCFOR�C��� ��m�O}M.  � @�T5(�U�#P, 1�֔, 3��45��N�PX_ASt�� �0��ADD����$SIZ��$VsAR���TIP/�).��A�ҹM�ǐ ��/�1�+ U"S�U!yCz���FRIF���J�S���5Ԓ�NFp�� �� � xp`SI��TE�C���C�SGL��TQ2�@&����� ��STM�T��,�P �&BW<uP��SHOW4����SV�$��; �Q�A00�@Ma }���� �����&અ�5��6��7��8
��9��A��O ���� ��Ӂ���0��F���  G��0G���0G��@�@G��PG��1	U1	1	1+	18	U1E	2��2��2��U2��2��2��2��U2��2��2��2	U2	2	2+	28	U2E	3��3��3��U3��3��3��3��U3��3��3��3	U3	3	3+	38	U3E	4�4��4��U4��4��4��4��U4��4��4��4	U4	4	4+	48	U4E	5�5��5��U5��5��5��5��U5��5��5��5	U5	5	5+	58	U5E	6�6��6��U6��6��6��6��U6��6��6��6	U6	6	6+	68	U6E	7�7��7��U7��7��7��7��U7��7��7��7	U7	7	7+	78	�7E��VP��UP}Ds�  �`xNЦ�5�YSLOt�� � L��d���A�aTA�0d���|�ALU:ed�~�C�UѰjgF!aID_YL�ÑeHI�jI��?$FILE_���df��$2�fSA>�� hO��`E_B�LCK��b$��hD_CPUyM�yA���c�o�d��Y����Rw �Đ
PW��!� oqLA��Sp=�ts�q~tRUN� �qst�q~t���qstܼq~t �T��AC�Cs��X -$�qLEN;��tH���ph�_�I��ǀLO�W_AXI�F1�q�d2*�MZ���ă���W�Im�ւ�aR�T#OR��pg�D�Y���LACEk�ւ�p8V�ւ~�_MA2�v�8������TCV��؁��T��ي�����t��V����V�Jj�R�MDA���J��m�u�b�
���q2j�#�U�{�lt�K�JK��VK;�h��H���3��J0�����JJ��JJ��A�AL��ڐ��ڐԖ42Օ5���N1���(ʋƀW�LP�_(�g�����pr�� `�`GROUw`��}B��NFLIC���f�REQUIRE3�EBU��qB���w�2����p���q5��p�� \��APKPR��C}�Y�
ް;EN٨CLO7�驇S_M��H���u�
��qu�� ���M�C�����9�_MG��C�Co��`M�в��N�BRKL�NOL�|�N�[�R��_LI�Nђ�|�=�J����P ܔ��������������D���6ɵ�̲8k��i���q���� ��
��q)��7�PATH3�L�B�L���H�wࡠ�J�CN��CA�Ғ�ڢB�I�N�rUCV�4a��C!�UM��Y,�����aE�p����ʴ���PAYLOA��J{2L`R_AN�q�Lpp���$�M��R_F2LSHR��N�LOԡ�Rׯ�|`ׯ�ACRL_G� �ŒЛ� ��Hj`߂�$HM���FLE�Xܣ�qJ�u� :��������������1�F1 �V�j�@�R�d�v�������E����ȏڏ� ���"�4�q���6�M� ��~��U�g�y�ယ	T��o�X��H����� �藕?�����ǟِ ݕ�ԕ����%�7���JJ�� � `V�h�z���`AT��l��@�EL�� Sj��J|�Ŝ�JEy�gCTR��~�TN���FQ��HAND_�VB-���v`�� $��F2M�����ebSW�bD�'���� $$MF�:�R g�(x�,4�%��0&�A�`�=��aM)F�A(W�Z`i�Aw�A��X �X�'pi�Dw�D��P2f�G�p�)STk��!4x��!N��DY�pנ M�9$`%Ц�H��H׀c�׎���0� ��P ѵڵ��������:D�J��� ����1��R�6��QASYIMvř���v��J�8��cі�_SH>��� �Ĥ�ED����������J�İ%��C�ID�.��_VI�!X�>2PV_UNIX�FThP�J��_R�5_Rc� cTz�pT�V��@���İ��߷��U ����dD���Hqpˢ��faEN�3�DI�����O4d�`J��) x g"IJAAȱz� aabp�coc�`a�pdq��a� ��OMM�E��� �b�RqT(`PT�@� S��a7��;�Ƞ�@�h�a�iT��@<� $DU�MMY9Q�$P�S_��RFC��$v �����Pa� XƠ���SuTE���SBRY��M21_VF�8$_SV_ERF�O��\LsdsCLRJtA���Odb`O�p �� D $GL3OBj�_LO���u��q�cAp�r�@aSYS�qADR``�`�TCH  � �,��ɩb�W_NAƇ��7�Ac�T�SR���l ���
*?�&Q�0" ?�;'?�I)?�Y)��X� ��h���x������)�� Ռ�Ӷ�;��Ív�?���O�O�O�DD�XSCSRE栘p����3ST��s}y`��R��/_HA�q�� TơgpTYP �b���G�aG�蕵�Od0IS_�䓀dАUEMd�# ����ppS�qa�RSM_�q*eUNEXCEP)fW�`S_}pM�x���g�z�8����ӑCOU��S��Ԕ 1�!�UE�&��Ubwr��PRO�GM�FL@$CUgpPO�Q��5��I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp��OUS�� �� @6p�v$BU�TTp�RpR�CO�LUMq�e��SE�RV5�PANE|H�q� � �@'GEU���Fy��?)$HELPõ)B/ETERv�)ෆ� ��A � ��0`��0��0ҰIN簊�c�@N��IH�1��_� �v��LN�r� �qprձ_ò=�$H���TEXl����F�LA@��RELVB��D`��������M��?,�ű�m�����"�USRVwIEW�q� <6p�`U�`�NFI<@;�FOCU��;�7PRI@m�`�Q�Y�TRIP�qm��UN<`Md� x#@p�*eWARN)e�6�SRTOL%���g��ᴰONCOR�N��RAU����T����w�VIN�Le�� $גPA�TH9�גCACH���LOG�!�LI�MKR����v���HwOST�!�bz�R��OBOT��d�IM>� �� ����Zq�Zq;�V�CPU_AVAIYL�!�EX	�!AN���q��1r��1r���1 �ѡ�p� � #`C����@$�TOOL�$��_wJMP� ���e$SS�����VSHIF��Nc߃P�`ג�E�ȐR�����OSUR��Wk`RADILѮ��_�a��:�9a��`a�r���LULQ$OUTPUT_BM����IM�AB �@�r�TILSCO��C7����� ��&��3��A��@�q���m�I�2G��4�V�pLe�}��yD�JU��N�WA�IT֖�}��{�%�! NE�u�YBO��� �� �$`�t�SB@T;PE��NECp�Jp^FY�nB_T��R�І�a$�[Yĭc	B��dM���F� `�p�$�pb�OP?�wMAS�_DO�!QT�pD��ˑ#�%��p!"DELAY�:`7"JOY�@(� nCE$��3@ �xm��d�pY_[�!"�`�"��[���P? �4�ZABC%�� � $�"R��
�ϐ�$$CLAS>������!ϐx4�� � VIRT]ќ�/ 0ABS����1� 5� < �! F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $�6HZi{0-�AX�L�pl��!�63  ��{tIN��qztP#RE�����v�p�u�LARMRECO�V 9�rwtN�G�� .;	 �=#�
�.�0PoPLIC��?5��p�Ha�ndlingTo�ol o� 
V�7.50P/23� �!�PB���
��_SWt� U�P�!� x�F0Ȭ�t���A� v�� 864�� ��it�y� N�2 7DA�5�� j� �QB@ϐo�No�neisͅ˰ ���T�]�!L�AAxyrP_�l�V�uT��s9�U�TO�"�Њt�y��HGAPON
0g�1z��Uh�D 1581����̟ޟxry����Q 1���p�,�蘦����;�@��q_��"=�" �c�.��H���D�HTTHKYX��"�-� ?�Q���ɯۯ5���� #�A�G�Y�k�}����� ��ſ׿1�����=� C�U�g�yϋϝϯ��� ��-���	��9�?�Q� c�u߇ߙ߽߫���)� ����5�;�M�_�q� �������%���� �1�7�I�[�m���� ������!����- 3EWi{��� ���)/A Sew����/ ��/%/+/=/O/a/ s/�/�/�/�/?�/�/ ?!?'?9?K?]?o?�? �?�?�?O�?�?�?O#O]���TO�E�W��DO_CLEAN���7��CNM  � �__/_�A_S_�DSPDR3YR�O��HIc��M@�O�_�_�_�_oo +o=oOoaoso�o�o���pB��v �u���a�X�t������9�PL�UGG���G��U�P�RCvPB�@���_�orOr_7�SEGF}�K[mwxq �O�O�����?rqLAP�_�~q�[� m��������Ǐُ�����!�3�x�TOT�AL�f yx�USE+NU�p�� �H����B��RG_STR�ING 1u�
_�Mn�S5��
ȑ_ITEM1Җ  n5�� � �$�6�H�Z�l�~��� ����Ưد���� ��2�D�I/O �SIGNAL̕�Tryout �ModeӕIn�p��Simula�tedבOut���OVERR~�P = 100֒�In cycl���בProg OAbor��ב���StatusՓ	�Heartbea�tїMH Fa�ul��Aler '�W�E�W�i�{ύϟ�p�������� �C Λ�A����8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|���WOR{pΛ��(ߎ� ���� ��$�6�H�Z� l�~�������������p�� 2PƠ �X ��A{��� ����/A Sew�����SDEV[�o� #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1?�C?U?g?y?PALTݠ1��z?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_�?GRI�`ΛDQ�? _l_~_�_�_�_�_�_ �_�_o o2oDoVoho@zo�o�o�o2_l�R� �a\_�o"4FX j|����������0�B�T��oPREG�>�� f��� Ə؏���� �2�D� V�h�z�������ԟ����Z��$ARG�_��D ?	����;��  	$Z�W	[O�]O��Z��p�.�SBN_CONFIG ;�ꎱ����CII�_SAVE  �Z�����.�TCE�LLSETUP �;�%HOM�E_IOZ�Z�%�MOV_��
�R�EP�lU�(�UTOoBACKܠ���FRA:\�z� \�z�Ǡ'�`�z���ǡi�I�NI�0z���~n�MESSAG����ǡC���ODE_!D������%�O�4��n�PAUSX!�~;� ((O>� �ϞˈϾϬ������ ����*�`�N߄�r��߶�g�l TSK � wͥ�_�q�UP3DT+��d!�AſWSM_CF���;���'�-�GRgP 2:�?� N��BŰA��%�XSC�RD1�1
7� 	�ĥĢ�������� ��*�������r��� ��������7���[� &8J\n��*�>t�GROUN�UϾ�UP_NA��:�	t��_ED��17�
 �%�-BCKEDT�-�2�'K�`D���-t�z�q�Yq�z���2t1�����q�k�8(/��ED3/���/�.a/�/;/M/ED4�/t/)?�/.?8p?�/�/ED5`??��?<?.�?O�?�?ED6O�?qO�?.MO8�O'O9OED7�O`O�_�O.�O\_�O�OE�D8L_,�_�^�-�_ oo_�_ED9�_�_]o�_	-9o�oo%oCR_ �9]�oF�o�k� � N�O_DEL��GE_UNUSE���LAL_OUT� ����WD_ABORﰨ~���pITR_RTNz��|NONSk����˥CAM_�PARAM 1�;�!�
 8
S�ONY XC-5�6 234567w890 ਡ�@���?��( А\�
���{�u���^�HR5q�8̹��ŏR57ڏ��Aff��KO�WA SC310�M
�x�̆�d @<�
���e� ^��П\����*��<��`�r�g�CE__RIA_I�!�5=�F��}�z�� ��_LIU��]�����<��F�B�GP 1��Ǯ�M�_�q�0��C*  ����C1*��9��@��G����CR�C]��d��l���s��R�����[�Դm��v���������� C����b(�����=�HE�`�ONFIǰ�B�G_PRI 1�{V���ߖϨϺ�����������CHKPwAUS�� 1K� ,!uD�V�@�z� dߞ߈ߚ��߾����� �.��R�<�b��ҍO��������_�MOR�� �>��BZ?����� 	 �����*�@�N�`�������$?��q?;�;����)K��9�P���ça�-:���	�

��M���pU��ð��<��,~��D�B���튒)
m�c:cpmidb�g�f�:�  K��¥�p�|/�  �������� �sV>��pj�pkUX�?��p��pE�Ug�/���p�Uf�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����o=L���*MC��1����?43���1��t�īCz�  BHH�CPU�eB��CF��;.<C����C5rY
K�D��nyDQ��D���>��D�;D���=�F��>F�$�G}RB�7Gz�0��Y	��Y!�&w�1����s���.�p���b���BDw�M@x8�ʊ1Ҩ����g@D��p@�0EYK�EX��EQ�EJ�P F�E�F�� G��>^�F E�� FB�� H,- Ge���H3Y��:��  >�33 s���~  n8�~@��5Y�E>�ðyA��Y<#�
"Q� ���+_�'RS/MOFS�p�.8���)T1��DE ���F 
Q��;�(P  B_<_���R����	op6C4RP�Y
s@ ]AQ��2s@C�0B3�MaCR{@@*cw��UT�p�FPROG %�z�o�oigI�q���v���ldKEY_TB�L  �&S�#� ��	
�� �!"#$%&'(�)*+,-./0�1i�:;<=>?�@ABC� GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�������������������s���p`LCK�lx4�p`�`STAT ���S_AUTO_D�O���5�IND�T_ENB!���R��Q?�1�T2}�^�S�TOPb���TRL^r`LETE��Ċ�_SCREEN ��Zkcs�c��U��MMEN�U 1 �Y  <�l�oR�Y1� [���v�m���̟���� �ٟ�8��!�G��� W�i��������ïկ ��4���j�A�S��� w�����迿�ѿ��� �T�+�=�cϜ�sυ� �ϩϻ�������P� '�9߆�]�o߼ߓߥ� �������:��#�p� G�Y��������� ��$����3�l�C�U� ��y����������� ���	VY)�_MA�NUAL��t�DB;CO[�RIGڇ
��DBNUM� ���B1 e
�PXWO_RK 1!�[�_�U/4FX�_�AWAY�i�G�CP  b=�Pj_CAL� #�j�Y���܅ `�_�  1">�[ , 
�m�g�&/~&lMZ�I�dPx@P@#ONT�IMه� d��`&�
�e�MOT�NEND�o�RECORD 1(�[qg2�/{�O��! �/ky"?4?F?X?�( `?�?�/�??�?�?�? �?�?)O�?MO�?qO�O �O�OBO�O:O�O^O_ %_7_I_�Om_�O�_ _ �_�_�_�_Z_o~_3o �_Woio{o�o�_�o o �oDo�o/�oS �oL�o����@ ���+�yV,�c� u��������Ϗ>�P� ����;�&���q��� 򏧟��P�ȟ�^�� ����I�[����� � ��$�6�������j�TOLERENC�wB���L���� CS_CFG �)�/'dM�C:\U�L%04�d.CSV�� cl��/#A ��CH��z� //.ɿ��(�S�RC_OUT �*��1/V�S�GN +��"���#�09-MA�Y-20 11:�33027-JA}Np�21:48+ P;�����/.��f�pa��m��PJP�����VERSIO�N Y�V�2.0.�ƲEF�LOGIC 1,^� 	:ޠ�=�ޠL��PROG�_ENB��"p�U�LSk' ����_?WRSTJNK ���"fEMO_OPT_SL ?	��#
 	R575/#=�����0��B����TO  ��ݵϗ��V_F E�X�d�%��PA�TH AY�A�\�����5+ICTZ�Fu-�j�>#egS�,��STBF_TTS��(�	d���l#!w��� MAU��z�^"MKSWX�.�<�4,#�Y�/�
!J� 6%ZI~m��$�SBL_FAUL�(�0�9'TDIAb[�1<�<� ����123456�7890
��P ��HZl~��� ����/ /2/D/�V/h/�� P� ѩ�yƽ/��6�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�?��,/�UMP���� �ATR���1O�C@PMEl�OOY_�TEMP?�È��3F���G�|DUNI���.�YN_BRK� 2_�/�EMG?DI_STA��]���ENC2_SCR 3�K7(_:_ L_^_l&_�_�_�_�_)��C�A14_�/o@o/oAoԢ�B�T5�K�ϋo~ol�{_ �o�o�o'9K ]o������ ���#�5��/V�h� z��л`~�����ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T���x��� ������ү����� ,�>�P�b�t������� ��ο����(�f� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��:� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ���������* <N`r���� ���&8J \n�������� ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? ��?�?�?�?�?OO ,O>OPObOtO�O�O�O��O�O�O�O__NoE�TMODE 16v�5�Q �d��X
X_j_|Q�PR�ROR_PROG7 %GZ%�@��_�  �UTABLE  G[�?oo�)oRjRRSEV_?NUM  �`WP��QQY`�Q_�AUTO_ENB�  �eOS�T_N�Ona 7G[�Q�Xb  *��`�J�`��`��`d`+�`p�o�o�o�dHISUc��aOP�k_ALM �18G[ �A��l�P+�ok}������o_Nb�`  G[�a�R
�:P�TCP_VER �!GZ!�_�$E�XTLOG_RE�Qv�i\�SI�Ze�W�TOL  ��aDzr�=�#דQXT_BW�D�p��xf́t�_D�I�� 9�5��d�T�asRֆSTE�P��:P�OP_�DOv�f�PFA�CTORY_TU�NwdM�EATU�RE :�5̀�rQHand�lingTool� �� \sfm�English� Diction�ary��rodu�AA Vis��� Master�����
EN̐n�alog I/O�����g.fd̐u�to Softw�are Upda�te  F OR��matic B�ackup��H5�96,�gro�und Edit�ޒ  1 H5Camera�F��OPLGX�e�ll𜩐II) nX�ommՐshw�n��com��co����\tp���pa�ne��  opl���tyle se�lect��al �C��nJ�Ցoniwtor��RDE���tr��Reli�ab𠧒6U�Diagnos(�푥��5528�u��h�eck Safe�ty UIF��E�nhanced �Rob Serv>%�q ) "S�r�User Fr[������a��xt. oDIO �fiG�s sŢ��endx��Err�LF� p$Ȑĳr됮� �����  !��FCTN_ Menu`�v-��ݡ���TP In�ېfac�  E�R JGC�p�בk Exct�gޠ�H558��ig�h-Spex�Sk�i1�  2
P���?���mmunic'�ons��&�l��ur�ې��ST xǠ��conn���2��TXPL��n{cr�stru�����"FATK�AREL Cmd�. LE�uaG�5�45\��Run-�Ti��Env��dG
!���ؠ++��s)�S/W��[��License�Z��� 4T�0�ogBook(Syڐ�m)��H54O�M�ACROs,\�/�Offse��Lo�a�MH������r�, k�MechS�top Prot����� lic/�M=iвShif����ɒMixx��)����xSPS�Mode Switch��7 R5W�Mo�:�=.�� 74 ����g��K�2h�ul�ti-T=�M���L�N (Pos�Regiڑ�������d�ݐt Fun��ǩ�.�����Nu�m~����� lne���ᝰ Adju�p�����  - =W��tatuw᧒}T�RDMz��ot��scove
 U�9���3����uest 49�2�*�o�����62~;�SNPX b Ҟ��8 J7`���Lgibr��J�48��D�ӗ� �Ԅ�
�6O��� Parts in VCCMt�32���	�{Ѥ�J�990��/I� �2 P��TMILKIB��H���P��AccD�L�
T�E$TX�ۨ�ap�1S�Te����pkCey��wգ�d���Unexce{ptx�motnZ�0�������є��� O���� 90�J�єSP CSX�C<�f��Ҟ� P�y�We}���PRI��>vr�t�me�n�� ��iP�ɰa�����vGr{id�play�İv��0�)�H1�M�-10iA(B2�01 �2\� 0�\k/�Ascii��l�Т�ɐ/�Coyl��ԑGuar�� 
�� /P-�ޠ"�K��st{Patt ��!S�Cyc�҂�orie��I�F8�ata- qu�Ґ�� ƶ��mH5�74��RL��am����Pb�HMI �De3�(b����P�CϺ�Passw�o+!��"PE? S1p$�[���tp��� �ven��Tw�N�p��YELLOW sBOE	k$Arc��'vis��3*�n0�WeldW�cia�l�7�V#t�Opd����1y� 2F�=a�portN�(�p�T1�T� �� f��xy]�&TX��tw�igj�1� b�� ct\�JPN� ARCPSU cPR��oݲOL� wSup�2fil� p&PAɰאcro�� "PM(����O$�SS� eвtexF�� r���=�t�OssagT��P���P@�Ȱ�锱�r�tW��H'>r�dp9n��n1
t�!� z ��ascbin4psyn���+Aj�M HEL��NCL VIS� PKGS PL;OA`�MB �,��4VW�RIPE� GET_VAR� FIE 3\t���FL[�OOL:� ADD R72�9.FD \j8�'�CsQ�QE��DV�vQ�sQNO WT�WTE��}PD  �^��biRFOR ��ECTn�`���ALSE ALA�fPCPMO-130  M" #h��D: HANG �FROMmP�AQf�r��R709 D�RAM AVAILCHECKSO!���sQVPCS S�U�@LIMCHK� Q +P~dFF P�OS��F�Q R5�938-12� CHARY�0�P?ROGRA W��SAVEN`AME.�P.SV��7��$�En*��p?FU�{�T�RC|� SHAD�V0UPDAT K�CJўRSTATI��`�P MUCH �y�1��IMQ MOTN-003���}�ROBOGUI�DE DAUGHp�a���*�tou�����I� Šhd�AT�H�PepMOVET��ǔVMXPAC�K MAY AS�SERT�D��YC�LfqTA�rBE ?COR vr*Q3r�AN�pRC OP�TIONSJ1vr�̐PSH-171ZZ@x�tcǠSU1��1Hp^9R!�Q�`_TP�P��'�j�d{t�by app w�a 5I�~d�PHI����p�aTEL�MXSPD TB5b�Lu 1��UB6@�qEmNJ`CE2�61���p��s	�may 1n�0� R6{�R�} �Rtraff)��� 40*�p��f�r��sysvar scr J7��cj`DJU��bH� V��Q/�PSET� ERR`J` 6�8��PNDANT� SCREEN UNREA��'�J`MD�pPA���pR`�IO 1���PFI��pB�pGROUN�PD��G��R�P�QnRSVIP !p�a�P�DIGIT VE�RS�r}BLo�UE�Wϕ P06  �!��MAGp�ab�ZV�DI�`� S�SUE�ܰ�EP�LAN JOT` 'DEL�pݡ#Z�@=D͐CALLOb�Q� ph��R�QIP�ND��IMG�R�719��MNT/��PES �pVL�c��Hol�0Cq���t�PG:�`C�M�c�anΠ��pg.v~�S: 3D mK�view d�` L�p��ea7У�b� �of �Py���AN�NOT ACCE�SS M��Ɓ*�tn4s a��lok�^�Flex/:�Rmw!mo?�PA?��-�����`n�pa �SNBPJ AUTO-�06f����T|B��PIABLE1q� 636��PLN�: RG$�pl;pNnWFMDB�VI��>�tWIT 9x�0@o��Qui#0�ҺP�N RRS?pUS�B�� t & r/emov�@ )�_�v�&AxEPFT_=�� 7<`�pP:�O�S-144 ��h� s�g��@OST�� � CRASH� DU 9��k$P�pW� .$��_LOGIN��8&��J��6b046 i�ssue 6 J�g��: Slow� �st��c (�Hos`�c���`I�L`IMPRWtSPOT:Wh:0�T��STYW ./�VM�GR�h�T0CAT.��hos��E�q�T�� �O�S:+p�RTU' k�-S� ,����E:��pv@�2��� t\hߐ��m� ��all��0� 9 $�H� WA͐���3 CNT0 T��� WroU�al�arm���0s�d �� �0SE1���r R{�OMEBp���K�7 55��REàSE�st��g   �  �KANJI��no���INISITALIZ-p��dn1weρ<��d�r�� lx`�SC�II L�fai/ls w�� ��`�YSTEa���o��PNv� IIH���1W��Gro>Pm ol\wpSh@�P��Ϡ?n cflxL@А�WRI �OF Lhq��p?�F�up��de-rela�_d "APo SY��ch�Abetwe>:0IND t0$FgbDO���r� `��GigE�#op�erabilf  �PAbHi�H`��c�l�ead�\etfp�Ps�r�OS 0�30�&: fig��GLA )P ��i��}7Np tpswx�-B��If�g�������5aE�a EX�CE#dU�_�tPCL{OS��"rob�+NTdpFaU�c�!����PNIO V750�Q1��QaN��DB ��P M��+P�QED�DET���-� \rk��O�NLINEhSBU�GIQ ߔĠi`Z�I�B�S apABC? JARKYFq�9 ���0MIL�`� �R�pNД �p0G+AR��D*pR��PN�"! jK�0cT�P�Hl#n�a�ZE }V�� TASK�$VP2(�4`
�!�$��P�`WIBPK0�5�!FȐB/��B�USY RUNN��� "�򁐈��R�-p�LO�N�DI�VY�CUL��f3sfoaBW�p����30	V��ˠIyT`�a505.�@{OF�UNEX�P�1b�af�@�E��S�VEMG� NML�q� D0pCC_SGAFEX 0c�08"q]D �PET�`N@N�#J87����RsP��A'�M�K�`K��H GUNCH�G۔MECH�pM�c� T�  y, �g@�$ ORY L�EAKA�;�ޢS�PEm�Ja��V�tG�RIܱ�@�CTLN�TRk�FpepnR�j50�EN-`#IN�����p �`�Ǒk!��T3/dqo��STO�0A�#�L��p �0�@�Q�АY0�&�;pb1TO8pP�s���FB�@Yp`�`DU��aO�supk��t4 � P�F� Bn�f�Q�PSVGN-q1��V�SRSR)J�UP�a2�Q�#D��q l O��QBRKCTR5Ұ�|"�-�r�<pc�j!IN=VP�D ZO� ���T`h#�Q�cHset�,|D��"DUAL�� w�2*BRVO1/17 A]�TNѫt8�+bTa2473��q.?��sAUz�i�B��complete���604.� �-�`hanc�U�� F��e8�� 	 ��npJtPd!q��`���� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� xP���R(}\xPe� aʰI���E��1��p�� j  �� xSP�'^P �A�AxP�q\ 5 sig��a��"AC;a��
�b�CexPb_p��.p�c]l<bHbcb_c�irc~h<n�`tl 1�~`xP`o�dxP�b]o2�� �cb�c�ixP>�jupfrm�dxP�o�`exe�a�oFdxPtped}o��u`>�cptlibxzxP�lcr�xrxP\�b�lsazEdxP_fm �}gcxP�x���o|sp��o�mc(��ob_jDzop�u6�wf���t��wms�1q��s1ld�)��jmc�o\��n��nuhЕ��|st�e��>�pl�qp�iwcck���uvf0uxߒ��lvisn��CgaculwQ
E� F  ! Fc.sfd�Qv�� qw����Data Ac_quisi��nF�<|1�RR631`��T}R�QDMCM ��2�P75H�1�P5k83xP1��71��k59`�5�P57<P xP�Q����(���Q̖�o pxP!da�q\�oA��@��y ge/�etdms�?"DMER"؟,�GpgdD���.�m��8�-��qaq.<᡾FxPmo��h���f{��u�`13��MACR�Os, Sksaf�f�@z����03�SR��Q(��Q6��1�Q9�ӡ�R�ZSh��PxPJW643�@7ؠ6�P,�@�PRS�@���e x�Q�UС PIK�Q52 PTLC�W���xP3 (��p/O��!�Pn �xP�5��03\sfm�nmc "MNM�Cq�<��Q��\$AcX�FM���ci,Ҥ��X����cdpq+�
�s�k�SK�xP�SH560,P��,�y��refp "RE�Fp�d�A�jxP	�o�f�OFc�<gy�to�TO_����ٺ���+je�u��caxis2�xPE��\�e�q"ISDT�c��]�prax ���MN��u�b�isde܃h�\�w�xP�! isbasi5c��B� P]��QoAxes�R6��8����.�(Ba�Q�ess��xP����2�D�@�z�atis ���(�{�����~��m��FMc�u�{�<
ѩ�MNIS��ݝ ����x����ٺ���x� j75��De�vic�� Interfac�RȔQJ754��� xP�Ne`��xP�ϐ`2�б����dn� �"DNE���
t�pdnui5UI��ݝ	bd�bP>�q_rsofOb~
dv_aro��u�����stchkc��z	 �(�}onl��G!ffL+H�J(��"l"�/�n�b��z�h�amp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!�2��xpc_2pcc{hm��CHMP_�|8бpevws��2�쳌pcsF��#C� SenxPacrao�U·�-�R6�P�d�xPk�����p��g8T�L��1d M�2`���8�1c4ԡ�3 qem��GEM,\i(�>�Dgesnd�5��`�H{�}Ha�@sy����c�Isu�xD��Fmd��I��7�4���u����AccuCal �P�4� ��ɢ7ޠBU0��6+6f�6��C99\aFF q�S(�U��2�
X�p�!Bdf��cb_�SaUL��  �� ?�ܖt�o��otplus\tsrnغ�qb��Wp��t���1��T�ool (N. �A.)�[K�7�Z�(P�m����bfc�ls� k94�"Kp4p��qtpap�� "PS9H�stpswo��p�L7��t\�q����D�yt 5�4�q��w�q��� ��M�uk��rkey�����s��}t�sfoeatu6�EA��� cf)t\Xq�����̜d�h5���LR0C0�md�!�587���aR�(����2V���8c?u3l\�pa�3}H�&r-�Xu���t,�� �q "�q�Ot� �~,���{�/��1c�}����y�p�r��5� ��S�XAg�-�y���W�j874�- i�RVis���Queu�� Ƒ�-�6H�1���(����u����tӑ����
�tp�vtsn "VTCSN�3C�+�� v\p�RDV����*�pr�dq\�Q�&�vs�tk=P������n�m&_�դ�clrq8ν���get�TX��Bd���aoQϿ�0qstr�D[� ��at�p'Z����npv��@�enlIP0��`D!x�'�|���sc ����tvo/��2�q���vb����q ���!���h]��(�� Control^�PRAX�P5��g556�A@59�P[56.@56@5A��J69$@982� J552 IDVR7�hqA���16��H���La�� ���Xe�frlpa�rm.f�FRL��am��C9�@(F�����w6{���A<��QJ643�� �50�0LSE
�_pVAR $SG�SYSC��RS_?UNITS �P�2��4tA�TX.$V�NUM_OLD �5�1�xP{�50�+�"�` Funct���5tA� }��`#@��`3�a0�cڂ��9���@H5נ� �P���(�A����۶�}����ֻ}��bP�Rb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`��2�1���96����@�%C�� Aف��J�bIncr�	����\����1o5qni4�MNINp	xP�`���!��Hour�  � �2�21 ��AAVM���0y ��TUP ��J545 ���6162�V�CAM  (��CLIO ���R6�N2�MS�C "P ��STYL�C�2�8~ 13\�NRE "FHRM �SCH^�DC�SU%ORSR �{b�04 �oEIOC�1 j o542 � os| ~� egist������7�1��MASK�93�4"7 ��OCO) ��"3�8��12���� 0 HB���� 4�"39N� �Re�� �LCH=K
%OPLG%��3"%MHCR.%M�C  ; 4? ��6 6dPI�54�s� �DSW%MD� pQ�K!637�0�0p"��1�Р"4 �6~<27 CTN K V� 5 ���"7���<25�%/�T�%FRDM� �Sg!���930 FB( NB�A�P� ( HLB o Men�SM$@<jB( PVC ��s20v��2HTC�~CTMIL��~\@PAC 16U��hAJ`SAI \@EL�N��<29s�U�ECK �b�@FR3M �b�OR����IPL��Rk0CS�XC ���VVF�naTg@HTTP ��!26 ��G��@obIGUI�"%IPGS�r� H863 qb�!�07rΈ!34 �r�84 \so`! Qx`CC�3 Fb�21�!9s6 rb!51 ����!53R% 1!s(3!��~�.p"9js �VATFUJ775�"��pLR6^RP�W;SMjUCTO�@xT158 F!80���1�XY ta3!770� ��885�UO	L  GTSo
�{` �LCM �r| TS�S�EfP6 W�\@C�PE `��0VR�� l�QNL"��@001 imrb�c3 =�b�0���0�`�6 w�b-P- Ru-�b8n@5EW�b9 �Ґa� ���b�`�ׁ�b2 2000$��`3��`4*5�`A5!�c�#$�`7.%~�`8 h605? ;U0�@B6E"aRpm7� !Pr8 t��a@�tr2 iB�/�1vp3�vp5 �Ȃtr9Σ�a4@-�p�r3 F��r5`&�re`u��r7 ��r8�U�p9 \h�738�a�R2DK7"�1f��2&�y7� �3 7iCЊ�4>w5Ip�Or6�0 C�L�1bEN�4 I�pyL�uP��@LN�-PJ8�N�8Ne�N�9 H�r`�E"�b7]�|���8�В����9 2��a`0�qЂ5�%U097 0��@1�0����1 (�q�3 5R���0���mpU��0�0�7*�H@x(q�\P"RB6�q124�b;��@���f@06� x�3 p�B/x�u ��x�6 /H606�a1� ����7 6 ���<p�b155 ����}7jUU162 ��3 g��4*�6?5 2e "_��PF�4U1`���B1��z�`0'�174 �q���P�E186 R� ��P�7 ��P�8�&�3 (�90 B/�s191����@�202��6 30���A�RU2� d���2 b2h`��4Ģ᪂2�4���19�v Q�2��u2d�TRpt2� ��H�a2hPd�$�5���!U2�pD�p
�2�p��@5�0H-@��8 @�9��TX@�� �e5�`rb26Af�2^R�a�2 Kp��1y�b5Hp�`

�5�0@�gqGA��F�a52ѐ�Ḳ6�K60ہ5� ׁ2��i8�E��9�EU5@�ٰ\�q5hQ`S�2
ޖ5�p\w�۲�pJh �-P��5�p1\t�ZH�4��PCH�7j��phiw�@��P�x�~�559 ldu�  P�D���Q�@�������� �`.��P>��8��581�"�q58�!AM۲T�A iC�a589��@�x�����5 �a��12@׀0.�1���,�2��8��,�!P\h8��Lp� ��,�7��6�08�40\��ANRS 0C}A��p��{��ran��FRA ��Д�е���A% ���ѹ�Ҍ�����( ����Ќ���З��� ������ь����$�!G��1��ը���������� xS�`q�  �����`�64��M��iC/50T-H������*��)p46��� C���N����m75s�֐� Sp��b4�6��v����ГM-71?�7�З�����42������C��-��а�70�r�E��/h����O$���rD���c7c7C@�q��Ѕ���L���/��2\imm7c7�g������`���(��e����� "�������a r�L�c�T,�Ѿ�"��,�� ��x�Ex�m77t����k���a5�����)�iC��-HS-� B
_�@>���+�Т�7U��]���Mh7�s�7������-9~?�/260L_� �����Q������4��]�9pA/@���q�S�х鼔��h621��c��92������.�)92c0�g$�@ �����)$��5$����pylH"O"
�21p���t?�350� ���p��$�
��� �350!���0���9�U/0\m9��M9A3��4%� s��3M$��X%yu���"him98 J3����� i d�"m4~�103p�� ����h794̂�&R���H�0����\���g� 5AU��՜��0���*2@��00��#06�`�АՃ�է!07{r ��������kЙ @����EP�#�� ����?��#!�;&�07\;!�B1P��߀A��/ЁCBׂ2��!�:/��?�ҽCD2C5L����0�"l�2BL
#��B��\20�2_�r�re ���X��1��N����A$@��z��`C�p0U��`��04��DyA�\�`fQ����sU���\�5  ���� p�^P��<$85���+�P=�ab1l��1LT��lA8�!uDnE\(�20T��J�1 e�bH85���b����5[�16Bs��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3� � ��b�s��-`�_�Wa8�_����6I	$2�X5�1�U85��R�p6S����/�/+q��!�q��`�6o��58m[o)�m6sW��Q��?��set06�p ��3%H�5��10�p$����g/�JrH~��  ��A�856����F�� ���p/2��h�܅�✐)�5��̑v0��(��m6��Y�!H�ѝ̑m�6�Ҝ���a6�DM����-S�+��H2������ ��� �r̑��✐0��l���p1���Fx���2�\t6h T6H����Ҝ�'V l���ᜐ�V7ᜐP/����;3A7��@p~S��������4�`@圐�V���!3��2�PM[��%ܖO�7chn��vel5�p���Vq���_arp#���̑�.���2l_�hemq$�.�'�6415���5���?�� ��F�����5g�L�ј[���1��𙋹y1����M7NU�@�М��eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h����� �u���㜐��`ZS�!ܑ4���M-����S�$̑�ք �� �0��<�����07shJ�H�v�À�sF ��S*󜐳���̑�� �vl�3�A�T�#��`QȚ�Te��q�pr��,��T@75j�5�dd� ̑1�(UL�&�(�,����0�\�?���̑�a��? xSP���a��e�w�2��(�	�2�C��A/���\�+px�����21 (ܱ�CL S����B�̺��7F���?�<�lơ1L����c� ��b�u9�0����e/q���O���9�K��r9 (��,�Rs�ז�x5�G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O����1!41w���2<T@� _std��G��y� �ң�H� jdgm����w0\� �1 L���	�P�~�W*�b��t 5������%3�,���E{�������L��5\L��3�L�|#~���~!���4�#��O����h�L6A������2璥���44������[6\j4s��·���#��ol�E"w�8Pk�����?0 xj�H1�1Rr�>��6]�2a�2Aw�P ��2��|41�8��ˡ���{� �%�A<���  +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R� �ˑb�W���Fs��� �)�ѐ�!���a�1��ڛ�5��16�16�C��C����0\imBQ��d����b���\B5�-���DiL ���O�_�<ѠPEtL�E�RH�ZǠPgω�am1l��u���̑��b�<����<�$�T �̑�F����Ȋ�D�pb��X"��hr��pw� ���^P���9�0\� j971\kckrcfJ��F�s�����c��e "CTME�r��������a�`main.p[��g�`run}�_vc�#0�w�1O�ܕ_u����bctm�e��Ӧ�`ܑ�j7�35�- KAREL Use {�	U���J��1��
�p� Ȗ�9�B@���L�9��7j[�a�tk208 "KP��Kя��\��9���a��̹����cKRiC�a�o ��kc�q J�&s�����Grſ� fsD��:y��s�ˑ1X3\j|хrdtB�,� ��`.v�q�� ��sǑIf�Wfj52��TKQuto S�et��J� H5nK536(�932�Z��91�58(�9�BA�1(�74O,A$�?(TCP Ak��В/�)Y� �\t�pqtool.v��v���! co�nre;a#�Control Re��ble��CNRE (�T�<�4�2���D�)����S�552��q(g�� (򭂯4X�cO�ux�\sfuts�UTS`�i�栜����t�棂��? 68�T�!�SA OO+D6���������,!��6c+� ig.t�t6i��I0�TW8 ���la��vo58�o�bFå򬡯i�Xh��!Xk�0Y!�8\m6e�!6EC���v��6���������<16�A���A�6s����U�g�TX|ώ���r1�qR��˔Z4�T�����,#�eZp)g����<O NO0���uJ��tCR;�x�F�a� xSP�f���prdsuchk �1��2&&?���	t��*D%$�r(��@���娟:r��'�s�q8O��<scrc�C�<\At�trldJ"�o�\�V����Pa�ylo�nfir1m�l�!�87��7� �A�3ad�! ��?ވI�?plQ��3���3"�q��x p�l�`���d7��l�calC�uDu���;���mov�����i'nitX�:s8O�p�a�r4 ��r67A4�|�e GenerGatiڲ���7g2�q$��g R� (#Sh��c ,|�bE��$Ԓ\�:�"��4��4�4�. sg��5�F$d6�"e;Qp "SH�AP�TQ ngcr pGC�a(�&"<� ��"GDA¶��r6�"aW�/�$�dataX:s�"t�pad��[q�%tput;a__O7;a�o8(�1�yl+s�r�?�:H�#�?�5x�?�:c O��:y O�:�IO�s`O%g�qǒ�?�@08\��"o�j92;!�P�pl.Colli=s�QSkip#��@ 5��@J��D��@\ވP�C@X�7��7��|s2��ptclsF�LS�DU�k?�\_ ets�`�< \�Q��@���`dc�KqQ�FC;��J,�n��` (��4eN����T�{��� 'j(�c�����/IӸaxȁ��̠H������зa�e\mc�clmt "CL�M�/��� mate�\��lmpALM0�?>p7qmc?����2vm�q��%�3s���_sv90�_x_m#su�2L^v_� K�o�{in�8(3r<�c_logr�N�rtrcW� �v_3�~yc��d��<�te��derv$cCe� Fiρ�R��Q�?�l�enter߄|��d(Sd��1�TX�+�fK�r�a99sQ9x+�5�r\tq\�� "FNDR����STDn$�LANG�Pgui��D⠓�S����Ơ�sp�!ğ֙uf �ҝ�s����$�����e+�=����������ࠓ���w�H�r\f�n_�ϣ��$`x�tc�pma��- TC�P�����R638� R�Ҡ��38
��M7p,���Ӡ�$Ӏ��8p0Р�VS,�>�tk��99�a��B3�� �PզԠ��D�2�����UI��t���hqB���8��������p���rqe�ȿ��exe@ 4φ�B���e38�ԡG��rmpWXφ�var@�φ�3N������vx�!ҡ��q��RBT $cO�PTN ask �E0��1�R MA�S0�H593/�9�6 H50�i�48
0�5�H0��m�Q�QK��7�0�g�Pl��h0ԧ�2�ORD�P��@"��t\mas��0�a��"�ԧ�����k�գR�����¹`m��b��7�.f���u�d��r��splayD�E���1>w�UPDT Ub���887 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q `�䗣�#��К�`2�� vlv��Ù�`$�>�b���! S���Easy/К�U�til��룙�51G1 J�����R7 Θ�Nor֠��inGc),<6Q�� �`�c��"4�[���98Q6FVRx So����q�nd6����P�� 4�a\ (��
  ����D���d��K�bdZ����men7���- Me`tyFњ�Fb¨0�TUa�57	7?i3R��\��5�u?��!� n����f������l\mh�Ц�űE|Ghmn�	��<\HO���e�1�� l!D��y��Ù�\|�p����B���Ћmh�@��:.aG! ���/�t�55�6�!X�l�.us��Y/k)�ensubL���eK�h�� �B\1;5�g?y?�?�?D��?*r�m�p�?Ktbox  O2K|?�G��C?A%�ds���?1ӛ#�  �TR��/��P�4B�`��U�P�V�P"�Q�P0@�U�PO��P�"�T3�U@�P�f�Pk"�2}�4�T@�P�f�P2�"�Q5�S��Q���R?Ă�Q3t.��P׀al��P+O�P517��IN�0a��Q(}g��PESTf3ua�PB�l��ig�h�6�aq��P? � xS��`�  n�0mbum�pP�Q969g�6!9�Qq��P0�baAp|�@Q� BOX��,>vche�s�>v�etu㒣=wffse�3���]�;u0`aW��:zol�sm�<ub�a-��]D�K�ibQ�c����Q<twaǂ� tp�Q҄Tar�or Recov�b�O�P�642 ����a�q��a⁠Q3Erǃ�Qry�з`�P'�T�`�aar�������	{'�pak971��71��m���>�pjot��PXc���C�1�adb -�ail��nag���b�QR629�a�Q��b��P  �
�  �P��$$C�L[q ���t������$�PS_DIGIT�.��"�!� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv��������*璬1:PRODUCT�Q0\PGSTK�bqV,n�99��\���$FE�AT_INDEX���~��� 搠ILECO_MP ;��)���"��SETU�P2 <�~��  N !��_AP2BCK� 1=�  #�)}6/E+%,/i/��W/�/~+/�/ O/�/s/�/?�/>?�/ b?t??�?'?�?�?]? �?�?O(O�?LO�?pO �?}O�O5O�OYO�O _ �O$_�OH_Z_�O~__ �_�_C_�_g_�_�_	o 2o�_Vo�_zo�oo�o ?o�o�ouo
�o.@ �od�o���M �q���<��`� r����%���̏[��� ����!�J�ُn��� ����3�ȟW������ "���F�X��|���� /���֯e������0� ��T��x������=� ҿ�s�ϗ�,ϻ�9��b�� P/ 2>) *.VRiϳ�!�*�������ߌ��PC�7�!�OFR6:"�c������T��߽�Lը���ܮx���*.F��>� �	N�,�k���ߏ��STM @�����Qа���!��iPendant Panel���H��F���4�������GIF��������u����JPG &P��<�����	PANEL1.DT��������2�Y�G��
3w�� ���//�
4�a/��O///�/�
T�PEINS.XM)L�/���\�/�/��!Custom Toolbar?��PASSWO�RD/�FRS�:\R?? %P�assword ?Config�?� �?k?�?OH�6O�?ZO lO�?�OO�O�OUO�O yO_�O�OD_�Oh_�O a_�_-_�_Q_�_�_�_ o�_@oRo�_voo�o )o;o�o_o�o�o�o* �oN�or��7 ��m��&��� \�����y���E�ڏ i������4�ÏX�j� �������A�S��w� ����B�џf����� ��+���O������� ��>�ͯ߯t����'� ��ο]�򿁿�(Ϸ� L�ۿpς�Ϧ�5��� Y�k� ߏ�$߳��Z� ��~�ߢߴ�C���g� ����2���V����� ����?����u�
� ��.�@���d������ )���M���q����� <��5r�%� �[�&�J �n��3�W ���"/�F/X/� |//�/�/A/�/e/�/ �/�/0?�/T?�/M?�? ?�?=?�?�?s?O�? ,O>O�?bO�?�OO'O �OKO�OoO�O_�O:_ �O^_p_�O�_#_�_�_ Y_�_}_o�_�_Ho)f��$FILE_D�GBCK 1=���5`��� ( �)
�SUMMARY.�DGRo�\MD:�o�o
`Dia�g Summar�y�o�Z
CONSLOG�o�o�a
J��aConsol�e logK�[��`MEMCHEC�K@'�o�^qM�emory Da�ta��W�)}�qHADOW���P��sSha�dow Chan�gesS�-c-�?�)	FTP=���9����w`qmme?nt TBD׏�W�0<�)ETHERNET̏�^�q��Z��aEthe�rnet bpfi�guration�[��P��DCSVR�Fˏ��Ïܟ�q%��� verif�y allߟ-c1�PY���DIFF�ԟ��̟a��p%��diffc���q¡�1X�?�Q�� �����X��CHGD��¯ԯi��p!x��� ���2`�G�Y�� ��� ��GD��ʿܿq��p8���Ϥ�FY3h�O�a��� ��(σGD������y��p��ϡ�0�UPDA�TES.�Ц��[�FRS:\������aUpdates� List���kP�SRBWLD.C	M.��\��B��_p�PS_ROBOWEL���_����o�� ,o!�3���W���{�
� t���@���d����� /��Se���� �N�r� = �a�r�&�J ���/�9/K/� o/��/"/�/�/X/�/ |/�/#?�/G?�/k?}? ?�?0?�?�?f?�?�? O�?OUO�?yOO�O �O>O�ObO�O	_�O-_ �OQ_c_�O�__�_:_ �_�_p_o�_o;o�_ _o�_�o�o$o�oHo�o �o~o�o7�o0m �o� ��V�z �!��E��i�{�
� ��.�ÏR�������� ��.�S��w������ <�џ`������+��� O�ޟH������8����߯n����$FI�LE_��PR����������� �MDON�LY 1=4�� 
 ���w�į ��诨�ѿ������� +Ϻ�O�޿sυ�ϩ� 8�����n�ߒ�'߶� 4�]��ρ�ߥ߷�F� ��j�����5���Y� k��ߏ���B����� x����1�C���g��� ����,���P����������?��Lu�VISBCKR�<�a�*.VD|�4 �FR:\���4 Vision� VD file � :LbpZ� #��Y�}/$/ �H/�l/�/�/1/ �/�/�/�/�/ ?�/1? V?�/z?	?�?�???�? c?�?�?�?.O�?ROdO O�OO�O;O�O�OqO _�O*_<_�O`_�O�_�_%_�_�MR_G�RP 1>4��L�UC4  B��P	 ]�ol`��*u����RHB ��2� ��� ��� ���He�Y�Q`o rkbIh�oJd�o�Sc��o�oK�uL��)�J��F��5U�aSm�|��o�o E����Eà�E����.5�9q��l>���}@��bA�qTlq?eݐA�l�xq�0~�� F@ �r�d�a}J��N�Jk�H9��Hu��F!��/IP�s}?�`��.9�<9���896C'�6<,6\b��}B��B���C{��B���>B�B��� �"7�A����B��A���VA�SA��#���, A�PA�����|�ݏx����%���p�A6Β@U��{ �v�a�������П�� ��ߟ��<�'�hz;BH�P �a`�Q��QAK�@������ǯ�P
6�PJ��P�\�˯�o�o�B��P5���@�3�3@���4�m�T�U�UU��U�~w�>u?.�?!x�^���ֿ���3��=[�z�=�̽=�V6<�=�=��=$q��~���@8�i7G���8�D�8?@9!�7ϥ��@Ϣ���cD�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p������������� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__/  D�UPE_�Hly_�\@@m_B�=��vR/��I�O�SMT*�G���
�o�o+l�$HOST�C�1H�I� Ĺ�zMSM��l[bo�	1�27.0�`1�o  e�o�o�o #z�oFXj|�l6�0s	anonymous�����F�)Bao�&�&��o�x��o������ ҏ�3��,�>�a� O����������Ο�U %�7�I��]����f� x��������ү��� �+�i�{�P�b�t��� ���������S� (�:�L�^ϭ�oϔϦ� �������=��$�6� H�Zߩ���Ϳs����� ������ �2���V� h�z��߰������� ��
��k�}ߏߡߣ� ���߬���������C� *<Nq�_�� ����-�?�Q�c� eJ��n���� ���/"/E� X/j/|/�/�/� %'/?[0?B?T?f? x?��?�?�?�?�?? E/W/,O>OPObO�KDa�ENT 1I�K� P!�?�O  �P�O�O�O�O�O#_ �OG_
_S_._|_�_d_ �_�_�_�_o�_1o�_ ogo*o�oNo�oro�o �o�o	�o-�oQ u8n����� ���#��L�q�4� ��X���|�ݏ���ď�֏7���[���B�?QUICC0��h�z�۟��1ܟ��ʟ+��2,���{�!?ROUTER|�X��j�˯!PCJO�G̯��!19�2.168.0.�10��}GNAME� !�J!RO�BOT�vNS_C�FG 1H�I ��Aut�o-starte�d�$FTP�/ ���/�?޿#?��&� 8�JϏ?nπϒϤ�ǿ ��[������"�4�G�#������������ �����������&�8� J�\�n������� ������/�/�/F��� j��ߎ����������� ��0S�T��x �����!�3�� G,{�Pbt�� C����/� :/L/^/p/�/��� 	/�/=?$?6?H? Z?)/~?�?�?�?�/�? k?�?O O2ODO�/�/ �/�/�?�O�/�O�O�O 
__�?@_R_d_v_�_ �O-_�_�_�_�_oUO gOyO�O�_ro�O�o�o �o�o�o�_&8 Jmo�o����� o)o;oMoO!��oX� j�|�����oď֏� ���/���B�T�f�x����^�ST_ERR� J;�����PDUSIZ  ���^P����>ٕW�RD ?z����  guest���+�=�O��a�s�*�SCDMN�GRP 2Kz�;Ð��۠�\��K�� 	P01.14 8�q�   y���B    �;����{ ����������������������~ �ǟI��4�m�X�|�� � i  � � 
���� �����+��������
���l�.Vx����"�l�ڲ۰s�d��������_GROU��L.�� ��	��۠�07K�QUPD � ���PČ�T�Yg�����TT�P_AUTH 1�M�� <!i?Pendan����<�_�!KAREL:*����݇KC%�5�G���VISION SCETZ���|��� �ߪ���������
�W�.�@��d�v���C?TRL N��������
�FF�F9E3���F�RS:DEFAU�LT�FAN�UC Web S_erver�
�� ����q��������������WR_CON�FIG O�� ����IDL_�CPU_PC"���B��= �BH�#MIN.�BGNR_IO��� ����% NPT_SI�M_DOs}T�PMODNTOL�s �_PRTY��=!OLNK 1P���'�9K]o�MAS�TEr �����O_gCFG��UO��|��CYCLE����_ASG 19Q���
 q2/ D/V/h/z/�/�/�/�/��/�/�/
??y"N�UM���Q�I�PCH��£RTRY_CN"�u���SCRN������� ���R���?��$J2�3_DSP_EN������0OBP�ROC�3��JO�GV�1S_�@��8�?�';ZO'?}?0CPOSREO~�KANJI_� Ϡu�A#��3T ����E�O�ECL_L�M B2e?�@EYLO�GGIN��������LANGUA�GE _�=�� }Q��LG�2U������ �x������PC � �'0������MC�:\RSCH\0�0\˝LN_DISP V��������TOC�4D�z\=#�Q�?PB?OOK W+��`o���o�o���Xi��o�o�o�o�o~}	x(y��	ne�i��ekElG_BUF/F 1X���}2����Ӣ��� ���'�T�K�]��� ��������ɏۏ����#�P��ËqDCS� Zxm =���%|d1h`���ʟܟ|�g�IO 1[+G �?'����'� 7�I�[�o�������� ǯٯ����!�3�G� W�i�{�������ÿ׿z�El TM  ��d��#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝߜ�t�SEV�0m.�TYP�� �0�$�}�ARS"�(_|�s�2FL 1\��0���������0�����5�TP<P����DmNGNA�M�4�U�f�UPSF`GI�5�A�5s��_LOAD@G �%j%@_M�OV�u����MAXUALRMB7�P8 ��y���3�0]&q
��Ca]s�3�~��� 8@=@^+ �Z�v	��V0+�P1�A5d�r���U����� �E(iTy� ������/ / A/,/Q/w/b/�/~/�/ �/�/�/�/??)?O? :?s?V?�?�?�?�?�? �?�?O'OOKO.OoO ZOlO�O�O�O�O�O�O �O#__G_2_D_}_`_ �_�_�_�_�_�_�_o 
ooUo8oyodo�o�o �o�o�o�o�o�o-���D_LDXDIS�A^�� �MEMO�_APX�E ?��
 �0y� ���������ISC 1_�� �O����W�i� ����Ə�����}� �ߏD�/�h�z�a��� ����������� @���O�a�5������� �����u��ׯ<�'� `�r�Y������y�޿ �ۿ���8Ϲ�G�Y� -ϒ�}϶ϝ�����mπ����4��X�j�#�_MSTR `��~}�SCD 1as}�R���N�������� 8�#�5�n�Y��}�� �����������4�� X�C�|�g��������� ������	B-R xc������ �>)bM� q�����/� (//L/7/p/[/m/�/ �/�/�/�/�/?�/"? H?3?l?W?�?{?�?�?��?n�MKCFG �b���?��LT�ARM_�2cRu;B �3Wp|TNBpMETPUOp��2����NDS?P_CMNTnE@8F�E�� d���N��2A�O�D�EPO�SCF�G�NPS�TOL 1e-�4=@�<#�
;Q�1 ;UK_YW7_Y_[_m_�_ �_�_�_�_�_o�_o Qo3oEo�oio{o�o�a��ASING_CH�K  �MAqODAQ2CfO�7J�e�DEV 	Rz	�MC:'|HSI�ZEn@����eTA�SK %<z%$�12345678�9 ��u�gTRI�G 1g�� l<u%���3����>svvYPaq��kE�M_INF 1h�9G `�)AT&FV0�E0(���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ���ڄH�� ����G�ֈAO�w� 2�������џ ���� ����͏ߏP��t��� ����]�ί����� (�۟�^��#�5��� ��k�ܿ� ϻ�ů6� �Z�A�~ϐ�C���g� y��������2�i�C� h�ό�G߰��ߩ��� �ϫ��������d�v� )ߚ��߾�y����� ���<�N��r�%�7� I�[������9�& ��J[�g��>�ONITOR�@G� ?;{   	?EXEC1�3�U2�3�4�5�T�p�7�8�9�3�n�R�R�R RRR(R@4R@RLR2YU2e2q2}2�U2�2�2�2�U2�3Y3e3���aR_GRP_SOV 1it��q(�5�
��5��m۵MO~q_DC�d~�1PL_NAM�E !<u� ��!Defaul�t Person�ality (f�rom FD) ��4RR2k! 1j�)TEX)TH��!�AX d�?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO�O�O�Ox2-?�O�O �O__0_B_T_f_x_�b<�O�_�_�_�_�_ �_o o2oDoVoho&x�Rj" 1o�)&0=\�b, �9��b��a @D�  &�a?��c�a?�`�a�aA'�6�ew�;�	l�b	 ��xJ�p��`�`	p �< �(p�� �.r� K��K ��K=*��J���J���JV��kq`q�P��x�|� @j��@T;f�r�f��q�acrs�I5�� ��p���p�r��ph}�3��´7  ��>��p�h�`z��Ꝝ�"�Jm�q� H�N��ac��$�dw���  �  �P� Q� �� |  а�m�Əi}	'� � ��I� �  �����:�È~�È=���(��#�a	���I  ?�n @H�i~�ab�Ӌ�b�$w���"N0��  '�Ж�q�p@2��@Ǔ���r�q5�C��pC0C�@ C�����`
��A1q  � @B�V~X�
nwB0h�A��p�ӊa�p�`���aDz����֏���Я	�pv��( �� -��I��-�=��A&�a�we_q�`�p� �?�ff ���m��� �����Ƽ�!@ݿ�>N1�  P�apv(�` ţ� �=�qst��/?���`x`�� �<
6b<߈�;܍�<�ê�<� <�&P�ό�AO��c1��ƾ��?fff?O�?y&��qt@�.���J<?�`�� wi4����dly�e߾g ;ߪ�t��p�[ߔ�� �ߣ����� ����6�wh�F0%�r�!�߷�1ى����E��� E�O�G+� F�!���/���?�e�P���t���lyBL�cB��Enw4��� ����+��R��s���������h�Ô�>��I�mXj�F��A�y�weC�p�������#/�*/c/N/wi�����fv/C�`� CHs/�`
=$�p�<!�!������'�3A�A��AR1AO�^?�$�?����±
=ç>�����3�W
�=�#�]�;e��׬a@����{�����<��>(�B�u���=B0��?����	R��z�H�F�G����G��H�U`�E���C�+���}I#�I���HD�F���E��RC�j�=�>
I���@H�!H�(� E<YD0 w/O*OONO9OrO]O �O�O�O�O�O�O�O_ �O8_#_\_G_�_�_}_ �_�_�_�_�_�_"oo oXoCo|ogo�o�o�o �o�o�o�o	B- fQ�u���� ���,��P�b�M� ��q�����Ώ���ݏ �(��L�7�p�[��� ���ʟ���ٟ����6�!�Z�E�W���#1(� ��9�K���<ĥ �����Ư!3�8���!�4Mgs��,�I�B+8�J��a���{�d�d������ȿ���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ��ϰ�������  %��  ��h�Vߌ�z߰�&ڀg�/9�$������� 7����A�S�e�w�  ��������������2 F��$�&Gb��������!C���@����8�����F�� DzN�� F?�P D�������)#B�'9K]�o#?���@@*v
4$8�8��u8�.
 v ���!3EW i{����:�� ��ۨ�1���$MSKCFM�AP  ��� ����(.�ONREL  �!9��EXCFENBE'q
#7%^!FNCe/�W$JOGOVLI�ME'dO S"d�K�EYE'�%�R�UN�,�%�S?FSPDTY0g&<P%9#SIGNE/W$�T1MOT�/T!��_CE_GRP� 1p��#\ x��?p��?�?�?�? �?O�?OBO�?fOO [O�OSO�O�O�O�O�O _,_�OP__I_�_=_ �_�_�_�_�_oo�_�:o�TCOM_�CFG 1q	-оvo�o�o
Va_A�RC_b"�p)U?AP_CPL�ot$�NOCHECK {?	+ � x�%7I[m ���������!�.+NO_WAI�T_L 7%S2NT�^ar	+�s�_7ERR_12s	)9�� ,ȍޏ��x����&��dT_M�O��t��, ���*oq�9�PARAuM��u	+��`a�ß'g{�� =?��345678901��,��K�]�9� i�������ɯۯ��&g������C��cU�M_RSPACE�/�|����$OD�RDSP�c#6p(O�FFSET_CAsRT�o��DISƿ���PEN_FIL�E尨!�ai��`OPTION_IO�/���PWORK 5ve7s# ��Vŀؤ��p�4�p�	C ���p��<����RG_DSBL  ��P#��ϸ�RIENTTOD �?�C�� !=#���UT_SIM�_D$�"���V~��LCT w}��h�iĜa[�1�_PEsXE�j�RATv�Ш&p%� ��2^3j)TEX)TH�)�X d3����� ��%�7�I�[�m�� �������������!�3�E���2��u��� ������������c�<d�ASew� ��������썒^0OUa0o(ҿ�(����>u2, ���O ~H @D�  [?�aG?��cc��D][�Z�;��	ls��xoJ���������< ���� ��2�H�(��H3k7H�SM5G�22G���Gp
͜��'f�/-,2�C%R�>�D!�M#{|Z/��3�����4y H "�c/u/��/0B_���{�jc��t�!�/ �/�"t32�����/6  ���P%�Q%��%�|�T��S62�q?'e	'�� � �2I�� �  �=�+==��ͳ?�;�	�h	�0�I  ?�n @�2�.��Ov;��ٟ?&gN [OaA''�uD@!:� Cb@C�@F#H!��/�O�O sb
��Ab@�@�@�H�@�e`0Bb@QA�0Yv: �13Uwz$oV_�/z_e_�_�_�	��( �� -�2�1�1ta��Ua�c���:A-����.  �?�ff ���[o"o�_U�`oDXÜQ8���o�j>�1'  Po�V(���e�F0�f�Y���L�?�����xb�P<�
6b<߈;�܍�<�ê<� <�&�,/aA�;r�@Ov0P�?fff?�0?&�ip�T@�.{r�?J<?�`�u#	 �Bdqt�Yc�a� Mw�Bo��7�"�[� F��j�������ُ� ���3����,����(�E�� E�~�3G+� F��a ��ҟ�����,��PP�;���B�pAZ� >��B��6�<OίD��� P��t�=���a�s���<��6j�h��7o��>�S��O��0���Fϑ�A�a�_���C3Ϙ�/�%?��?���������#	�Ę��P �N||CH���Ŀ�������@I�_�'�3�A�A�AR1�AO�^?�$��?��� �±
�=ç>�����3�W
=�#�\ U��e���B��@���{����<����(�B��u��=B�0�������	�b�H�F�G����G��H��U`E���C��+��I#��I��HD��F��E��R�C�j=[�
�I��@H�!�H�( E<YD0߻������ ��� �9�$�]�H�Z� ��~������������� #5 YD}h� ������
 C.gR���� ���	/�-//*/ c/N/�/r/�/�/�/�/ �/?�/)??M?8?q? \?�?�?�?�?�?�?�? O�?7O"O[OmOXO�O |O�O�O�O�O�O�O�Ot3_Q(�������b��gUU���W_i_2�3�8�x�_�_2�4Mgs�_��_�RIB+�_�_�a���{�m iGo5okoYo�o}l��%P'rP�nܡݯ�o�=_�o�_�[R�?Q�u���  �p���o��/� �S��z
uүܠ�������ڱ�������8����  /�M��w�e��������l2 �F�$��Gb���t��a�`�p�S�C�y�@p�5�G�Y�۠�F� Dz��� F�P D�!�]����پ��ʯ�ܯ� ��~�?��W�@@�?�K��K���K���
 �|�������Ŀ ֿ�����0�B�TϸfϽ�V� ���{���1��$PAR�AM_MENU �?3���  DE�FPULSEr��	WAITTMO{UT��RCV��� SHELL�_WRK.$CU�R_STYL���	�OPT��P�TB4�.�C�R_DECSN���e�� ߑߣ���������� �!�3�\�W�i�{�����USE_PRO/G %��%����.��CCR���e�����_HOST �!��!��:���T �`�V��/�X��>��_TIME��^���  ��GDE�BUG\�˴�GI�NP_FLMSKĻ���Tfp����PG�A  ����)CyH����TYPE��������� �� -?hc u������� //@/;/M/_/�/�/ �/�/�/�/�/�/??�%?7?`?��WORD� ?	=	R}Sfu	PNSU�Ԝ2JOK�DR�TEy�]TRACECTL 1x3���� �`/ 	&�`�`�>��6DT Qy3��%@�0D � � `2@,�6D-6D.6D/6D026D16A�c2@�` 8BV�8BR�8BM 8BJ��8BF�8B6D6D	�6D
6D6D6D�6D6D6D^�8B�6D6D6D6D(6D�8B6D6D~P�8B6DV�8Bj�8B�6D6DҀ8B�8B!�6D"6D#6D�8B%�6D&6D'6D(6D)6D*6D5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m� �������Ǐن.A� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� �r����� ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ����������� �*��$PG�TRACELEN�  )�  �_�(��>��_UP z����m�u�Y��n�>�_CFG M{m�W�(�n����PКӂ�DEF�SPD |��l�aP��>�IN�пTRL }���(�8����PE_C�ONFI��~m�O�mњ��ծ��LID����~=�GRP 1���W��)�A ����&ff(�A+�33D�� D]�� CÀ A@1��Ѭ(�d�Ԭ���0�0�� 	 �1�ح֚��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P; t_�������  Dz (�
H�X~i� �����/�/�D///h/S/�/��
�V7.10bet�a1��  �A�E�"ӻ��A (�� ?!G�^�!>���"�����!���!BQ��!A\� �!���!*2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?O O:O%O7OpO[O�OO �O�O�O�O�O_�O6_ !_Z_E_~_i_�_�_�_ �_�_�_'o2o�_Vo AoSo�owo�o�o�o�o �o�o.R=vx1�/�#F@ �y �}��{m��y=�� 1�'�O�a��?�?�?�� ����ߏʏ��'�� K�6�H���l�����ɟ ���؟�#��G�2� k�V���z�������� o��ίC�.�g�R� d����������п	� ��-�?�*�cώ�� �Ϯ������B� ;�f�x�������DϹ� �߶��������7�"� [�F�X��|����� ������!�3��W�B� {�f��������� ��� ��/S>wb t������ =OzόϾψ� ���ϼ� /.�'/R� d�v߈߁/0�/�/�/ �/�/�/�/#??G?2? k?V?h?�?�?�?�?�? �?O�?1OCO.OgORO �OvO�O�O���O�O�O __?_*_c_N_�_r_ �_�_�_�_�_o�_)o Tfx�to��� /�o/>/P/b/ t/mo�|��� ����3��W�B� {�f�x�����Տ���� ���A�S�>�w�b� ���O��џ������ +��O�:�s�^����� ��ͯ���ܯ�@oRo do�o`��o�o�o��ƿ �o���*<N�Y� �}�hϡό��ϰ��� �����
�C�.�g�R� ��v߈��߬�����	� ��-��Q�c�N�ﲟ ���l�������� ;�&�_�J���n����� ������,�>�P�: L���������� ��(�:�3��0i T�x����� /�///S/>/w/b/ �/�/�/�/�/�/�/? ?=?(?a?s?��?�? X?�?�?�?�?O'OO KO6OoOZO�O~O�O�O �O�O*\&_8_r����_�_��$P�LID_KNOW�_M  ��� Q�TSV� ���P��?o"o4o �OXoCoUo�o R�S�M_GRP 1�T�Z'0{`�@�`)uf�e�`
�5�  �gpk'P e]o�����`�����SMR�cŅ�mT�EyQ}?  yR����������폯� ��ӏ�G�!��-��� ��������韫���ϟ �C���)������������寧���QST^�a1 1��)����P0� A  4��E2�D�V�h����� ��߿¿Կ���9�� .�o�R�d�vψ��Ϭ�(�����2�0� Q'�<3��3�/�A�S��4l�~ߐߢ߂�5���������6 
��.�@��7Y�k�}���8�������~�MAD  �)��PARN_UM  !�}o\+��SCHE� S��
��f���S��UP�Df�x��_CMP_�`H�� ��'�UER_C;HK-���ZE�*<RSr��_�Q_#MOG���_�X��_RES_G�� !���D�>1b U�y�����@/�	/���� +/�k�H/g/l/��� �/�/�/�	��/�/�/ �X�?$?)?���D? c?h?����?�?�?��V 1��U�ax�@�c]�@t@(@�c\�@�@D@�c[�*@��THR_INRr�J�bz�Ud2FMASS?O� ZSGMN>OqCM�ON_QUEUE� ��U�V P~P UX�N$ UhN�FV�@END�A��I�EXE�O�E��BE��@�O�COPTIO��G��@PROGR�AM %�J%��@�?���BTASK�_IG�6^OCFG� ��Oz��_�PD�ATA�c��[@Ц2=�DoVohozo �j2o�o�o�o�o�o�);M jINFO[��m��D� �������1� C�U�g�y���������@ӏ���	�dwpt�l� )�QE DIT� ��_i��^WE�RFLX	C�RG�ADJ �tZA	�����?נʕFA��?IORITY�GW}���MPDSPNQ�����U�GD��O�TOE@1�X�� (!AF:@E�� c�Ч!tc�pn���!ud|����!icm����?<�XY_�Q��X���Q)� *0�1�5��P��]� @�L���p�������� ʿ��+�=�$�a�H��ϗ�*��PORTT)QH��P�E���_CARTREP�PX��SKSTA��H�
SSAV�@��tZ	2500H863���_x�
�'�U�X�@�swP�tS�ߕߧ���URGeE�@B��x	WF��#DO�F"[W\��������WRUP_DELAY �X�>��R_HOTqX	B�%�c���R_NORMALq^R��v�SEMI�����9�_QSKIP'��tU;r�x 	7�1� 1��X�j�|�?�tU�� ������������ $J\n4��� �����4F X|j���� ���/0/B//R/�x/f/�/�/�/tU�$�RCVTM$��D]�� DCR'����Ў!C`N�C��d�C��o?���>��L<�|�{:��g�&���/���%��t����|���}'�:�o?�� �<
6b<���;܍�>u.��?!<�&�?h?�?�?�@>��? O O2ODOVOhOzO�O �O�O�O�O�?�O�O_ _@_+_=_v_Y_�_�_ �?�_�_�_oo*o<o No`oro�o�o�o�_�o �o�o�o�o8J- n��_����� ��"�4�F�X�j�U ������ď���ӏ� ��B�T��x����� ����ҟ�����,� >�)�b�M��������� ���ïկ�Y�:�L� ^�p���������ʿܿ � ����6�!�Z�E� ~ϐ�{ϴϗ�����-� � �2�D�V�h�zߌ� �߰���������
��� .��R�=�v��k�� ���������*�<� N�`�r���������� ������&J\ ?������� �"4FXj|���!GN_ATC� 1�	; �AT&FV0E�0�ATDP�/6/9/2/9��ATA�,�AT%G1%�B960�+�++�,�H/,��!IO_TYPE'  �%�#t��REFPOS1 �1�V+ x�u/�n�/j�/
= �/�/�/Q?<?u??�?�4?�?X?�?�?�+2 1�V+�/�?�?\O��?�O�?�!3 1� O*O<OvO�O�O_�OS4 1��O�O�O�_�_t_�_+_S5 1�B_T_f_�_o	o|Bo�_S6 1��_��_�_5o�o�o�oUoS7 1�lo~o�o�o�H3l�oS8 1�%_����SMASK 1�V/  
?�M��'XNOS/�r�������!MOTE  �n��$��_CFG �����q���"PL_RANG������POWER �����SM_D�RYPRG %�o�%�P��TAR�T ��^�UME_PRO-�?�����$_EXEC_E�NB  ���GSPD��Րݘ��gTDB��
�RM�.
�MT_'�T�����OBOT_N�AME o�����OB_ORD_NUM ?��b!H863  �կ�����PC_TI�MEOUT�� xޚS232Ă1��� LTE�ACH PENDcAN��w��-���Maint�enance CGons���s�"��~�KCL/Cm�Ț

���t�ҿ No Use-p��Ϝ�0�NPO�\򁋁��.�oCH_L�������q	��s�MAVGAIL�����糅���SPACE1 ;2��, j�߂ �D��s�߂� �{~S�8�?�k� v�k�Z߬��ߤ��ߚ � �2�D���hߊ�|� ��`��������� � �2�D��h��|� ��`���������y���2����0�B��� f�����{���3);M_ ������/� /44FXj |*/���/�/�/?(??=?5Q/c/u/ �/�/G?�/�/�?O�? $OEO,OZO6n?�? �?�?�?dO�?�?_,_@�OA_b_I_w_7�O �O�O�O�O�_�O_(o�Ioo^oofo�o8 �_�_�_�_�_�oo6o Ef){����G �o� t���
M� � ��*�<�N�`�r����� ��w���o�収���d.��%�S�e�w� ����������Ǐَ�� �Θ8�+�=�k�}��� ����ůׯ͟���� %�'�X�K�]������� ��ӿ������#��E�W� `� @�������x�����\�e���������� �R�d߂�8�j߬߾� �ߒߤ���������� 0�r���X�����������8����
��ύ�_MODE�  �{��S E��{|�2�0�����3�	S|)�CWORK_AD޳�B�(+R  �{�`� �� _INTVAL����d���R_OPT�ION� ���H VAT_GRPw 2��upG(N�k |��_���� �/0/B/��h�u/T�  }/�/�/�/�/�/�/ ?!?�/E?W?i?{?�? �?5?�?�?�?�?�?O /OAOOeOwO�O�O�O �OUO�O�O__�O=_ O_a_s_5_�_�_�_�_ �_�_�_o'o9o�_Io oo�o�oUo�o�o�o�o �o�o5GYk- ���u���� �1�C��g�y���M� ����ӏ叧�	��-� ?�Q�c����������� ����ǟ�;�M��_����$SCAN�_TIM��_%�}�R �(�#�((�<04Wd d 
�!D�ʣ��u��/�����U�"�25�����dA�8�"H�g��]	����������dd�x�  �P���� ��  8� ҿ�!���D��$�M�_� qσϕϧϹ�������p�ƿv���F�X��/� ;��ob��pm��?t�_DiQ̡>  � l�|� ̡ĥ�������!�3� E�W�i�{������ ��������/�A�S� e�]�Ӈ��������� ����);M_ q������� r���j�Tfx �������/ /,/>/P/b/t/�/�/�/�/�/�%�/  0 ��6��!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O*�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko�O�OJ�o�o�o�o �o�o�o 2DV hz������0�
�7?  ;�>� P�b�t���������Ǐ ُ����!�3�E�W��i�{�������ß �ş3�ܟ��&�8� J�\�n�����������a�ɯ����,�� �+�	12345678�ү 	� =5����f�x��������� ����
��.�@�R� d�vψϚ�៾����� ����*�<�N�`�r� �߳Ϩߺ�������� �&�8�J�\�n�ߒ� ������������"� 4�F�u�j�|������� ��������0_� Tfx����� ��I>Pb t������� !/(/:/L/^/p/�/@�/�/�/�/�/�2 �/?�#/9?K?]?�iCz  Bp˚_   ��h2���*�$SCR_G�RP 1�(�U�8(�\x}d�@ �� �'�	 �3 �1�2�4(1*�&�I3��F1OOXO}m���D�@�0ʛ)����HUK�LM-10iA 890?��90;��F;�M61C D�:�CP��1
\&V�1	�6F@��CW�9)A7Y	(R@�_�_�_�_�_�\���0i^�oOUO >oPo#G�/���o'op�o�o�o�oB�0!�rtAA�0*�  @�Bu&Xw?��ju�bH0{UzAF@ F�`�r ��o�����+� �O�:�s��mBqrr��0��������B�͏b� ���7�"�[�F�X��� |�����ٟğ���N��@�AO�0�B�CU
L����E�jqBq>HE�̔�$G@�@pϯ B���G�I
E�0�EL_DEFAU�LT  �T���E��M�IPOWERFL�  
E*��7�W7FDO� *��1�ERVENT 1O���`(�� �L!DUM_E�IP��>��j!?AF_INE�¿�C�!FT���丿�!o:� ���a�!RPC_OMAINb�DȺPϜ��t�VIS}�Cɻ�����!TP��P�U�ϫ�d��E�!
�PMON_PROXYF߮�e4ߑ���_ߧ�f����!R?DM_SRV�߫�9g��)�!R�Iﲰ�h�u�!
v�M�ߨ�id���!R�LSYNC��>��8���!ROS��4��4��Y�(�}� ��J�\����������� ��7��["4F �j|����!��Eio�ICE�_KL ?%�� (%SVCPRG1n>���3�"�3���4//"�5./3/�6V/[/�7~/�/��D�/�	9�/�+�@��/� �#?��K?��s? � /�?�H/�?�p/ �?��/O��/;O� �/cO�?�O�9?�O �a?�O��?_��? +_��?S_�O{_� )O�_�QO�_�yO�_ ��Os����>o �o}1�o�o�o�o�o�o �o;M8q\ �������� �7�"�[�F��j��� ����ُď���!�� E�0�W�{�f�����ß ���ҟ���A�,� e�P���t���������ί�y_DEV ���MC�:�@`!�O�UT��2��REC 1�`e�j�� �� 	  �����˿���ڿ��
 �`e���6� N�<�r�`ϖτϦ��� ��������&��J�8� n߀�bߤߒ��߶��� ����"��2�X�F�|� j������������ ��.�T�B�x�Z�l� ������������, P>`bt�� ����(L :\�d���� � /�$/6//Z/H/ ~/l/�/�/�/�/.��/ ?�/2? ?V?D?f?�? n?�?�?�?�?�?
O�? .O@O"OdORO�OvO�O �O�O�O�O�O__<_ *_`_N_�_�_x_�_�_ �_�_�_oo8oo,o no\o�o�o�o�o�o�o �o�o "4jX �������� ��B�$�f�T�v��� ���������؏���>�,�b�P�r���p�V� 1�}� P
���!��� �y���TYPE\���HELL_CFOG �.��Ϗ  	�����RSR������ӯ�� �����?�*�<�u� `������������+����%�3�PE��Q�\�ӐM�Lo�p��d��2Ӑ�d]�K�:�HK 1�H� u����� ��A�<�N�`߉߄� �ߨ������������&�8��=�OMM ��H���9�FTOV_ENB&�1��OW_REG_U�I��8�IMWAI�T��a���OUTr������TIM��w���VAL��>��_UNIT��K��1�MON_ALI�AS ?ew� ( he�#������ ����Ӕ��);M ��q����d� �%�I[m �<����� �!/3/E/W//{/�/ �/�/�/n/�/�/?? /?�/S?e?w?�?�?F? �?�?�?�?�?O+O=O OOaOO�O�O�O�O�O xO�O__'_9_�O]_ o_�_�_>_�_�_�_�_ �_�_#o5oGoYokoo �o�o�o�o�o�o�o 1C�ogy�� H����	��-� ?�Q�c�u� ������� ϏᏌ���)�;�� L�q�������R�˟ݟ �����7�I�[�m� �*�����ǯٯ믖� �!�3�E��i�{��� ����\�տ����� ȿA�S�e�wω�4ϭ� �����ώ����+�=� O���s߅ߗߩ߻�f� ������'���K�]� o���>�������� ���#�5�G�Y��}����������o��$S�MON_DEFP�RO ������ �*SYSTEM�*  d=��R�ECALL ?}��� ( �}3�copy frs�:orderfi�l.dat vi�rt:\tmpb�ack\=>in�spiron:4804��r��o��}*.mdb:*.*CU
Y��6�	.x.:\�8@R�n���/.a6H_^�// �-?Qb/t/�/�/ �F/��/�/??) �M�/p?�?�?�8?�J?��? OO�%
x�yzrate 61 �?�?�?nO�O�O�%.GR(1228 HOZO�O�O_"/4/ �/�Ga_s_�_�_�/E_ �HY_�_�_o!?3?FO �C�_no�o�o�?6oHo �@^o�o&_8_�_ �_m��_�_�_Z ���"o4o�oXoi� {����o�oC��o��� �O0Oԏe�w���8�O�O�!064�OY� ����!�3���˟ݟ�n��������I2076G�Y�����!3 ���a�s������E� ��Y�����!�3�F� £ݿnπϒϥ�6�H� Š^�����&�8��� ܿm�ߑߤ���ȿZ� �����"�4���X�i� {��ϲ�C������� ��0�B�T�e�w��� �߮�I������� ,��P�as���� ;��`�(��@��o��&� ���desktop-�mbmd4ji:95248�Y�� /!3����o/�/�/&�!�@'10008 P/�/�/??*�;.�@��/�#i?{?�? �2��I?�,a?�?�OO$��$SNP�X_ASG 1�����9A�� P 0 �'%R[1]�@1.1O �?�$�%dO�OsO�O�O�O �O�O�O __D_'_9_ z_]_�_�_�_�_�_�_ 
o�_o@o#odoGoYo �o}o�o�o�o�o�o�o *4`C�gy �������	� J�-�T���c������� ڏ�����4��)� j�M�t�����ğ���� ��ݟ�0��T�7�I� ��m��������ǯٯ ���$�P�3�t�W�i� �������ÿ���� :��D�p�Sϔ�wω� �ϭ��� ���$��� Z�=�dߐ�sߴߗߩ� ������ ��D�'�9� z�]��������� 
����@�#�d�G�Y� ��}������������� *4`C�gy ������	 J-T�c��� ���/�4//)/ j/M/t/�/�/�/�/�/��/�/?0?4,DPA�RAM �9E}CA �	��:�P�4�0$HOF�T_KB_CFG�  q3?E�4PI�N_SIM  9K�6�?�?�?�0,@�RVQSTP_DSB�>�21On8J0�SR ��;� �& MULTI�ROBOTTAS�K=Oq3�6TO�P_ON_ERR�  �F�8�APT�N �5�@�A�BRINGo_PRM�O J0�VDT_GRP �1�Y9�@  	 �7n8_(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2Dkhz��� ����
�1�.�@� R�d�v���������Џ �����*�<�N�`� r���������̟ޟ� ��&�8�J�\����� ������ȯگ���� "�I�F�X�j�|����� ��Ŀֿ����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�tߛߘߪ߼����� ����(�:�a�^�p� ����������� � '�$�6�H�Z�l�~���������������3VP�RG_COUNTƛ6��A�5EN�B�OM=�4J_�UPD 1��;8  
q2�� ���� )$6 Hql~���� �/�/ /I/D/V/ h/�/�/�/�/�/�/�/ �/!??.?@?i?d?v? �?�?�?�?�?�?�?O OAO<ONO`O�O�O�O �O�O�O�O�O__&_ 8_a_\_n_�_�_�_YSDEBUG" ʇ �Pdk	�PSP�_PASS"B�?�[LOG �V�m�P�Xξ_  �g�Q
�MC:\d�_b_MPCm��o�o��Qa�o �vfSA/V �m:dUb��U\gSV�\T�EM_TIME �1�� (�`��S�2o	T1S�VGUNS} #'�k�spASK_?OPTION" ��gospBCCF�G ��| 8�b�{�}`��� �a&��#�\�G���k� ����ȏ������"� �F�1�j�U���y��� ğ���ӟ���0��T�f��UR���S��� ƯA������ ��D� �nd��t9�l������� ��ڿȿ�����"� X�F�|�jϠώ��ϲ� ��������B�0�f� T�v�xߊ��ߦؑ��� ����(��L�:�\� ��p���������� � �6�$�F�H�Z��� ~������������� 2 VDzh�� �������4 Fdv���� ��//*/�N/</ r/`/�/�/�/�/�/�/ �/??8?&?\?J?l? �?�?�?�?�?�?�?�? OO"OXOFO|O2�O �O�O�O�OfO_�O_ B_0_f_x_�_X_�_�_ �_�_�_�_oooPo >otobo�o�o�o�o�o �o�o:(^L np�����O� �$�6�H��l�Z�|� ����Ə؏ꏸ���� 2� �V�D�f�h�z��� ��ԟ����
�,� R�@�v�d��������� ίЯ���<��T� f�������&�̿��ܿ ��&�8�J��n�\� �π϶Ϥ�������� ��4�"�X�F�|�jߌ� �ߠ����������� .�0�B�x�f��R��� ���������,��<� b�P�������x����� ����&(:p ^�������  6$ZH~l ��������/ &/D/V/h/��/z/�/��/�/�/�&0�$T�BCSG_GRP� 2��%��  �1 
? ?�  /?A? +?e?O?�?s?�?�?�?��?�;23�<d�, �$A?1	� HC���6>�@E�5CL  �B�'2^OjH4Jݸ�B\)LFY g A�jO�MB��?F�IBl�O�O�@�JG|_�@�  D	�15_ __$YC-P{_F_$`_j\��_�]@0�> �X�Uo�_�_6oSoo�0o~o�o�k�h�0	V3.00'2�	m61c�c	�*�`�d2�o�e>əJC0(�a�i �,p�m-  �0�����omvu1JC�FG ��%� 1 #0vz��rrBrv�x�� ��z� �%��I�4� m�X���|�������� ֏���3��W�B�g� ��x�����՟����� ���S�>�w�b��� ��'2A ��ʯܯ��� ���E�0�i�T���x� ��ÿտ翢����/� �?�e�1�/���/�� �Ϯ��������,�� P�>�`߆�tߪߘ��� ���������L�:� p�^��������� ��� �6�H�>/`�r� ���������������  0Vhz8� �����
. �R@vd��� ����//</*/ L/r/`/�/�/�/�/�/ �/�/�/?8?&?\?J? �?n?�?�?�?�?���? OO�?FO4OVOXOjO �O�O�O�O�O�O__ �OB_0_f_T_v_�_�_ �_z_�_�_�_oo>o ,oboPoroto�o�o�o �o�o�o(8^ L�p����� ��$��H�6�l�~� (O����f�d��؏� ��2� �B�D�V����� ��n����ԟ
���.� @�R�d����v����� ���Я���*��N� <�^�`�r�����̿�� �޿��$�J�8�n� \ϒπ϶Ϥ������� ߊ�(�:�L���|�j� �߲ߠ���������� 0�B�T��x�f��� �����������,�� P�>�t�b��������� ������:(J L^������  �6$ZH~ l��^���dߚ  //D/2/h/V/x/�/ �/�/�/�/�/�/?
? @?.?d?v?�?�?T?�? �?�?�?�?OO<O*O `ONO�OrO�O�O�O�O �O_�O&__6_8_J_ �_n_�_�_�_�_�_�_ �_"ooFo��po�o ,oZo�o�o�o�o�o 0Tfx�H� ������,�>� �b�P���t������� ��Ώ��(��L�:� p�^�������ʟ��� ܟ� �"�$�6�l�Z� ��~�����دꯔo� �&�ЯV�D�z�h��� ����Կ¿��
��.π�R�@�v�dϚτ� s ���� ��������$TBJO�P_GRP 2����� O ?������������x/JBЌ��9�� �< �zX���� @����	 �C�� >t�b  C����>��͘Րդ��>̚йѳ33=��CLj�ff�f?��?�ffB@G��ь�����t�ц��>�(�\)��ߖ�E噙�;���hCYj��  �@h��B�  A�����f��C� � Dhъ�1���O�4�N����
�:���Bl^���j�i�l�l����A�ϙ�A�"��D��֊=qH������p�h�Q�;��A�j�ٙ7�@L��D	2��������$�6�>B�\p��T���Q�tsx�@33@���C����y�1����>G��Dh�������<���<{�h�@i� ��t� �	���K&� j�n|���p��/�/:/k/�ԇ����!��	V3�.00J�m61cI�*� IԿ��/��' Eo��E��E���E�F���F!�F8���FT�Fqe\�F�NaF����F�^lF����F�:
F�)�F��3G��G��G���G,I�!CH`��C�dTDU��?D��D���DE(!/E\��E��E�h��E�ME���sF`F+'�\FD��F`�=F}'�F���F�[
F����F��M;��;WQ�T,8�4` *Q�ϴ?�2���3�\�X/O��ESTP?ARS  ��	����HR@ABLE� 1����0��D
H�7 8��9
G
H�
H����
G	
H
�
H
HYE��
H�
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_Ht_�^:BS _� �J GoYoko}o�o�o�o�o �o�o�o1CU gy����`#oRL �y�_�_�_�_�O�O�O��O�OX:B�rNUM�  ����P��� V@P:B_?CFG ˭�Z��h�@��IMEBF_TT%AU��2@�GVERS�q���R 1���
 (I�/����b� �� ��J�\���j�|���ǟ ��ȟ֟�����0� B�T���x�������2��_���@�
��M�I_CHAN�� �� ��DBGLV����������ET�HERAD ?*��O�������xh�����ROUT�!��!������?SNMASKD��>U�255.���#������OOLOF/S_DI%@�u.��ORQCTRL �����}ϛ3rϧ� ����������%�7� I�[�:���h�z߯�A�PE_DETAI�"�G�PON_SV�OFF=���P_M�ON �֍�2���STRTCHK� �^�����VTCOMPAT���O�����FPROG� %^�%MU�LTIROBOT�Tݱ���9�PLA�Y&H��_INST+_Mް �������US�q��LCK����QUICKM�E�=���SCRE�Z�G�tps� ���u�z�����_��@@n�.�SR_�GRP 1�^�/ �O���� 
��+O=sa�쀚�
m���� ��L/C1g U�y����� 	/�-//Q/?/a/�/�	123456�7�0�/�/@Xt�1����
 �}i�pnl/� gen.htm�? ?2?�D?V?`Pan�el setupZ<}P�?�?�?�?�?�? �??,O>OPO bOtO�O�?�O!O�O�O �O__(_�O�O^_p_ �_�_�_�_/_]_S_ o o$o6oHoZo�_~o�_ �o�o�o�o�o�oso�o 2DVhz�1 '���
��.�� R��v���������Џ|G���UALRM��oG ?9� � 1�#�5�f�Y���}��� ����џן���,���P��SEV  �����ECFG ��롽�}A��   BȽ�
 Q���^���� 	��-�?�Q�c�u���Й��������� P�����I��?����(%D�6� �$�]� Hρ�lϥϐ��ϴ��π����#��G���� ��߿U�I_Y�H�IST 1�� � (�� ���3/SOFTP�ART/GENL�INK?curr�ent=edit�page,��,1����!�3��� �����menu��962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V