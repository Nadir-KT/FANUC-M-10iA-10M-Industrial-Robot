��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ����ALRM_�RECOV1   $ALMO�ENB��]ON�i�APCOUPwLED1 $[�PP_PROCE�S0  �1��GPCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y12 � u3�|4|GRG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WAx�471�:OFF_ �N�3DELHLO�Gn25Aa2?i1@N?�� -M��H W+0�$Y �$DB� 6COM�W!2MO� "0CyL]C.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2�X�D�#
 d �$CARD_E�XIST4$FSSB_TYP~uAHKBD_S�B֒1AGN Gn �$SLOT_N�UMJQPREV�,DBU� g1G ;1_�EDIT1 �� 1G=� S<�0%$EP�O$OP�A�ETE_OKRU�S�P_CRQ�$;4�V� 0LACIw1�RAPk �1�x@ME@$D�V�Q�Pv�A{�oQL� OUzR A,mA�0�!� B� OLM_O�^eR�"�CAM_;1 �xr$ATTqR4NP� ANN�@�5IMG_HEI�GHQ�cWIDTMH4VT� �UU0F_ASPECQw$M�0EXP�v�@AX�f�CFT� X $GR�� � S�!�@B@N�FLI�`t� UI�RE 3dTuGITC�HC�`N� S�d_�L�`�C�"�`ED(lpE� J�4S�0� ��zsa�!ip;G0� � 
$WARNM�0f�!,P� �s��pNST� CORyN�"a1FLTR�u�TRAT� T�p H0ACCa1��8�{�ORI
`"S�={RT0_S�BMֱpHG,I1 E[ Tp�"3I9��TY12`�K*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6��U7��8��94�qO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS�`�}Aw��"�tP_*0wOFSzR @� �RO_K8���aIT<�3��NOM_�0�1iĥ3nQCPT� �� $���AxP��K}EX�� �0g0�I01��p�
$TF�a��C$MD3��T�O�3�0U� �� K�Hw2�C1|�	EΡg0wE{vF�vF���p@�a2 m
P$A`PU�3N)#�dR*��AX�!sDETAI�3BUFV��p@1� |�p۶�pPIZdT� PP[�MZ��Mg�Ͱj�F[�SIMQSI�"0��A.�t���Pkx Tp�|zM��P�B�FAkCTrbHPEW7�`P1Ӡ��v��MCd�� �$*1JB8�p<�*1DECHښ��H���b� � �+PNS_EMP���$GP���,P_���3�p�@Pܤ��TC��|r��0�s��b��0�� �B���!
���J�R� ��SEGFRR��Iv �aR�Tkp9N&S,�PVF4��>� &k�Bv �u�cu��aE�� !2��p+�MQ��E�SIZ�3����T��P�����>�aRSINF��� ��kq���������LX�����F�CRCMu�3CClpG��p� ��O}���b�1��������2�V�DxIC��C ���r����P��{� SEV �zF_�եF�pNB0�?�p�����A�! �r �Rx����V�lp�2�@�aR�t�,�g�RTx #�5�5H"2��uAR���`CX�'$LG�p��B�1 `s�P�t�aA�0{�Уb+0R���tME�`0!BupCrRA 3tCAZ�л�pc�OT�#FC�b�`�`FNp��8�1��ADI+�a %��b�{��p$�pSp�c�`S�P��a,Q�MP6�`Y�3��M�'�pU��aU � $>�TITO1��S�S�!��$�"0�D�BPXWO��!���$SK��2
&�@DB�"�"@�;PR� 
� ����# >�q1M$��$��+�L9!$?(�V�%@?�A/��PC&_?R4gENE��'~?�(�� RE�pY2(�H �OS��#$L�3$$3R�h�;3�MVOk_D@!V�ROScrr�w�S����CRIGGER�2FPA�S��7�ET�URN0B�cMR_���TUː[��0EkWM%���GN>`���RLA���Eݡ<�P�&$P�t�'�@4a��C�DϣV��DXQ��4�1��MVG�O_AWAYRM�O#�aw!�D�CS_)  `IS#� �� �s 3S�AQ汯 4Rx�@ZSW�AQ�p�@1UW��NcTNTV)�5RV
a�����|c�éWƃ��J�B��x0��SAFE�ۥ�V_SV�bEX�CLUU�;��ONL��cYg�~az��OT�a{�HI_V�? ��R, M�_ �*�0� ��_z�2�� RCdSGO  +�rƐm@�A�c~b���w@��V�i�b�fANNUNx0�$�dKIDY�UABc�@ Sp�i�a+ �j�f�ΰ�APIx2,��$F��b�$ѐOT�@A� $DUMMY ��Ft��Ft±� 6�U- ` !�HE�|s��~bc�B@ �SUFFI��V4PCA�Gs5Cw�6Cq���DM�SWU. 8!�KgEYI��5�TM�10�s�qoA�vINޱE��!, / D��H7OST�P!4����<���<�°<��p<�E�M'���Z�� SBL�� UL��0  ��	����DT��01 � $|��9USAMPL�@��/���決�$ I@|갯 $SUBӄ���w0QS�����#��SAV�����c�S< X9�`�fP$�0E!�� YN_B�#2 M0�`DI�d�pO|��m��#$F�R_I�C� �ENC2s_Sd3  ��< 3�9���� cgp����4�"��2�A9��ޖ5���`ǻ�@Q@K&D-!�a�AVER�q��λ�DSP
���PC�_�q��"�|�ܣ�V7ALU3�HE�(��M�IP)���OP5Pm �TH�*�D�S" T�/�Fb�B;�d����d D�qм�16 H(rLL_DUǀ�a�@��0k���֠OT�"U��/���@@NOAUkTO70�$}�Hx�~�@s��|�C ����C� 2v�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3�T�3a�3n�4|¸�'����9 A<���z�ΓKI��0��H硵BaFEq@{@�: ,��&a?3 P_P?��>�J����E�@��r��RP��;fp$T�P�$VARI�����,�UP2Q`< W�߃TD��g���П`��������BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P"@��Fl@``>t ;��6����ST����T ��M ����0	��i� ��F���������kRt �����FORCEUyP�b܂FLUS
p�H(N��� ��6bD_CM�@E�7N�� (�v�P��REM� Fa��@j����
K�	N���EcFF/���@IN�Q�OV��OVA��	TROV DyT)��DTMX: e �P:/��Pq�XvXpCLN _�p���@ ��	_|��_QT: �|�&PA�Q	DI���1���0�Y0RQm�_�+qH���M���CL�d#�RIV{�ϓN"�EAR/�IO�P�CP��BR��C�M�@N 1b 3GgCLF��!DY�(ء�a�#5T�DG����� �%%�FSS� )�? P(q1�1��`_1"811R�EC13D;5D6O�GRA���@��i���PW�ON2EBUG�S�2��C`gϐ_E A� ��?����TE�RM�5B�5��O�RIw�0C�5tio�SM_-`���0�D�5o�TA��9EIUP��Fg� -QϒA�P|�3�@B$SEGGJv� EL�UUSEPNFI��pBx��1x@��4>DC$UF�P��$���Q�@C���G�0T�����SwNSTj�PATۡ<g��APTHJq�A�E*�Z%qB\`F�{E���F�q�pARxPY�aS�HFT͢qA�AX_�SHOR$�>��6 �@$GqPE���O#VR���aZPI@P@$�U?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi� [Y)��G�@R��i�e԰�i�R�!P�uAScYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UaP���P���WOR�@�M��k0SMT��G��GR��3�a�PA�@��p5�'�H� � j�A�T�OCjA7pP]Pp$OPd�O��C�%��p�O!��RE.pR�C�AO�?��Be5pR�EruIx'Q�G�e$PWR) IMdu�RR_$sp�5�.�B Iz2H8�=��_ADDRH�H_LENG�B�q�q:��x�R��So�J.�SS��SK������ ��-�SE*���rmSN�MN1K	��j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ���p�Q� ��OUPW3��b_>�I��!q�a1 ��������|��� �����-���:���i+IOX2S=�D�e�x�]���L $��<p�!_OFF[r_�oPRM_�N�a�TTP_�H��M; (�pOBJ�"�p�G�$H�LE�C|��ٰN � 9�.*�AB_�T��
��S�`�S��LV��K�RW"duHITCOmU?BGi�LO�q����d� Fpk��GpSS� ���HW�h�wA��O.��`I�NCPUX2VISIO��!��¢.�á�<�á-� �IOL]N)�P 87�R'�^[p$SL�bd oPUT_��$dp��Pz �� F_�AS2Q/�$L D���D�aQT U�0]PA������PHY`G灱Z���5�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp����x��ٶ�1UJ���S����NE�WJsOG�G �DIS��b&�KĠ��3T |���AV��`_�CTR<!S^�FLAGf2r�;LG�dU �n�:���3LG_SIZ���ň��=���FD��I����Z �ǳ� �0�Ʋ�@s��-ֈ�-ր=�-���-��0-�ISGCH_��Dq��N?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHrܭ�I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn���_BWUFF1XY��PT�$�� �v���fĵ�1�A�rYY���P �����pOS1J�2�3���_�>0Z �  ��apiE�*��IDX�d	P�RhrO�+��A&+ST��R��Yz�<!� Y$EK&C K+���Z&m&KF�1[ L��o�0��]P�L�6pwq�t^����tN�V�7�_ \ �`��瀰�7��#�0�C��] ��CL�DP��;eTRQL�I�jd.�094FLAGz�0r1R3�DM��R7��LDR5<4R5ORG.���e2(`���V��8.��T<�4�d^ A�q�<4��-4R5S�`�T00m��0DFRCLMC!D�?�?3I�@��MIC��d_ Yd���RQm�q��DSTB	�  ؏Fg�HAX;b |�H�LEXCESZr��rBMup�a`��B;d �
qC`��`5a��F_A�J���$[�O�H0K�db q\��ӂS�$MB���LIБ}SREQU�IR�R>q�\Á�XD�EBU��PT�ML� MP�c�ba��Ph؃ӂ!BoAND�ф�`�`d�҆�c�cDC1��IN�����`@�(h?Nz�@q��o����RPST8� �e�rLOC�RYI�p�EX�fA�px��AoAODAQP�7f X��ON��[rMF�����f)�"I�`�%�e��T���FX�@�IGG� g �q��"E�0��#���$R�a%;#7y��Gx�VvCPi�DATAw�pE:�y�[�Eѭ��NVh t $+MD�qIё)�v+�tń�tH�`�P�u�<|��sANSW}��t(�?�uD�)�b��	@Ði �@CU���V�T0�eRR2�j Dɐ�Qނ�B?d$CALI�@F��G�s�2�RIN���v�<�INTE���kE���,��b����_Nl��ڂ���kDׄRm�DIVFiFDH�@ـn��$V��'c!$��$Z������~�[��oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS�@#2L  �Ė83ಀ����� ��PAT!H��������3̒Vp�A_�Q�.�4�B��Cᐈ�_MGh��$DDQ���G�$FWh��p��m������b�DE��PPAB�NԗROTSPE!ED����00J�Я�8��@��̐$US�E_��P��s�S�Y��c�A kqYNru@Ag��OFF�qn�MOUN�NGg��K�OL�H�INC *��a��q��Bj�L@�BENCS��q�BđX���D��IN#"I̒0��4�\BݠVEO�w�>Ͳ23_UPE�߳/LOWL���00����D���Bp���� �1RCʀƶMO3SIV�JRMO���@�GPERCH  �OV��^��i� <!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸUPp������TRKr�>"AYLOA'a��  Q-�̒<�1Ӣ`0 ���RTI$Qx�0 MO ���МB R�0J��D���s�H����b�DU�M2(�S_BCKLSH_C̒��>� =�q�#�U��ԑ���2�<t�]ACLALvŲp�1n�P�CHK00:'%SD�RTY4�k���y�1�q_6#2�_�UM$Pj�Cw�_�S�CL��ƠLMT_OJ1_LO��@���q��E�����๕�幘SPC��7���L���PCo���H� ȰPU�m�C/@�"XT\_�c�CN_��N��Le���SFu���V��&#����9�̒��=�C�u�SH6#��c��� �1�Ѩ�o�0�͑
��f_�PAt�h�_Ps�W�_10��4�R�01D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�sR0Hљ��_W��-ԁ_=��C��I��I*�I�II�F�`�aJLA.�1[�VC��0�D�BO1U�@i�B\JRKU��~	@DBL_SMd�:BM%`_DLC�BGRV��C��I���H_� �*CcOS+\�(LN� 7+X>$C�9)I�9)u*c,)�Z2 HƺcMY@!�( "TH&-��)THET0�N�K23I��"=�A C-B6CB=�C�A�B�(261C�616SB8C�T25GTS QơC��aS$" �4c#<�7r#$DUD�EX��1s�t��B�6���AQ�|r�f$NE�DpI B U�\B5��$!��!�A�%E(G%(!LCPH$U�2׵�2SX pCc%pCr%�2�&�C�J�&!�VAHV6H3�YLUVhJVuKV�KV�KUV�KV�KV�IHAH@ZF`RXM��wXuKH�KUH�KH�KH�KH�I�O2LOAHO�YWNO�hJOuKO�KO�KO*�KO�KO�&F�2#1�ic%�d4GSPBA?LANCE_�!�c�LEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%�Ċ1ky�UTO_<?�jT1T2Cy��2N&�v�ϰctw�gѠp�0Ӓ~���T��O����� INSEGv�!�REV�v!���gDIF��1l�w6�1m
�OB�q
����MIϰ1��L�CHWAR����A�B&u�$MEC�H,1� :�@�U�AX�:�P��Y�G$�8pn� 
Z��|���RO�BR�CR̒��N�'�MSK_�`�f�p P Np_���R����΄ݡ�1 ��ҰТ΀ϳ��΀"��IN�q�MTC�OM_C@j�q � L��p��$ONORE³5����$�r 8� GRl�E�SD�0ABF��$XYZ_DAx5A���DEBU�qXI��Q�s �`$�wCOD�� ���k�F�f�$BU�FINDXР � ��MOR��t $-�U��)��rФB���͓�Gؒu� � $SIMULT ��~�� ����OBJE�` �AD�JUS>�1�AY_	Ik��D_����C��_FIF�=�T � ��Ұ��{��p� ��З��p�@��D�FRiI��ӥT��RO� Ұ�E�{�͐OPsWO�ŀv0���SYSBU�@ʐ$�SOP����#�U<"��pPRUN�I�PA�DH�D����_OU�=��qn�{$}�IMAG��iˀ�0P�qIM��Ơ�IN�q���RGOVRDȡ:���|�aP~���Р�0L_6p0���i��RB���0e��M���EDѐ*F� ��N`M*�����̰SL�`ŀw �x $OVSL�vSDI��DEX�m�g�e�9w�����V� ~�N���w�����h�ǖȳ�M�J͐��q<��� x HxˁE�F�ATUS�Ѕ�C�0àǒ��BSTM����If����4����(�ŀy DBˀEz�g���PE�r������
���EXE ��V��E�Y�$Ժ ŀgz @ˁ��UP{�fh�$�p��XN����9�H� �P�G"�{ h $GSUB��c�@_��|01\�MPWAI��P����LO��<�F��p�$RCVF�AIL_C�f�B�WD"�F���DEF�SPup | L�ˀ`�D�� U�UCNI��S���R`Ь��_L�pP��%���P�ā}��� @B�~���|��`ҲN�`�KET��y���Pԙ $�~���0SI�ZE��ଠ{���S�<�OR��FORMAT/p � F���r�EMR��y�UX8����PLI7�ā�  $�P�_SWI������_PL7�AL_� �ސR�A��B��(0C��Df�$mEh����C_=��U� � � 1���~�J3�0��^��TIA4��5��6��MOM������� �B�AD`��*��* PU70NRW��W ��U����� A$PI�6���	�� )�4l�}69��Q�|��c�SPEED�PGq�7�D�>D�� ���>tMt[��SAM�`痰>��MOV���$�@�p�5��5�D�1�$2�������{�2��Hip�IN?,{� �F(b+=$�H*�(_$<�+�+GAMM�f�1>{�$GET��Đ�H�D����
^pLI�BR�ѝI��$H�I��_��Ȑ*B6Eď�*8A$>G086LW =e6\<G9�686��R���ٰV��$�PDCK�Q�H�_����;"��z�.%��7�4*�9� ��$IM_SR�O�D�s"���H�"�L	E�O�0\H��6@�R� �ŀ�P~�qUR_SCR����AZ��S_SAV�E_D�E��NO��CgA�Ҷ��@�$�� ��I��	�I� %Z[ � ��RX" ��m�� �"�q�'"�8� Hӱt�W�UpS���%���L;@���O㵐 .'}q��Cg���@ʣȳ���S�M�AÂ� ?� $PY��g$WH`'�NGp� ��H`��Fb��Fb��Fb��PLM���	� 0h�H�{�X��O��z�Zp�eT�M���� pS��C��O__0_�B_�a��_%�� | S����@	�v��v  �@���w�v��EM��%� �Cfr�B�ːt��ftP��PM���QU� �U�Q���Af�QTH=�H{OL��QHYS�3ES�,�UE��B���O#��  ��P�0�|�gAQ���ʠu���O��ŀ�ɂv�-�8�A;ӝROG��a2D�E�Âv�_�Ā^Z�INFO&��+�h���b�R�OI��� ((@SLEQ /�#������o���S`c0O�0�051EZ0NUe�_��AUT�Ab�COPAY��Ѓ�{��@M���N�����1�P�
� ���RGI�����X_�Pl�$�����`
�W��P��j@�G����EXT_CY�CtbR��p�����h�_NA�!�$�\�<�RO�`]��� � m��P�OR�ㅣ���SReVt�)����DI �T_l���Ѥ{�ۧ�Шۧ �ۧ5٩6٩7�٩8����S�B쐒���$�F6���PL�A�A^�TAR ��@E `�Z������<��d� ,(@FL�q`h��@YNL���Mz�C���PWR���쐔e�DELA�Ѱ�Y�pAD#q�Q�QSKIP��� ĕ�x�O�`NT2!� ��P_x��� ǚ@�b�p1�1� 1Ǹ�?� �?��>���>�&�>�3�>�9��J2R;쐖 46��EX� TQ���� ށ�Q���[�KFд��w�RDCIf� �U`�X}�R�#%M!�*�0�)��$RGEA�R_0IO�TJBFcLG�igpERa�TC݃������2T�H2N��� 1�� �Gq TN�0 ����M����`Ib���AREF:�1�� l�h���ENAB��lcTPE?@���!(ᭀ�� ��Q�#�~�+2 H�W���2�Қ���"�4�F�X�����3�қ�{��������j�4�Ҝ��
��.�@�R�
j�5�ҝu�������(����j�6�Ҟ���(:L��7�ҟ�o�����j�8�Ҡ��"4F�j�SMSK�� Q �+@��E�A���REMOTE������@ "1��Q�IO�5"%I��Pt����POWi@쐣  �����X�gpi������Y"$DSB_SIGN4A�Qi�̰�C���tRS232�%�Sb�iDEVI�CEUS#�R�RP�ARIT�!OP�BIT�Q��OWCONTR��Qⱬ��RCU� M�SU_XTASK�3NB���0�$TATU�P#H�"@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�U�PDl�ARB�SP|%0���� !m$USA���az9�L�ERI�0f��p�RY�5~"_�@f�P8�1�!�6WRK���D9�F9ХFRIgEND�Q4bUF���&�A@TOOLHFM�Y5�$LENG�TH_VT��FI!R�pqC�@�E� IOUFIN�R����RGI�1�AIT�I:�xGX��I�FG2�7G1a����3�B��GPRR�DA��O_0� o0e�I1RER�đ�3&���TC���AQ�JV�G|�.2���F��1�!d�9Z�8+5�K�+5��E�y�L0�4�OX �0m�LN�T�3Hz��89��%�4J�3G��W�0�W�RdD�Z��Tܳ��K��a3d��$cV C2���1��I1H��02K2sk3K3 Jci�aI�i�a�L���SL��R$Vؠ�BV�EVk��A bQ*R��� �,6Lc���9V`2F{/P:B��PS_�Et�$rr�C�ѳg$A0��wPR���v�U�cSk�� {��$�1��� 0���VX`�!�tX`��0P��Ё�
�5SK!�� �-qR��!0�4��z�NJ AX�!h��A�@LlA��A�THIC�1�������1�TFE���q>�IF'_CH�3A�I0�����G1�x������t9�Ɇ_JF҇�PR(���RVA=T�� �-p���7@����DO�E��CsOU(��AXIg��OFFSE+�TRIG�SK��c������e�[�K�Hk���8��IGMAo0�A-���ҙ�ORG_UNsEV��� �S�~쐮d �$��z����GROU���ݓTO2��!ݓDSP��JOG'��#	�_P'�2OR����>P6KEPl�IR��0�PM�RQ�AP��Q��E�0q�e���ScYSG��"��PG��BRK*Rd�r�3�-��������ߒ<pADx��ݓJ�BSOC�� N�DUMMY�14�p\@SV�PD�E_OP3SFS�PD_OVR��bٰCO��"�OR-��N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA��"LCHDL�R�ECOV��0�Wb�@M�յ�RO3���_�0� @܄ҹ@VERE�$7OFS�@CV� 0BWDG�ѴC��2j��
�TR�!��E�_FDOj�MB_�CM��U�B �BL =r0�w�=q�tVfQ�Ґx0sp��_�Gxǋ�A�M��k�J0������_�M��2{�#�8$�CA�{Й���8$�HBK|1c��IO␅.�:!aPPA "�N�3�^�F���:"�?DVC_DB�C��@d�w"����!��1����ç�3����ATIEO� �q0�UC�&CAB�BS@�PⳍP�Ȗ��_0~c�SUBCPUq��S�Pa aá�}0�S�b��c��r"ơ$HW_C���:c��Ic�A�A-�l$UNI5T��l��ATN�f�����CYCLųN�ECA��[�FLT?R_2_FI���(��}&��LP&�����o_SCT@SF_��aF����G���FS|!�¹�CHAA/���8��2��RSD�x"�ѡb�r�: _T��PcRO��O�� EM��_��8u�q 1u�q��DI�0e�?RAILAC��}RMƐLOԠdC��:a�nq��wq����PRJ��SLQ�pfC��z30	��FUNCŢ�rRINkP+a�0 ̆�!RA� >R �
Я�ԯWAR��BLFQ��A0�����DA�����LDm0�a�B9��nqBTI�vrbؑ���PRIA,Q1�"AFS�P�!������`%b���Mr�I1U�DF_j@ؖ�y1°LME�FA��@HRDY�4��P�n@RS@Q�0"�MULSEj@f�b�q� �X��ȑ����$.A$�1�$c1Ó���7� x~�EGvpݓ��q!AR����0�9>B�%��AXE.��ROB��W�A4�_�-֣SY���!6���&S�'WR���-1���STR��5�:9�E�� 	5B��=QB90�@6�������OT�0o 	$�ARY8�w20�Ԛ�	%�FI��;�$LINK�H��1%�a_63�5�q�2XYZ"��;�qH�3@��1�2�8{0	B�{D��� CFI��6G��
�{�_J��6��3NaOP_O4Y;5�FQTBmA"�BC
�z�DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ �@�5<:7�� W1�?0K�Mc��68Cb�vrb�4�ORQ��X�>8�#op ������wq�Uf����N�TOVE�Q��M;����E#�UK#�UQ"�VW �ZQ�W���Tυ� ;� ����QH�!`�ҽ��U��Q�WkeK#kecXE)R��	GE	0��S�dAWaǢ:D���0�7!�!AX�rB !{q��1uy-! y�pz�@z�@z6P z\Pz� z1v� y�y�+y�;y� Ky�[y�ky�{y�x�y�q�yDEBU��$����L�!º2WG`  AB!�,�r�SV���� 
w� ��m���w����1���1 ���A���A��6Q��\Q����!�m@��2CLAB3B�U������S = ÐER|���� � $�@ڳ Aؑ!p�PO���Z�q0w�^�_M�RAȑ� d r T�-�ERR�L�TYz�B�I�qV3@�cΑTOQ�d:`L� �d2ᕴP��|˰[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	V FZN_wCFG_!� 4�� ?º�|�ų����@�Ȳ�W ���\$� �n���Ѵ��9c�Q���(�FA�He�,�XEDM�(�����!s��Q�g�P{R�S�HELLĥ�� 56�B_BAS�!�RSR��ԣo ��#S��[��1r�%���2ݺ3ݺ4ݺ5*ݺ6ݺ7ݺ8ݷ���ROOI䰝0�0NLK!�CAB� ���ACK��IN��T�:�1�@�@ z�m�_�PU!�CO� ��OU��P� Ҧ) ��޶���TPFWD_�KARӑ��RE�~��P��(��QU�E�����P
��CSTOPI_AL������0&���㰑�0S#EMl�b�|�M��dЛTY|�SOK�}�D�I�����(���_�TM\�MANRQ�ֿ0E+�|�$K�EYSWITCH�&	���HE
�B�EAT����E� LQEҒ���U��FO������O_HOM��O�REF�PPARz��!&0��C+�9OA�ECO��B<�rIOCM�D8�µ����8�` � �D�1����U��&�M�H�»P�CFORC���� ��OM>�  � @V��*|�U,3P� 1-�`ʀ 3-�4��NP�X_ASǢ� 0�ȰADD����$�SIZ��$VA�Rݷ TIP]�\�2�A򻡐��Ȑ]�_� �"S꣩!C<ΐ��FRIF⢞�aS�"�c���NF�ҸV ��` � x�`S�I�TES�R6SSKGL(T�2P&���AU�� ) STMTdQZPm 6BW�P�*SHOWb���SV�\$�� ���A00P�a� 6�@�J�T�U5�	6�	7�	8�	9�	A�	� �!�'��C@�F�0u �	f0u�	�0u�	�@�u[Pu%121�?1L1Y1f1�s2�	2�	2�	2��	2�	2�	2�	2�22%222�?2L2Y2f2�s3P)3�	3�	3��	3�	3�	3�	3�33%323�?3L3Y3f3�s4P)4�	4�	4��	4�	4�	4�	4�44%424�?4L4Y4f4�s5P)5�	5�	5��	5�	5�	5�	5�55%525�?5L5Y5f5�s6P)6�	6�	6��	6�	6�	6�	6�66%626�?6L6Y6f6�s7P)7�	7�	7��	7�	7�	7�	7�77%727�?7,i7Y7Fi7�s�VP�UPD>��  ��|�԰��YSLOǢ� � z��и����o�E��`>�^t��АAcLUץ����CU��z�wFOqID_L��ֿuHI�zI�$F�ILE_���t���$`�CKuSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_ �TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅��L~�_Vj��'����� ` �GGROU�pD��B�NFLIC��R�EQUIREa�E�BUA��p����2�¯�����c��� \��APPR���C���
�EN��CLOe��S_!M v�,ɣ�
���o� ���MC�8&���g�_MG�q��C� �{�9���|�B;RKz�NOL��|�:� R��_LI|���$��k�J����P
��� ڣ�����&���/���Q6��6��8����|���� ���8�%�W�2�e�PATHa�z�p�z�=�vӴ��ϰ�x�CN=�CaA�����p�IN��UC��bq��CO�U�M��YZ������qE�%���2������PA�YLOA��J2L�3pR_AN��<�L���F�B�6�R�{�R_?F2LSHR��|�LOG��р��ӎ���ACRL_u��������.���H�p�$yH{���FLEX
��s�J�� :�/����6�2���0��;�M�_�F16�� ��n���������ȟ��Eҟ�����,�>� P�b���d�{�����@�������5�T��X��v���Eť mFѯ��������&�/�A�S�e�D�J>x�� � ������j�4pAT����n��EL  �%øJڪ��ʰJE��CTYR�Ѭ�TN��F&���HAND_VB�[
�pK�� $�F2{�6� �rS�Wi�D�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�(#�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������uN���2�H̟�����"CqENL� a�DI��>�Obt8C�Dpx�� ��2IxQA����q��-���s �� ����� ���OMME���rr�QTVpPT@�P ���qe�i�����P�x ��yT�Pj�� $DUMMY}9�$PS_��RFq�  ��:�� ���!~q� �X����K�STs��ʰSBR��M21�_Vt�8$SV_�ERt�O��z���C+LRx�A  O�r?p�? Oր � D $GLOB���#LO��Յ$�o���P�!SYSA�DR�!?p�pTCH>M0 � ,��ސ�W_NA���/�e�$%SR��l (:]8:m� K6�^2m�i7m�w9m� �9���ǳ��ǳ���ŕ ߝ�9ŕ���i�L� ��m��_�_�_�TDџXSCRE�ƀӚ� ��STF����}�pТ6�1] _:v AŁ� T����TYP�r�K��u�!u���O�@I�S�!��t.D�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J��*��AI=�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� D�C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!$1VSHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3��H���w�2u�b�V�rzu��%�DJU��~|#�WAIT�������%ONE���YBOư ?�� $@p%�vC�SBn)TPE��NEC��x"�$t$��.�*B_T��R��% �qR� ���sB�%�tM�+Z�t�.�F�R!�݀��OPm�MAS��_DOG�OaT	�D����C3S�	�O2DELAY���e2JO��n8E��Ss4'#�J�aP6%�����Y_��O2$��2���5���`? sqZA�BCS��  �$�2��J�
� �$�$CLAS�����AB�sp'@@�VIRT��O.@A�BS�$�1 <E�� < *AtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v���8��M@[�AXLրK��*B�dC  ���IqN��ā��PRE������LAR�MRECOV �<I䂥�NG�� �\K	 A  � J�\�M@PPLIMC�?<E�E��Handl�ingTool ��� 
V7.5�0P/28[�  o�����
�w_SW�� UP*A7� ��F0ڑ���AG@�� S20��*A���:�ާ�X�FB �7DA5�� �N'@��y@��None������� ��T���*A4y�+xl�_��V����:g�UTOB���������HGAPO�N8@��LA��U��D� 1<EfA����������� Q 1שI Ԁ��Ԑ�:�i�n��܍�#BGB �3��\�HE�Z��r�HTTHKY ��$BI�[�m����� 	�c�-�?�Q�o�uχ� �ϫϽ��������_� )�;�M�k�q߃ߕߧ� ���������[�%�7� I�g�m������� ������W�!�3�E�c� i�{������������� ��S/A_ew �������O +=[as�� �����K//'/ 9/W/]/o/�/�/�/�/ �/�/�/G??#?5?S? Y?k?}?�?�?�?�?�? �?COOO1OOOUOgO yO�O�O�O�O�O�O?_�	__-_K_Q_��(�T�O4�s���DO_C�LEAN��e��SN�M  9� ��9oKo]ooo�o�D?SPDRYR�_%�HI��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ|��g�PLUGGҠ��Wߣ��PRC�`B�`9��o�=�OxB��oe�SEGF��K������o%o�����#�5�m���LAP �oݎ����������џ �����+�=�O�a�>��TOTAL�.����USENUʀ�׫ �X���R(�RG�_STRING �1��
��M��Sc�
��_�ITEM1 �  nc��.�@�R�d�v� ��������п������*�<�N�`�r��I/O SIGN�AL��Try�out Mode��Inp��Simulated��Out��O�VERR�` = �100�In �cycl���P�rog Abor������Stat�us�	Hear�tbeat��M?H FaulB�K�AlerUم�s߅� �ߩ߻��������� �S���Q�� f�x���������� ����,�>�P�b�t�p������,�WOR�� ����V��
.@ Rdv����� ��*<N`PO��6ц��o �����//'/ 9/K/]/o/�/�/�/�/��/�/�/�/�DEV �*0�?Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�OPALTB��A�� �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_�oo(o:o�OGRI �p��ra�OLo�o�o�o �o�o�o*<N `r������`o��RB���o�>� P�b�t���������Ώ �����(�:�L�^�xp����PREG�N ��.��������*� <�N�`�r����������̯ޯ���&�����$ARG_��D �?	���i���  w	$��	[}��]}���Ǟ�\�SB�N_CONFIG� i��������CII_SAV/E  ��۱Ҳ�\�TCELLSE�TUP i�%�HOME_IO��͈�%MOV_8�2�8�REP����V�UTOBACK�
�ƽF�RA:\�� X�Ϩ���'` ���x������ �� ��$�6�c�Z�lߙ���������������� �!凞��M�_�q�� ���2��������� %�7���[�m������ ��@�������!3E$���Jo��p�����INI�@���ε��MESSAG����q�>�ODE_D$��ĳ�O,0.��PA�US�!�i� ((Ol���� ���� /�// $/Z/H/~/l/�/�'a~kTSK  qx�����UPDT%��d0;WSM�_CF°i��еU�'1GRP 2�h�93 |�B��A|�/S�XSCRD+1;1
1; ����/�?�?�? OO$O ��߳?lO~O�O�O�O �O1O�OUO_ _2_D_�V_h_�O	_X���GR�OUN0O�SUP�_NAL�h�	ܢĠV_ED� 1�1;
 �%-B?CKEDT-�_`�!oEo$���a�o�����ߨ���e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[8�5GED4�n�#�� ~�j���ED5Z��Ǐ6� ~��8�}���ED6�����k�ڏ ~G���!�3�ED7��Z��~� ~�8V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W�Ư�
}3�����CR o�����3�տ@ϯ�����P�PNO_DE�L�_�RGE_UN�USE�_�TLAL_OUT q��c�QWD_ABO�R� �΢Q��ITR�_RTN����N'ONSe����CAM_PARA�M 1�U3
 �8
SONY �XC-56 234567890�H� � @����?���( Щ�V�|[r؀~�X�HR5k�|U�Q��ο�R57����A�ff��KOWA SC310M|[�r�̀�d @6�|V��_�Xϸ� ��V��� ���$�6���Z�l��CE_RIWA_I857ЍF�1��R|].��_LIO4W=� ���P<~�F<�GwP 1�,����_GYk*C*�  ��C1� 9J� @� G� �CL�C]� d� l� s��R� ��[�m�� v� � �� ��� C�� �"��|W��7�HEӰON�FI� ��<G_P_RI 1�+P� m®/���������'CHKPAU�S�  1E� ,�>/P/:/t/^/�/ �/�/�/�/�/�/?(?@?L?6?\?�?"O������H�1_MO�R�� �XaB�iq-���5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`ϖ�S:�(����Yp0�_)o�S`�BBia�P�_mo8j�(�aKoo�o9i�(�E�og�o�o�m�o�f�oGq:I�ZDE�F f8��)��R6pbuf.txAtm�]n�@�����# 	`(Ж�A=L����zMC�21B�=��9���4�=��n׾�Cz  B�HBCCPUeB��_B�y;���>C���C�nSZE@E?{h�D]^Dْ�?r����D���^��G	��F���F��Cm�	fF�O�FٓΫSY���vqGR���Em�(�.����1(��<�q�G�)x2��Ң �� a��D�j���E�e��X��EQ�EJ�P F�E�F�� G���F�^F E�� F�B� H,- Ge��H3Y����  >�33 ����xV  n42xQ@��5Y��8B� A�AST<#�
�� �_'�%��wR_SMOFS���~�2�yT1�0DE ��O c
�(�;�"�  <�6�z��R���?�j�C4R��SZm� W���{�m�C��B-G�CR�`@$�q��T{��FPROG %i����c�I��� �����f�KEY_TB�L  �vM�u� ��	
�� �!"#$%&'(�)*+,-./0�1c�:;<=>?�@ABC�pGHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������p���͓���������������������������������耇�������������������s��!j�LCK��x.�j���STAT����_AUTO_D�O���W/�IND�T_ENB߿2R���9�+�T2w�XS�TOP\߿2TRL^l�LETE�����_SCREEN �ikcs�c��U��MMEN�U 1 i  <g\��L�SU+� U��p3g������ ������2�	��A�z� Q�c������������� ��.d;M� q������ N%7]�m ���/��/J/ !/3/�/W/i/�/�/�/ �/�/�/�/4???j? A?S?y?�?�?�?�?�? �?O�?O-OfO=OOO �OsO�O�O�O�O�O_��O_P_Sy�_MA�NUAL��n�DB;COU�RIG��ٟDBNUM�p���<���
�QPXWO_RK 1!R�ү��_oO.o@oRk�Q_�AWAY�S��G�CP ��=��df_CAL�P�db�RY��������X_�p 1"��� , 
�^@���o xvf`MT��I^�rl@�:sON�TIM�����ɼZv�i
õ�cMO�TNEND���dR�ECORD 1(�R�a��ua�O� �q��sb�.�@�R� �xZ�������ɏۏ 폄���#���G���k� }�����<�ş4��X� ��1�C���g�֟�� ������ӯ�T�	�x� -���Q�c�u������� ���>����)Ϙ� Mϼ�F�࿕ϧϹ��� :�������%�s`Pn&� ]�o��ϓ�~ߌ���8� J�����5� ��k� ���ߡ��J�����X� �|��C�U������ ����0�����	���dbTOLEREN�CqdBȺb`L��͐PCS_CFG� )�k)wd�MC:\O L%0?4d.CSV
�`�c�)sA �CH
� z�`)~����hMRC_OUT� *�[�nS�GN +�e�r���#�10-MA�Y-20 09:�26*V15-JA}Nj10:51�k P/Vt��)~�`pa��m��PJP���VERSIO�N SV�2.0.8.|EF�LOGIC 1,^�[ 	DX�P�7)�PF."PROG�_ENB�o�rj U�LSew �T�"_?WRSTJNEp�V��r`dEMO_OPT_SL ?	�e�s
 	R575)s7)�/??*?�<?'�$TO  ��-��?&V_@pE�X�Wd�u�3PA�TH ASA�\�?�?O/{ICTZ�aFo`-�gd>segM%&A�STBF_TTS��x�Y^C��SqqF��PMAU� t/XrMKSWR.�i�a.|S/�Z!D_N�O 0__T_C_x_g_�_�t�SBL_FAUL�"0�[3wTDIAbU 16M�ap�A�123456�7890gFP ?BoTofoxo�o�o�o �o�o�o�o,>�Pb�S�pP�_ ���_s�� 0`� ����)�;�M�_� q���������ˏݏ�|)UMP�!� �^�TR�B�#+��=�PMEfEI�Y_�TEMP9 È��3@�3A v�UNI��.(YN_BRK� 2Y)EMG?DI_STA�%W�ЕNC2_SCR 3��1o"�4� F�X�fv���������#��ޑ14���@�)�;�����ݤ5�����x�f	u� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/߭P�b� t�� ��xߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N���r��� ������������ &8J\n��� �����"`� FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/4?,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O?�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�O�O�o �o�o
.@Rd v������� ��*�<�N�`�r��� �o����̏ޏ���� &�8�J�\�n����������ȟڟ����H�E�TMODE 16v��� ���ƨ
R�d�v�נR�ROR_PROG7 %A�%�:߽��  ��TABLE  A�������#�L�RRSEV_?NUM  ��Q���K�S���_�AUTO_ENB�  ��I�Ϥ_N�Oh� 7A�{��R�  *����J��������^�+��pĿֿ迄�HISO��͡I�}�_ALM �18A� �;�����+�e�wωϐ�ϭϿ��_H���  A���|��4��TCP_VER �!A�!����$E�XTLOG_RE�Q��{�V�SI�Z_�Q�TOL  �͡Dz��A= Q�_BWD���иr���n�_DI�� 9��}�z�͡<m���STEP����|4��OP_DO����ѠFACTO�RY_TUN�d�G�EATURE �:����l��Handlin�gTool �� � - CEn�glish Di�ctionary���ORDEA�A Vis�� M�aster���9�6 H��nalo�g I/O���H�551��uto �Software� Update � ��J��mati�c Backup~��Part&��ground E�dit��  8\�apCame�ra��F��t\j�6R�ell���LwOADR�omm���shq��TI" ��co��
! yo���pane��� 
!��ty�le selec]t��H59��nD�~��onitor��48����tr��R�eliab���a�dinDiagnos"����2��2 ual Che�ck Safet�y UIF lg�\a��hance�d Rob Se�rv q ct\���lUser F�rU��DIF��E�xt. DIO 6��fiA d��wendr Err YL@��IF�r�ನ  �П�90��F�CTN Menu�Z v'��74� T�P In��fac�  SU (�G=�p��k E�xcn g�3��High-Sper wSki+�  sO��H9 � mmuni]c!�onsg�te�ur� ����V��y��conn���2��EN��Inc=rstru����5.fdKA�REL Cmd.� L?uaA� O~�Run-Ti� 'Env����K� ��u+%�s#�S/W���74��Licen�seT�  (A�u* ogBook�(Sy��m)��"�
MACR�Os,V/Off�se��ap��MH�� ����pfa5�M�echStop �Prot��� d��b i�Shif����j545�!x�r ��#��,���b ode Swiwtch��m\e�!�o4.�& pr�o�4��g��M?ulti-T7G����net.P{os Regi���z�P��t Fu9n���3 Rz1���Numx �����9�m�1�  Adju<j��1 J7�7�*� ����6tatu�q1EIKRD�Mtot��scove�� ��@By<- }uest1�$G�o� � U5\SNPX b"���<YA�"Libr��㈶�#�� �$~@h�p�d]0�Jts i?n VCCM����ĕ0�  �u!��2 �R�0�/I�08~��TMILIB�M� J92�@P�A�cc>�F�97�TgPTX�+�BRSQselZ0�M8 Rm��q%��692��Unexceptr �motnT  CcVV�P���KC�����+-��~K  I�I)�VSP CSXC�&.c�� e�"��� t�@We�w�AD Q�8bv9r nmen�@�KiP� a0y�0��pfGridAplay !� nh�@*��3R�1M-10iA�(B201 �`2�V"  F���sci�i�load��8�3 M��l����G�uar�d J85��0�mP'�L`���s�tuaPat�&]$C�yc���|0ori�_ x%Data'Pqu���ch�1���g`� j� RLJa�m�5���IMI �De-B(\A�cP"� #^0C  e�tkc^0assw�o%q�)650�Ap�U�Xnt��PvKen�CTqH�5�0�YELLOW� BO?Y��� Arc�0vis��C�h�WeldQci�al4Izt�Op�� ��gs�` 2@�a6��poG yRjcT1 NE�#HTf� xyWb��! �p��`gd`���p\� �=P��JPN ARCP*PR�A�� �OL�pSup̂fil�p��J�� n��cro�670�1�C~E�d��SS�pe.�tex�$ �P� �So7 t� ssa%gN5 <Q�BP:� 2�9 "0�QrtQCr��P�l0dpn������rpf�q�e�ppm�ascbin�4psyn�' pstx]08�HEL�NCL VIS �PKGS �Z@M�B &��B J8�@IPE GET_VAR FI?S_ (Uni� LU��OOL: ADD��@29.FD�TC4m���E�@DVp����`A�ТNO WT?WTEST �� ��!��c�FOR ^��ECT �a!� �ALSE ALA�`�CPMO-13�0��� b D: H�ANG FROM�g��2��R709� DRAM AV�AILCHECK�S 549��m�V�PCS SU֐L_IMCHK��P�0~x�FF POS� �F�� q8-12 CHARS��ER6�OGRA ���Z@AVEH�AME��.SV��Вאqn$��9�m "y��TRCv� SHA�DP�UPDAT �k�0��STATI���� MUCH ����TIMQ MOTN-003���@OBOGUI�DE DAUGH໱�b��@$tou�� �@C� �0��PA�TH�_�MOVE�T�� R64��V�MXPACK M�AY ASSERyTjS��CYCL`��TA��BE CO�R 71�1-�AN���RC OPTI�ONS  �`��A�PSH-1�`fi	x��2�SO��B��XO򝡞�_T��	�i�j�0j��du�byz �p wa��y�٠H�I������U�pb X?SPD TB/�F�_ \hchΤB0����END�CE�06�\Q�p{ sma'y n@�pk��L} ��traff#��	� ��~1fro�m sysvar/ scr�0R� ��Nd�DJU���H��!A��/��SET GERR�D�P7�����NDANT S�CREEN UNREA VM �P�D�D��PA���R~�IO JNN�0��FI��B��GRwOUNנD Y��Т٠�h�SVIP� 53 QS��DI�GIT VERS���ká�NEW�� �P06�@C�1IMCAG�ͱ���8� �DI`���pSSU�E�5��EPLAN� JON� DELL���157QאD��CALLI���Q��m���IPND}�IMG N9 PZ�{19��MNT/���ES ���`LocR Hol߀=��2�P�n� PG:��=�M��can����С�: 3D mE2view d X���ea1 �0b�po;f Ǡ"HCɰ��ANNOT AC�CESS M c�pie$Et.Qs �a� loMdFle�x)a:��w$qmo+ G�sA9�-'p~0̿�h0pa��eJ AUTO-�0��!�ipu@Т<ᡠIA�BLE+� 7�a F�PLN: L�p�l m� MD<�V�I�и�WIT H�OC�Jo~1Qu�i��"��N��US�B�@�Pt & r�emov���D�vAxis FT_7�PGɰCP:�O�S-144 � h� s 268QՐO�ST�p  CRA�SH DU��$P~��WORD.$��LOGIN�P��P�:	�0�046 i�ssueE�H�:� Slow st�c�`6�����z��IF�IMPR��SPOT:Wh4����N1STY��0V�MGR�b�N�CA�T��4oRRE�� �� 58�1��:N%�RTU!Pe -M .a�SE:�@pp���$AGpL��m@�all��*0a�OC�B WA���"3 �CNT0 T9DW�roO0alarm8�ˀm0d t�M��"0�2|� o�Z@O�ME<�� ��E%  ;#1-�SRE��M��st}0g   �  5KANJI~5no MNS@��INISITA7LIZ'� E�f�cwe��6@� dr�@� fp "��SC�II L�afai�ls w��SY�STE[�i�� � � Mq�1QGro8�m n�@vA�����&��n�0q��R�WRI OF L|k��� \ref"��
�up� de-r�ela�Qd 03�.�0SSchőb�etwe4�INDo ex ɰTPa�#DO� l� �ɰ�GigE�sope�rabil`p l�,��HcB��@]�lye�Q0cflxz�8Ð���OS {�����v4pfigi GL�A�$�c2�7H� wlap�0ASB� �If��g�2 l\�c�0�/�E�� �EXCE 㰁�P����i�� o0��G�d`]Ц�fq�l lsxt��EFal����#0�i�O�Y�n�CL�OS��SRNq1NT^�F�U��FqKP~�ANIO V7/�¥�1�{����DBa �0��ᴥ�ED��DET|�'� �b�F�NLINEb�B�UG�T���C"RL�IB��A��ABC? JARKY@���� rkey�`IL����PR��N��ITG+AR� D$�R �Er *�T��a�U�0��h�[�ZE V�� TASK p7.vr�P2" .�XfJ�srn�S谥d�IBP	c���B/��BUS��UNN�� j0-�{��cR�'���LOE�DIVS�CULs$cb����BW!��R~�W`�P�����IT(঱t�ʠ�OF��UNE�Xڠ+���p�FtE���SVEMG3`N�ML 505� D�*�CC_SAFE��P*� �ꐺ� PE�T��'P�`�F  �!���IR����c Ri S>� K��K��H GUNCHGz��S�MECH��IM��T*�%p6u���tPORY LE�AK�J���SP�EgD��2V 74\GRI��Q�g��oCTLN��TRe `@�_�p ���EN'�IN������$���r��T3)�i�STO��A�s�L��͐X	���q��Y� ��CTO2�J m��0F<�K����DU�S��O���3 9�J F��&���SSVGN�-1#I���RSRwQDAU�Cޱ� �T6��g��� 3�]���BR�KCTR/"� �q\�j5��_�Q�S�qI{NVJ0D ZO�P ݲ���s��г�Ui ɰx̒�a�DUAL�� J50e�x�RV�O117 AW�T�H!Hr%�N�247�%�52��|�&aol� ���R���at�Sd��cU���P,�LER��iԗQ0�ؖ  S!T���Md�Rǰt�_ \fosB�A�0@Np�c����{�U���ROP 2�b�pB>��ITP4M��b !AUt c0< � �plete�N@�� z1^qR635� (AccuCa�l2kA���I) �"�ǰ�1a\�Ps ��ǐ� bЧ0P������ig\cba?cul "A3p_ �1��ն���eta�ca��AT���PC��`�����_p�.�pc!Ɗ��:�cicrcB���5�tl��Bɵ�:�fm+�Ί��V�b�ɦ�r�upf�rm.����ⴊ�x�ed��Ί�~�ped�A�D �}b�ptl�ibB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆Ϙ���c�Ӳ�5�1j>�����tcȐ�Ϣ	�r����mm 1���T�sl^0��T�m�ѡ�#�rm3��u8b Y�q�std}��3pl;�&�ckv�=߆r�vf�䊰��9�v1i����ul�`�04fp�q �.f���� daq; i Da�ta Acqui+si��n�
��4T`��1�89���22 DMCM oRRS2Z�75���9 3 R710,�o59p5\?T "��1 (D�T� nk@���� ����E Ƒȵ��Ӹ��etdmm ��ER�����gE��1�q\mo?۳�=( G���[(

�2�` �! �@JMAC�RO��Skip/Offse:�a���V�4o9� &qR6C62���s�H��
 6Bq8����9~Z�43 J77� =6�J783�o `��n�"v�R5�IKCBq2 PT�LC�Zg R�3; (�s, �������03�	зJ���\sfmnmc? "MNMC�����ҹ�%mnf�FM�C"Ѻ0ª etm�cr� �8����� ,��D���   874\prdq>�,jF0���axi�sHProcess Axes e�wrol^PRA
��Dp� 56 J81�j�59� 56o6�� ���0w�690 998� [!IDV�1��2(x2��2ont �0�
����m2����?C��etis "ISD��9�� F/praxRAM�P�8 D��defB�,��G�isbasicHB�@޲{6�� W708�6��(�Acw:������D
�/,��AMOX�� ��DvE ��?;T��>Pi� RACFM';�]�!PAM�V �W�Ee�U�Q'
bU�75�.�ceN�e� nterfa�ce^�1' 5&!5�4�K��b(Dev am±�/�#���/<�Tazne`"DNEWE����btpdnui� �AI�_s2�d_rsono���bAs�fjN��bdv_arFvf�xhpz�}w��shkH9xstc��gAponlGzv{�ff��r���z��3{q'Td>pcOhampr;e�p� ^5977��	܀�4}0��mɁ�/�����l�f�!�pcchmp�]aMP&B�� �m�pev�����p�cs��YeS�� M/acro�OD��16Q!)*�:$�2U"_,x��Y�(PC ���$_;������o��J�g�egemQ@GEM�SW�~ZG�gesn�dy��OD�ndda��S��syT�Kɓ�Csu^Ҋ���n�m��<�L��  ���9:�p'ѳ޲��spotplusp���`P-�W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\f�eatu 0FEA�WD�oolo�s�rn'!2 p���a؝As3��tT.� (?N. A.)��!�e!�J# (j�,`��oBIB�oD -��.�n��k9�"K���u[-�_���p� "PSEqW����?wop "sEЅ� &�:�J������y�|� �O8��5��Rɺ��� ɰ[��X������ـ%�(
ҭ�q HL �0k�
�z�a!�B�Q�"(g�Q����� ]�'�.�����&���<�0!ҝ_�#��tpJ�H� ~Z��j�����y���� ��2��e������Z�� ��V��!%���=�]�p͂��^2�@iRV� Kon�QYq͋JF0B� 8ހ�`�	(^>�dQueue���X�\1�ʖ`�+F1tpv�tsn��N&��ftupJ0v �RDV�	�f��J1 Q���v��en��kvst�k��mp��btk�clrq���get����r��`kack�XZ��strŬ�%�st0l��~Z�np:!�`����q/�ڡ6!l��/Yr�mc�N+v�3�_� ����.�v�/\jF���� �`Q�΋ܒ�N50 (FRA��+�����fraparm���Ҁ�} 6�J6�43p:V�ELSE�
#�VAR $�SGSYSCFG�.$�`_UNITS 2�DG~°@�4�Jgfr��4A�@FRL-��0ͅ�3ې���L �0NE�:�=�?@�8 �v�9~Qx304��;�BPRSM~QA��5TX.$VNUM_OL��5��DJ�507��l� Functʂ"qwAP��琉�3 H�ƞ�kP	9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TP�PR���QA�prnaSV�ZS��AS8D�j510U�-�`cAr�`8 ��ʇ�DJR`�jYȑH  ��Q �PJ6�a2�1��48AA�VM 5�Q�b0 �lB�`TUP xb?J545 `b�`�616���0V�CAM 9�CwLIO b1�s5 ���`MSC8��
rP R`\s�STYL MNI�N�`J628Q  �`NREd�;@�`�SCH ��9pDCSU Mete�`�ORSR Ԃ�a0�4 kREIO�C �a5�`542�b9vpP<�nP�a�`�R�`7�`�M?ASK Ho�.r�7 �2�`OCO :��r3��p�b�p���r0X��a�`13\�mn�a39 HR�M"�q�q��L�CHK�uOPLG� B��a03 �q.��pHCR Ob�pC�pPosi�`fP6� is[rJ554��òpDSW�bM�D8�pqR�a37 }Rjr30 �1�s4 �R6�m7��52�r5 �2.�r7 1� P6����Regi�@T^�uFRDM�uSaq�%�4�`930�uS�NBA�uSHLB�̀\sf"pM�N{PI�SPVC�oJ520��TC�`�"MNрTMIL��IFV�PAC �W�pTPTXp6�.%�TELN N� Me�09m3�UECK�b�`U�FR�`��VCOR^��VIPLpq89q�SXC�S�`VVF��J�TP �q��Rw626l�u S�`�Gސ�2IGU�I�C��PGSt�\ŀH863�S�q������q34sŁ6�84���a�@b>�3� :B��1 T��9�6 .�+E�51 �y�q53�3�b1 ̛��b1 n�jr9 <���`VAT ߲�q�75 s�F��`�sA�WSM��`TOP u�ŀR52p���a�80 
�ށXY �q���0 ,b�`8855�QXрOLp}��"pE࠱tp�`LCyMD��ETSS�挀6 �V�CPEs oZ1�VRCd3�
�NLH�h��0011m2Ep��3 f��p���4 /165CR��6l���7PR���008 tB��9 o-200�`U0�p�F�1޲1 ��޲2 L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�J�?7 rbcfA�L��8\PC����"�32�m0u�n�K�Rٰn�5� 5EW
n�99 z��40 kB���3 ��6ݲ�`00�iB/��6�u��7�u��8 µ������s�U0�`�t �1 0�5\rb��2 E@���K���j���5˰��60��a�HУ`:Ł63�jAF�_���F�7 ڱ݀H�8�eHЋ�&�cU0��7�p���1u��8u��9 c73������D7� r��5t�97 ��E8U�1��2��1�)1:���h��1np�"���8(�U1��\pyl��,࿱v ��B�854��1V���D�-4��im��1�<����>br�3pr�48@pGPr�6 B����$�p��1����1�`͵�155ض157 �2��62�S����B��1b��2����1Π2"�2���B6`�1<c�4 7B�5i DR��8_�B/���187 uJ�8 ;06�90 rBn��1 (��202 /0EW,ѱ2^��2��90�U2�p�2��S2 b��4��2�a�"RB����9\�U�2�`w�l���4 6	0Mp��7������b�,s
5 ��3����<pB"9 3 ����l�`ڰR,:7 �2��V�2��5���2^H��a^9���qr�����n�5����5᥁""�8a�Ɂ}�5B���5����`UA���� ���86 �6 S�0�5�p�2�#�52�9 �2^�b1
P�5~�2`���&P*5��8��5��u�r!�5��ٵ544��%5��R�ąP nB^,z�c (�4���L���U5J�V�5��1�1^��%�����5 b21��gA���58W82� r�b��5N�E�589�0r� 1�95  �"������c8"a��|�L ���!J"5|6���^!�6��B�"8P�`#��+�8%�6B��AME�"1 iCN��622�Bu�6V���d� 4��84�`A�NRSP�e/S� C�5� �6� ��� \� �6� �V� 3�t��� T20CA�R��8� Hf� 1D�H�� AOE� ��� ,�|�� a�0\�� �!64K���ԓrA� �1 (M{-7�!/50T� [PM��P�Th:1�C��#Pe� �3�0� 5>`M75T"� �D�8p� �0Gc� u�4|��i1-710i�1B� Skd�7j�?6�:-HS,� �RN�@��UB�f�X�=m7C5sA*A6an���!X/CB�B2.6A �0 ;A�CIB�A�2�QF1�U�B2�21� /70�S� �4����Aj1��3p���r#0 B2\m*A@C��;bi"�i1K�u"A~AAU� imm7c7��ZA@HI�@�Df�A�D5*A��E� 0TkdR1�35�Q1�"*�@�Q�1�QC )P�1*A�5*A�EA�5XB�4>\77
B7=Q �D�2�Q$B�E7�C�D%/qAHEE�W7�_|` jz@� 2�0�Ejc�7�`�E"l7�@7@�A
1�E�V~`�W2%Qr�R9ї@0L_�#�����"A���b��H3s=rA/2�R5nR 4�74rNUQ1ZU�A�sw\m9
1M92L2��!F!^Y�ps� 2c1i��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHsXBSt62�q`s������ ��Pxq3530_*A3I)�2�db�u0�@� '4TX�m0�pa3i1A3s0Q25�c��st�r�VR1%e�q0
��j1 ��O2 �A�UEiy�@.�‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?P Q��qA!Pvs� 5	1 5aU���?PŅ���ဝQ9A6�zS*�7�qb5�1����Q��'00P(��V7]u�a itE1���ïp?7� �!?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ�޵y00\ry�"R�2BL�tN  ���� �1D�Aʑ2�qeR�5���_b�3�X]1m1l�cqP1�a�E�Q� 5�F����!5���@M-16Q�� f���r���Q�e� ��� PN�L�T_�1��i1��945�3��@�e�|�b1l>F1u*AY2�
�R8�Q����RJ�J13�D}T� 85
Qg� /0��*A!P�*A�Ð�d����2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt]1 ^u�ajrI�B����~`�|I�b��yI�\m�Qb�I�uz�A�c3Apa\9q� B6S��S��m���}�85`N�N�  �(M�� �f1���6����161j��5�s`�SC���U��A����5\se�t06c����10��y�h8��a6��6x��9r�2HS �� �Er���W@}�a��IlB���Y�ٖ�m�u �C����5�B��B��h`�F���X0���A :���C�M��AZ��@��4�6i����� e�O�-	���f1��F  �ᱦ�1F�Y	���GT6HL3��U66~`Ȗ��U�dU�9D20Lf0��Qv� ��fjq ��N������0v
� ���i	�	��72l�qQ2������� \�chngmove�.V��d���@2l_arf	�f ~��6������9C��Z���~���kr41@ S���0��V��t�����U�p7nu�qQ%�A]��V�1\"�Qn�BJ�2W� EM!5���)�#:��64��F�e50S �\��0�=�PV�� �e������E������m7shqQSH"U��)��9�!A���(���� �,���ॲTR11!��,�60e=��4F�����2��	 R-����������@�Ж��4���LS0R�)"�!lOA��Q�X) %!� 16�
U /��2�"2�E�9p���2>X� SA/i��'�
7F�H�@!B�0�� �D���5V��@2cV E��p��T��pt갖��1L~E�#�F�Q��9�E�#De/��RT��59���	�A�EiR���|����9\m20챃20��+�-u�19r4 �`�E1�=`O9`� �1"ae��O�2��_\$W}am41�4�3��/d1c_std ��1)�!�`_T��r~�_ 4\jdg�a �q�PJ%!~`-�r�+�bgB��#c300D�Y�5j�QpQb1�`bq��vB��v25�Up�����qm43�  �Q<W�"PsA��e ����t�i�P�W .��c�FX.�e4�kE14�44�~o6\j4�443sxj��r�j4up�� �\E19�h�PA�T�= :o�APf��coWol!\�2a��2A;_	2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a�:88J9X�l5�m�1a첚��*���(85�&�������P6���R,52&A����,fA9IfI50\u�z�OV
�v��}E�֖J���Y>� 16�r�C�Y��;��1��L ���Aq�&ŦP1��vB�)e�m�����1pĻ �1D�ʹ27��F�KAREL �Use S��FC�TN��� J970�FA+�� (�Q޵0�p%�)?�Vj9F?(��j�Rtk208 C"Km�6Q�y�j��iæPr�9�s#��v��krcfp�RCF�t3���Q��kcctme�!ME�g����^6�main�dV�� ��ru��kDº��c���o����J�dt��F �»�.vrT�f�����E%�!��\5�FRj73B�K����UER�HJ�O  �J�� (ڳF���F �q�Y�&T��p�F�z��19�tkvBr���V�Bh�9p�E�y�<�k�������;�v���"CT��f����)�
І ��)�V	�6���!� �qFF��1q���=��� ��O�?�$"���$���je���TCP A�ut�r�<520 �H5�J53E19�3��9��96�!8���9��	 �B574V��52�Je�(�� Se%!Y�����u���ma�Pqtool��ԕ������co�nrel�Ftro�l Reliab�le�RmvCU!��H51����� a�551e"�CNRE¹I�c�&���it�l\sfut?st "UTա��"X�\u��g@�i�D6Q]V0�B,Eѝ6A� �Q�)C���X���Yf�I�1|6s@6i��T6IU��vR��d�
$e%1��2�C58�E6��8�Pv�iV�4OFH58SOeJ� mnvBM6E~O58�I �0�E�#+@�&�F�0 ���F�P6a���)/++��</N)0\tr1x�����P ,��ɶ��rmaski�ms�k�aA���ky'd�h�	A	�P�sDisp_layIm�`v��~��J887 ("A��+Heůצprd�s��Iϩǅ�h�0p�l�2�R2��:�Gt�@��PRD�TɈ�r��C�@Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��Px^@�P�firmQ� ���Pp�2�=bk�6�r��3��6��tppl��PL���O�p<b�ac�q	��g1J�U�d0�J��gait_9e���Y�&��Q���	�S�hap��erat�ion�0��R6�7451j9(`sGen�ms�42-f�Ár�p�5����2�rsgl�E��p�G���qF�205p�5S���ՁN�retsap�BP�O��\s� "GC�R�ö? �qngda�G��V��st2axU��Aa]��b�ad�_�btpu�tl/�&�e���tp�libB_��=�2.p����5���cird��v�slp��x�hex��v�re?�Ɵx�gkey�v�pm���x�us$�6�gcr��F������[�q27�j92�v�ollismqSk�9O��>�� (pl.���t��p!o��29$Fo8���cg7no@�tptwcls` CLS�o�b�\�km�ai_
�!s>�v�o	�t�b��x�ӿ�E�H��6~�1enu501�[�m��utia|$c�almaUR��Ca�lMateT;R5	1%�i=1]@-��/V�� ��Z�� �fq1�9 "K9E�L����z2m�CLMTq��S#��et �LM�3!} �F�c�ns�pQ�c���c_mo4q��� ��c_e���F��su��ޏ �_ �x@�5�G�join�@i�j��oX���&cW0v	 ���N�ve��C�clm�&Ao# �|$�finde�0�STD ter� FiLANiG���R��
��8n3��z0Cen���r,������J��� �� ���K��Ú�=�К�_Ӛ��r� "FNDR�� 3��}f��tguid��`��N�."��J�tq��  �������������J����_������c���	m�Z��\fndr.��n#>
B2�p��Z�CP Ma�����38A��� c
��6� (���N�B ������� 2�$�	81��m_���"ex�z5�.Ӛ��c���bSа�ef�Q��	��RBT~;�OPTN � +#Q�*$�r*$��*$r *$%/s#C�d/.,P�/|0*ʲDPN���$���$*�Gr�$ko Exc�'IF�$�MASK�%93 {H5�%H558�$_548 H�$4-1��$��#1(�$�0 E�$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3��9j0"M�49�4 � ��4�4tp�sh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E�\���5�A�4��3a�dq\�5K979�":E�ajO l "�DQ^E^�3i�Dq� ��4ҲO ?R�? ��q�5��T��3rAq�O�Lst�5~��7�p�5��REJ#�2�@a�v^Eͱ�F���4��.��5y N� �2il�(in�4��31 aJH1�2Q4�251ݠ��4rmal� �3) �REo�Z_�æOx�����4��^F�?onor Tf��7_ja�UZҒ4l��5rmsAU�Kkg���4�$HCd\�fͲ�e�ڱ�4�REM���4y�ݱ"u@�RER593�2fO��47Z��5lity,�U��e"DGil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe�=$��^�
E��u�IAymptm�U��BU��vste�y\�3��me� b�DvI�[�Qu�:F�U�b�*_�
E,�su$��_ Er��oxx���4huse�E-�?�sn�������FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��� b���(��1�� �c��Y�R�� �>�P� ��W��������'��0ɵ�[��͂����  � ,�N@� �A��bumpšf��B*�Box%��7Aǰ�60�BBw���MC� u(6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`���)���\bbk968� "�4�ω�bb��9va69����etbŠ��X�����#ed	�F��u�f�& �sea"������'�\��,���b�ѽ"�o6�H�
�x�$�f���!y���Q[�!� tperr�f�d� TPl0o� R/ecov,��3D���R642 � 0���C@}s� N@��(NU�rro���yu2�r��  �
�  ����$$�CLe� �������������$~z�_DIGIT��.������ .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ oo$j��+c:PRODUCTM��0\PGSTKD��V&ohozf99���D���$F�EAT_INDE�X��xd���  
�`IL�ECOMP ;����#��`�cS�ETUP2 <��e�b�  �N �a�c_AP2�BCK 1=�i  �)wh0?{%&c����Q� xe%�I�m�� �8��\�n����!� ��ȏW��{��"��� F�Տj���w���/�ğ S���������B�T� �x������=�үa� �����,���P�߯t� �����9�ο�o�� ��(�:�ɿ^���� �ϸ�G���k� �ߡ� 6���Z�l��ϐ�ߴ� ��U���y����D� ��h��ߌ��-���Q� ��������@�R��� v����)�����_��� ��*��N��r� �7��m�@&�3\�i
pP� 2#p*.V1Rc�*��`� /��PC/|1/FR6:/"].��/+T�`�/ �/F%�/�,�`r/?��*.F�8?	�H#&?e<�/�?;STM �2�?�.K �?��=iPen�dant Panel�?;H�?@O�7�.O�?y?�O:GIF �O�O�5�OoO�O_:JPG _J_�56_�O�_�_�	PANE�L1.DT�_@�0�_�_�?O�_2�_�So�WAo�_o�o�Z3 qo�o�W�o�o�o)�Z4�o[�WI���
TPEINSO.XML��0�\���qCust�om Toolb�ar	��PAS�SWORDy�FRS:\L�� �%Passwo�rd Config���֏e�Ϗ�B 0���T�f�������� ��O��s������>� ͟b��[���'���K� �򯁯���:�L�ۯ p�����#�5�ʿY�� }��$ϳ�H�׿l�~� Ϣ�1�����g��ϋ�  ߯���V���z�	�s� ��?���c���
��.� ��R�d��߈���;� M���q������<��� `������%���I��� �����8����n ���!��W�{ "�F�j| �/�Se��/ �/T/�x//�/�/ =/�/a/�/?�/,?�/ P?�/�/�??�?9?�? �?o?O�?(O:O�?^O �?�O�O#O�OGO�OkO }O_�O6_�O/_l_�O �__�_�_U_�_y_o  o�_Do�_ho�_	o�o -o�oQo�o�o�o�o @R�ov��; �_���*��N� �G������7�̏ޏ m����&�8�Ǐ\�� ���!���E�ڟi�ӟ ���4�ßX�j����� ���įS��w�������B�#��$FIL�E_DGBCK �1=��/���� ( ��)
SUMMA�RY.DGL����MD:������Diag Sum�mary��Ϊ
C?ONSLOG������D�ӱCon�sole log�E�ͫ��MEMCHECK:�!ϯ����X�Memory� Data��ѧ��{)��HAD�OW�ϣϵ�J����Shadow C?hangesM�'��-��)	FTAP7Ϥ�3ߨ���Z��mment TB�D��ѧ0=4)�ETHERNET��������T�ӱE�thernet �\�figurat�ionU�ؠ��DCSVRF�߽߫������%�� ve�rify all���'�1PY���DIFF�����[����%��diff]������1R�9�K���� ���X=��CHGD������c��r�����2ZAS� ��GD����k��z��FY�3bI[� �/"GD����s/����/*&UPDATES.� ��/��FRS:\��/�-ԱUpda�tes List��/��PSRBWLOD.CM(?���"�<?�/Y�PS_ROBOWEL��̯�? �?��?&�O-O�?QO �?uOOnO�O:O�O^O �O_�O)_�OM___�O �__�_�_H_�_l_o �_�_7o�_[o�_lo�o  o�oDo�o�ozo�o 3E�oi�o�� �R�v���A� �e�w����*���я `���������O�ޏ s������8�͟\�� ���'���K�]�쟁� ���4���ۯj����� �5�įY��}���� ��B�׿�x�Ϝ�1� ��*�g�����Ϝ��� P���t�	�ߪ�?��� c�u�ߙ�(߽�L߶� �߂���(�M���q�  ���6���Z���� ��%���I���B������2�����h�����$FILE_� P�R� ��������M�DONLY 1=�.�� 
 � ��q��������� �~%�I�m �2��h� �!/�./W/�{/
/ �/�/@/�/d/�/?�/ /?�/S?e?�/�??�? <?�?�?r?O�?+O=O �?aO�?�O�O&O�OJO �O�O�O_�O9_�OF_�o_
VISBCK�L6[*.VD�v_�_.PFR:\��_�^.PVis�ion VD file�_�O4oFo\_ joT_�oo�o�oSo�o wo�oB�of�o �+����� ��+�P��t���� ��9�Ώ]�򏁏��(� ��L�^�������5� ��ܟk� ���$�6�ş�Z��~�����
M�R_GRP 1>�.L��C4 w B���	 W������*u����RHB ���2 ��� ��� ���B� ����Z�l���C���D�ি����Ŀ��K���L5ȦJ����F�5UT?��Q�n�����ֿ G,�F�I�/E���.���9:�]�@��'�A&�#�A�f�?�f��A~��r��E�� F@ ��������J��NJ�k�H9�H�u��F!��IP�s�?����(��9�<9��896C'�6<,6\b� �+�&�(�a�L߅�X���A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�P=��P��K���ܿ� �B���/ ��@�33�:��.�g&�@U�UU�U��q	>u?.�?!rX���	�-=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7��:����D�@ ?D�� Cϥ��C������Q�,/� �����/M��/q��/ �/�/�??:?%?^? p?[?�??�?�?�?�?  O�?�?6O!OZOEO~O iO�O�O�O�OW�ߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������0�[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U�� 
//./�v���/ ���/�/�/�/�/� !?3?E?W?i?�/?�? �?�?�?�?�?��� AO�?eO�/�O�O�O�O �?�O�O__+_NO�O J_s_�_�_�_�_
OO .OoB_'ovOKo]ooo �oP_>o�o�o�o�oo �o5GYk}�_ �_�_��8o�� 1�C�U�$y������� �ӏf���	��-�?� ����Ə���ϟ �����;�M�_� q���.�(���˯ݯ� �P�b�t�����m��� ������ǿٿ����� !�3�E�h��{ύϟ� �����$�6�H�J�/� ~�S�e�w߉ߛ�jϿ� �������*߬�=�O��a�s��YT_ER�R J5
���P�DUSIZ  j��^J����>��?WRD ?t���  guest}��%�7��I�[�m�$SCDMNGRP 2Ktw�������V$�K�� 	�P01.14 8~��   y�����B   � ;����� ����������
 �������?�����~����C.gR|����  i  ��  
��������� +�������
���l �.r���"�l��� m
d����|��_GROU��]L�� �	�����07EQUPD'  	պ�J��TYa ����T�TP_AUTH �1M�� <!iPendany���6�Y!K?AREL:*��
-KC///A/ �VISION �SETT�/v/� "�/�/�/#�/�/
? ?Q?(?:?�?^?p>�CTRL N�����5�
�.?FFF9E3�?��FRS:DEF�AULT�<F�ANUC Web Server�:
�����<kO}O�O�O�O�O��WR_C�ONFIG OΡ� �?��ID�L_CPU_PC�@�B��7P�;BHUMIN(\��~<TGNR_IO�������PNPT_�SIM_DOmV�w[TPMODNT�OLmV �]_PR�TY�X7RTOLN/K 1P����_�o!o3oEoWoio�RMASTElP��R��O_CFG�o�iU�O��o�bCYCL�E�o�d@_ASG� 1Q����
  ko,>Pbt�� �������sk.�bNUM����K@�`IPCH�o��`RTRY_CN@xoR��bSCRN����Q��� �b�`�b�R���Տ��$�J23_DSP_�EN	����OBPROC�U�i�JOGP1SY@~��8�?�!��T�!�?*�POSR�E�zVKANJI�_�`��o_�� ��T��L�6͕����CL�_LGP<�_���EY�LOGGIN�`���LANG?UAGE YF7R�D w���LG���U�?⧈�xR� �����=P��'0��$ N�MC:\RSCH�\00\��LN_DISP V��`
��������OC�R�.RDzVTA{�OGBOOK W
{���i��ii��X �����ǿٿ����1�"��6	h������e�?�G_BU_FF 1X�]��2	աϸ����� ������!�N�E�W� ��{ߍߺ߱�����������J���DC�S Zr� =����^�+�ZE���������a�IO 1[�
{ ُ!� � !�1�C�U�i�y����� ����������	- AQcu��������EfPTM  �d�2/ASe w������� //+/=/O/a/s/�/8�/��SEV���]�TYP`�/??y͒�RS@�"��×�FL 1\
������?�?�?`�?�?�?�?/?TP6���">�NGN�AM�ե�U`�UP�S��GI}�𑪅�mA_LOAD�G� %�%DF_MOTN���O�@�MAXUALRM <��J��@sA�Q����QWS ��@C �]m�@-_���MP2�7�^
{� ر�	�!�P�+ʠ�;_/��R1r�W�_�WU�W�_ ��R	o�_o?o"oco Noso�o�o�o�o�o�o �o�o;&Kq\ �x������ �#�I�4�m�P���|� ��Ǐ���֏��!�� E�(�i�T�f�����ß ��ӟ���� �A�,� >�w�Z�������ѯ�� ��د���O�2�s� ^�������Ϳ���ܿ��'��BD_LDX�DISAX@	��M�EMO_APR@E� ?�+
  � *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT ��Q�c�Ϝ߇��ߧ� ����w����>�)�b� t�[����{����� �����:���I�[�/� �����������o��� ��6!ZlS� �s����2 �AS'�w�� ��g��.//R/�d/�_MSTR �`�-w%SCD 1am͠L/�/H/�/ �/?�/2??/?h?S? �?w?�?�?�?�?�?
O �?.OORO=OvOaO�O �O�O�O�O�O�O__ <_'_L_r_]_�_�_�_ �_�_�_o�_�_8o#o \oGo�oko�o�o�o�o �o�o�o"F1j Ug������ ���B�-�f�Q����u�����ҏh/MKC_FG b�-�~�"LTARM_���cL�� �σQ�N�<�METsPUI�ǂ���)�NDSP_CMN�Th���|�  	d�.��ς�ҟܔ�|�POSCF�����PSTOL 1�e'�4@�<#�
5�́5�E�S�1�S� U�g�������߯��ӯ ���	�K�-�?���c��u�����|�SING_CHK  ��^;�ODAQ,�f���Ç��DEV }	L�	MC:!̟HSIZEh��-���TASK %�6�%$123456789 �Ϡ��TRIG 1g�+ l6�%���ǃ`�����8�p�YP[�� ��EM_INF� 1h3� �`)AT&�FV0E0"ߙ�)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ������H�����A���AI�q�,��|���� ���ߵ�����J� ��n������W����� ������"����X� �/����e��� ���0�T;x� =�as��/� ,/c=/b/�/A/�/ �/�/�/��?�� �^?p?#/�?�/�?s? }/�?�?O�?6OHO�/ lO?1?C?U?�Oy?�O �O3O _�?D_�OU_z_�a_�_�ONITO�R��G ?5�  � 	EXEC�1Ƀ�R2�X3�X4��X5�X���V7�X8
�X9Ƀ�RhBLd�R Ld�RLd�RLd
bLdb Ld"bLd.bLd:bLdFb�Lc2Sh2_h2kh2�wh2�h2�h2�h2��h2�h2�h3Sh3�_h3�R�R_GRP_SV 1in����(ͅ�
�3w�8��r�ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A��W�@<�P�R�
h�B�b�A��j���a��:��Dzۀ���߹�����j���( �� -��C���'�7��&���q�Y������ �?�ff ���gy ������q+q��
>N+�  PƱj�(�� ��7	���|�/?����xZ�p�<
6b<߈�;܍�<�ê�<� <�&Jσ�AI�ɳ+����?fff?I�?y&�k�@�.��J<?�`� q�.�˴fɺ�/�� 5/����j/U/�/y/ �/�/�/�/�/?�/0?q��F�?l??��?/�?+)�?�?�E��� E�I�G+� F��?)O�?�9O_OJO�OnO�Of�BL޳B�?_h�.��O �O��%_�OL_�?m_�?��__�_�_�_�_�
��h�Îg>��_Co�_goRodo�oF�GA�ds�q�C�op�o�o|�����$]Hq���D��fpC���pCHm�ZZ7t���6q�q�����N'�3A�A��AR1AO�^?�$�?�K��0±
=ç>�����3�W
�=�#�W��e���9�����{����<���(�B�u�����=B0�������	L��H��F�G���G���H�U`E���C�+����I#�I���HD�F���E��RC�j=���
I��@�H�!H�( E<YD0q �$��H�3�l�W��� {��������՟��� 2��V�A�z���w��� ��ԯ�������� R�=�v�a��������� ���߿��<�'�`� Kτ�oρϺϥ����� ���&��J�\�G߀� kߤߏ��߳������� "��F�1�j�U��y� ������������0�@�T�?�Q����(�1g��3/E�����5������q�3�8�����q4�Mgs&IB�+2D�a���{�^^	���P���uP2P7Q4_A��M0bt��R����X��/   �/ �b/P/�/t/�/ *a@)_3/�/�/�%1a�?�/?;?M?_?q?  �?�/�?�?�?�?�O 2 F�$N�vGb�/�A��@X�a�`�qC��C@�o��O2���OF� �DzH@�� F�P D���O�O�ys<O!_3_E_W_i_~s?���@@pZ�.t22!:2~
 p_�_ �_�_	oo-o?oQoco�uo�o�o�o�o��Q ���+��1���$MSKCFMA�P  �5� �6�Q�Q"~��cONREL  �
q3�bE�XCFENB?w
8s1uXqFNC_Qt�JOGOVLIM�?wdIpMrd�bKE�Y?w�u�bRU�N�|�u�bSFSPDTY�avJu�3sSIGN?QtTO1MOT�Nq�b�_CE_GRP [1p�5s\r� ��j�����T��⏙� �����<��`��U� ��M���̟��🧟� &�ݟJ��C���7��� ����گ�������4��V�`TCOM_C_FG 1q}�V�p�����
P�_AR�C_\r
jyUA�P_CPL��ntN�OCHECK ?={ 	r ��1�C�U�g�yϋ� �ϯ���������	���({NO_WAITc_L�	uM�NTX��r{�[m�_E�RRY�2sy3�� &�������r��c� ��T_MO���t��, K��$�k�3�PARAM:��u{��V[ﰽ�!�u?�� =9@3�45678901 ��&���E�W�3�c������{������� �����=�UM_RSPACE ��Vv��$ODR�DSP���jxOF�FSET_CAR9Tܿ�DIS���PEN_FILE�� �q��c֮�OPT?ION_IO���PWORK v_�ms �P(��R�Q
�j.j	 ���Hj&6$� R�G_DSBL  ��5Js�\��R�IENTTO>p�9!C��PqfA� UT_SIM_D�
r�b� V� LCT ww�bc��|U)+$_PEXE�d&RATp �vju�p���2X�j)TUX�)TX�##X d-�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O�H2�/oO�O�O�O�O@�O�O�O�O_]�<^O ;_M___q_�_�_�_�_��_�_�_o���X�O�U[�o(��(����$o�,� ��IpB` @oD�  Ua?�[cbAa?��]a]�DWcxUa쪋l;�	lmb��`�x�J�`�����a�< ��`�� ��b, H(���H3k7HSM5�G�22G��ޏGp
��
�!���'|, CR�>��>q�GsuaT�o3���  �4sp�Bpyr  ]o�*SB_����j]���t�q� ���rna �,���_6  ��PUQ�|N�M��,k�!�	'� �� ��I� ��  ��%�=���ͭ���ba	����I  �n @��~���p�"���� �N	 W��  '!o�:q�pC	 C�@@sBq�|�:�� m�
�!�h@ߐ�n����Z��B	 �A���p�# �-�qbz�P���t�_�������( �� -��恊�n�ڥ[A]ё��b4�'!��(p �?�ff� ��
�����OZ�R��8��z���>΁  Pia��(�ವ@���ک�a�c�dF#?����x����<
6b�<߈;܍��<�ê<� �<�&�o&�)�A��lcΐI�*�?ff�f?�?&c���@��.uJ<?�`��Yђ^�nd ��]e��[g��Gǡd<� ���1��U�@�y�d� �߯ߚ����߼�	��߀-������&��"�E��� E��G+� Fþ������ �����&��J�5��
bB��AT�8�ђ�� 0�6���>���J�n�7��[m�0���h��1��>�M�I
�@F��A�[��C-�)��?�ؠ�� /�YĒ��0Jp��vav`CH/�������}!@I��Y�'�3A�A��AR1AO��^?�$�?�����±
=ç�>����3�W�
=�#����+e��ܒ�����{�����<���.(�B�u���=B0��?����	�*�H�F�G����G��H�U`�E���C�+��-I#�I���HD�F���E��RC�j�=U>
I���@H�!H�(� E<YD0 /�?�?�?�?�?O�? 3OOWOBOTO�OxO�O �O�O�O�O�O_/__ S_>_w_b_�_�_�_�_ �_�_�_oo=o(oao Lo�o�o�o�o�o�o�o �o'$]H� l������� #��G�2�k�V���z� ��ŏ���ԏ���1� �U�g�R���v������ӟ�������-��(ε�������<a����Q�c�,!3�8�}���,!�4Mgs����ɢI�B+կ篴a���{���A�/��e�S���w��P!�P�������7��ӯ�ϑ�R9�Kτϰoχϓϥ�  ��� �χ����)��M��ʀ�������{߉ߛ� ��ߒߤ�������  )�G�q�_�����2 F��$�&Gb���n�[ZjM!C�s�@�j/�A�S���F�� Dz��� F?�P D��W����)������������x?���@@*
9�E�E��uE��
  v������� *<N`�*P� ���˨�1���$PARAM_MENU ?-���  �DEFPU�LSEl	WAITTMOUT��RCV� �SHELL_WR�K.$CUR_S�TYL�,OsPT�/PTB./�("C�R_DECSN���,y/�/�/ �/�/�/�/?	??-?�V?Q?c?u?�?�US�E_PROG �%�%�?�?�3CC�R�����7_H�OST !�!�44O�:T̰�?PC�O)ARC�O�;_T�IME�XB�  ��GDEBUG�V@��3GINP_�FLMSK�O�IT�`��O�EPGAP 2�L��#[CH�O�H�TYPE��� �?�?�_�_�_�_�_o o'o9obo]ooo�o�o �o�o�o�o�o�o: 5GY�}��� ������1�Z���EWORD ?	�7]	RS`�	/PNS�$��sJOE!>�TEs@�WVTRACECToL 1x-��W ��Ӱ�|�ɆDT Qy-����D � ��,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�T�(�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_j��_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ�_ ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������//�"#�$PGTRA�CELEN  �#!  ���" �8&_UP z���g!�o S!h 8!_�CFG {g%Q#"!x!�$J �"� |"DEFSPD� |�,!!J ��8 IN TRLW }�-" 8�(�IPE_CONF�I� ~g%��g!�$�$�"8 L�ID�#�-74G�RP 1�7Q!��#!A ����&ff"!A+33�D�� D]� ?CÀ A@+6�!�" d�$�9�9*1*0?� 	 +9�-+6�? ´	C�?�;B@3AO�?OIO3O�mO"!>�T?��
5�O�O�N�O =��=#�
�O _�O_J_5_n_Y_�O�}_�_y_�_�_�_  #Dzco" 
oBo �_Roxoco�o�o�o�o �o�o�o>)b�M��;
V7.10beta1�$�  A�E}�rӻ�A " ޼p?!G��q>˙��r��0�q̽ͻqBQ��qAA\�p�q�4�q�p�"�BȔ2�D�V�h�Bw��p�?�?)2{ ȏw�׏���4�� 1�j�U���y�����֟ ������0��T�?� x�c�������ү���� !o�,�ۯP�;�M��� q�����ο���ݿ� (��L�7�p�+9��sF@ �ɣͷϥ� g%������+�!6I� [߆������ߵߠ��� ������!��E�0�B� {�f���������� ���A�,�e�P��� t���������� ��=(aL^�� �����'9 $]�Ϛ��ϖ��� ����/<�5/`�r� �ߖߏ/>�/�/�/�/ �/?�/1??U?@?R? �?v?�?�?�?�?�?�? O-OOQO<OuO`O�O �O�O�O���O_�O)_ _M_8_q_\_n_�_�_ �_�_�_�_o�_7oIo t���o�o���o �o�o(/!L/^/p/�/ {*o������ ���A�,�e�P�b� ���������Ώ�� +�=�(�a�L���p��� ���Oߟ񟠟� �9� $�]�H���l�~����� ۯƯ���#�No`oro �on��o�o�o�oԿ ���8J\ng�� ��vϯϚ�������	� ��-��Q�<�u�`�r� �ߖ��ߺ������� ;�M�8�q�\������ ��z������%��I� 4�m�X���|������� ����:�L�^���Z ����������� $�6�H�Swb �������/ /=/(/a/L/�/p/�/ �/�/�/�/?�/'?? K?]?H?�?��?�?f? �?�?�?O�?5O OYO DO}OhO�O�O�O�O�O �O&8J4_F_�� ��_�_��_�_" 4-o�O*ocoNo�oro �o�o�o�o�o�o) M8q\��� ������7�"� [�m��?����R�Ǐ�� �֏�!��E�0�i� T���x��������_ $_V_ �2�l_~_�_������R�$PLID�_KNOW_M � �T������SV �v�U͠�U��
��.�ǟR�=��O�����mӣM_G�RP 1��!`0*u��T@ٰo�ҵ�
���Pзj�� `���!�J�_�W�i� {ύϟϱ��������Ϭ߱�MR�����T��s�w� s��ߠ� �߯߅��ߩ߻����� A���'����� ����������=�� �#���������}���ء��S��ST��1 �1��U# ���0�_ A .��, >Pb����� ���3(iL ^p������2*���<-/3/)/;/M/A4f/x/�/�/5�/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?MA/D  d#`�PARNUM � w�%OS+CH?J ME
�G`A8�Iͣ�EUPD`OrE�
a�OT_CMPa_��B@�P@'˥~TER_CHK'U���˪?R$_6[RqSl�¯��_MOA@�_�U_�_RE_RES_G ��>� oo8o+o\oOo�oso �o�o�o�o�o�o�o�W �\�_%�Ue  Baf�S� ��� �S0����SR0� �#��S�0>�]�b��S��0}������RV 1񈟥��rB@c]���t�(@c\�����D@c[��$���RTHR_ICNRl�DA��˥d,�oMASS9� ZM��MN8�k�MON_�QUEUE ����˦��x� RDN�PUbQN{�P[��E�ND���_ڙEXE�ڕ�@BE�ʟ��OPTIOǗ�[���PROGRAM %��%��ۏ�O~��TASK_IAD�0�OCFG ��tO��ŠDATA����Ϋ@��2 7�>�P�b�t���,��� ��ɿۿ�����#�5ϼG���INFOUӌ�������ϭϿ��� ������+�=�O�a� s߅ߗߩ߻�������h�^�jč� y�ġ?PDIT ��ίc���WERFL�
��
RGADJ7 �n�A�����?����@���IOR�ITY{�QV���M�PDSPH�����U�z����OTOE�y�1�R� (!AF4�E�P]���?!tcph����!ud��!�icm��ݏ6�X�Y_ȡ�R��ۡ)� *+/ ۠�W:F� j�������%7[B�*���PORT#�BC�۠����_CARTREP
�R� �SKSTAz��ZS�SAV���n�	�2500H863����r�$!�R�
���q�n�}/�/��'� URGE�Bl��rYWF� DO{��rUVWV��$�A�W�RUP_DELA�Y �R��$R_'HOTk��%O]?��$R_NORMA�Lk�L?�?p6SEM�I?�?�?3AQSKkIP!�n�l#x 	1/+O+ ORO dOvO9Hn��O�G�O�O �O�O�O_�O_D_V_ h_._�_z_�_�_�_�_ �_
o�_.o@oRoovo do�o�o�o�o�o�o�o *<Lr`����n��$RCV�TM�����pDkCR!�LЈq�Cl�fC���C��>?�A��>:��<l���4M�b�����O
�n��������{��4Oi��O <
�6b<߈;����>u.�??!<�&{�b� ˏݏ��8�����,� >�P�b�t��������� Ο���ݟ��:�%� 7�p�S������ʯܯ � ��$�6�H�Z�l� ~�������ƿ���տ ���2�D�'�h�zϽ� �ϰ���������
�� .�@�R�d�Oψߚ߅� �ߩ���������<� N��r������� ������&�8�#�\� G�����}��������� ��S�4FXj| ������� ��0T?x�u ����'//,/ >/P/b/t/�/�/�/�/ �/�/�?�/(??L? 7?p?�?e?�?�?��? �? OO$O6OHOZOlO ~O�O�O�?�?�O�O�O �O __D_V_9_z_�_ �?�_�_�_�_�_
oo�.o@oRodovo�X�qG�N_ATC 1��� AT�&FV0E0�k�ATDP/6/�9/2/9�hA�TA�n,A�T%G1%B96}0�i+++�o�,�aH,�qIO�_TYPE  �u�sn_�oREFPOS1 1�P{� x�o�X h_�d_����� K�6�o�
���.���R�x���{{2 1�P{���؏V�ԏz����q3 1��$�6��p��ٟ���S4 1�����˟���n�|��%�S5 1�<��N�`�����<���S6 1�ѯ���/�𭿘�ѿO�S7 1�f�x���ĿB�-�f�>�S8 1������Y�������y�SM�ASK 1�P � 
9�G��XNO�M���a~߈ӁqMOTE  h�~t��_CFG �������рrPL_RA�NG�ћQ��POW_ER ��e����SM_DRYP_RG %i�%���J��TART ��
�X�UME_P�RO'�9��~t_E�XEC_ENB � �e��GSPD�������c��TDB����RM��MT�_!�T���`O�BOT_NAME� i���iO�B_ORD_NU�M ?
�\q�H863  a�T��������b�PC_TIMEO�UT�� x�`S2�32��1��k �LTEACH PENDAN ��ǅ�}���`�Maintena�nce ConsțR}�m
"{�dKCL/Cg��Z ���n� No Use}�	���*NPO��х����(CH_�L�������	��mMAVAILȰ�{��ՙ�SPACE1 2��| d��(>���&���p��M,8�?�ep/eT/ �/�/�/�/�W//,/ >/�/b/�/v?�?Z?�/ �?�9�e�a�=??,? >?�?b?�?vO�OZO�?��O�O�Os�2� /O*O<O�O`O�O�_��_u_�_�_�_�_[3 _#_5_G_Y_o}_�_ �o�o�o�o�o[4.o@oRodovo$�o �o����"�	�7�[5K]o��A� ���	�̏�?�&�T�[6h�z������� ^�ԏ���&��;�\�C�q�[7�������� ͟{���"�C��X�y�`���[8����Ư دꯘ��0�?�`�#��uϖ�}ϫ�[G ��i� �ϋ
G� ����$�6� H�Z�l�~ߐ��8 ǳ�@����߈��d(� ��M�_�q���� ��������?���2� %�7�e�w��������� �����������!�R E�W�����������?Q; `�� @0�@�ߖrz	�V_ �����
/L/^/ |/2/d/�/�/�/�/�/ �/?�/�/�/*?l?~? �?R?�?�?�?�?�?�?�?2O�?
��O[�_MODE  ��˝IS ���vO,*ϲ�O-_���	M_v_#dCWO�RK_AD�M�{P%aR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/$��:	d/JaR��WY��^���^R�^	r  P��� �  8��P�	�D��GYk}�� ������Qp/@/R//)P;�o\T��Q�pg-�t�_�DiKT��[  � lv%������/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OWW�#�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_olO~O d+No`oro�o�o�o�o �o�o�o&8J \n������u�  0�"0g�/� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q�����$o��˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�����Do ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������w
�  58�J�\�n߀� �ߜկ���������	� �-�?�Q�c�u������ ��-�� ��� �2�D�V�h�z���������������v���& ���%	12345�678�" 	�
�/� `r�������� (:L^p�� ����� //$/ 6/H/Z/l/~/��/�/ �/�/�/�/? ?2?D? V?h?�/�?�?�?�?�? �?�?
OO.O@Oo?dO vO�O�O�O�O�O�O�O __*_YON_`_r_�_ �_�_�_�_�_�_oo C_8oJo\ono�o�o�o �o�o�o�oo"4 FXj|���������	��s�3�E�W�{�Cz � Bp��   ��2���z�$S�CR_GRP 1��(�U8(�\�x^ @�  �	!�	 ׃���"� $� ��-��+��R�nw����D~������#����O����M-10iA 78909905 Ŗ~5 M61C >P4��Jׁ
� ���0�����#�1�	"�z�������4¯Ҭ ���c� ��O�8�J��� ����!�����ֿ��B�y�������r��A��$�  @���<� �R�?��d���H�y�u�O���F@ F�`�§�ʿ�϶� ������%��I�4�m� �<�l߃ߕߧ߹�B���\����1�� U�@�R��v����� �������;���*<=�
F���?�d�<��>m���@��:��� B����ЗЙ���EL_D�EFAULT  ������B�MIPOWERFL  �x$1 WFDO� $��ERVE�NT 1������"�pL!D?UM_EIP��8���j!AF_I�NE �=�!FIT���!���4 ��[!�RPC_MAIN�\>�J�nVI�Sw=���!�TP�PU��	d��?/!
PMON?_PROXY@/�Ae./�/"Y/�fz/��/!RDM_S�RV�/�	g�/#?!#R C?�h?o?K!
pM�/�i^?��?!RLSYN�C�?8�8�?O!�ROS�.L�4 �?SO"wO�#DOVO�O �O�O�O�O_�O1_�O U__._@_�_d_v_�_ �_�_�_o�_?ooco�iICE_KL �?%y (%SVCPRG1ho 8��e���o�m3�o�o"�`4 �`5(-"�`6PU�`7x}��`���l9��{ �d:?��a�o��a�o E��a�om��a���a B���aj叟a�� �a�5��a�]��a� ���a3����a[�՟�a �����a��%��aӏM� �a��u��a#����aK� ů�as���a��mob �`�o�`8�}�w����� ��ɿ���ؿ���5� G�2�k�VϏ�zϳϞ� ���������1��U� @�y�dߝ߯ߚ��߾� ������?�*�Q�u� `���������� ��;�&�_�J���n������������sj_�DEV y	��MC:Pϻ_OUT"�,REC 1q�Z� d  / 	 	�������
� �PJ�%6 (�&�[w֍,�*  �T - �- �A�- c|�P�� ���//B/0/f/ x/Z/�/�/�/�/�/�/ �/?�/?P?>?t?b? �?�?�?�?�?�?�?O OOLO:OpO�OdO�O �O�O�O�O�O�O$__ H_6_X_~_l_�_�_�_ �_�_�_�_ ooDo2o Tozo\o�o�o�o�o�o �o�o.R@v d����},� ���4�"�X�F�|� ��p�����֏ď�� ��0��@�f�T���x� ����ҟ�Ɵ���,� �<�b�P���h�z��� ���ί��(�:�� ^�L�n�p�������ܿ �п� �6�$�Z�H� jϐ�rϴϢ������� ���2�D�&�h�Vߌ� z߰ߞ����������� 
�@�.�d�R��ZjoV 1�w P��m��	>  � ��
T�YPEVFZN_CFG ��'d7�?GRP 1�A�c/ ,B� A� �D;� B����  B4R�B21HELL�:�(
� �X����%RSR ����E0iT� x�������/Sew�  ��%w��(���#��������2#�d�����HK 1��� �k/f/x/ �/�/�/�/�/�/�/? ?C?>?P?b?�?�?�?��?��OMM �����?��FTOV_�ENB ���+�HO�W_REG_UI�O��IMWAITrB�JKOUT;F���LITIM;E;���OVAL[OMC_UNITC�F+��MON_ALIA�S ?e�9 ( he��_&_8_J_ \_��_�_�_�_�_j_ �_�_oo+o�_Ooao so�o�oBo�o�o�o�o �o'9K]n ����t��� #�5��Y�k�}����� L�ŏ׏������1� C�U�g���������� ӟ~���	��-�?�� c�u�������V�ϯ� �����;�M�_�q� �������˿ݿ��� �%�7�I���m�ϑ� �ϵ�`�������ߺ� 3�E�W�i�{�&ߟ߱� �����ߒ���/�A� S���w����X�� ��������=�O�a� s���0����������� ��'9K]� ���b��� #�GYk}�: ������/1/ C/U/ /f/�/�/�/�/ l/�/�/	??-?�/Q? c?u?�?�?D?�?�?�? �?O�?)O;OMO_O
O �O�O�O�O�OvO�O_�_%_7_�C�$SM�ON_DEFPR�O ����`Q �*SYSTEM*�  d=OURECALL ?}`Y� ( �}4c�opy md:p�rgstate.�dg virt:�\temp\=>�192.168.�4�P46:302�0 0>_�_�_o}�3�Uconslo	g�_�_ �_eowo�oiio�_<oNo�o�o��f2�Uerrall.ls�o�n�o�ew�`9�Rfr�s:orderf�il.dat1umpback<Nt�����j0�Tb:*.*�� �b�t����c6��x9�P8144 W������.��*.d��ƎϏ�`�r���e
xyz=r�` 61 +�=� O�����e���� ӑ��ҟc�u����� 5�͇ٯ����"����̈ѯb�t���c4x��:\)���;�S�U�����
� }5��a ����H�ؿi�{ώ��� ��@�V��������� B���e�w߉ߜ�/�<� ҿ�����ϫ߽�P� a�s��Ϫ�3����� ����(���L�]�o� ���ߦ�9��������� �$��H�Yk}�� ��+=O���>)�6788 �� cu����5�6� ���"��5�b/�t/�/�����8976 W/�/�/�/��/ �)�/`?r?�?���;? M?�?�?O'�4�? �?cOuO�O��5/�' �O�O�O/"/�O�(�O b_t_�_����:DV_��_�_o�_�_6  �_goyo�o�O�O9_T_ �o�o	_�o@_�oc u��_-o?o�_�� �o��No_�q��� �o�o1�oݏ���&��J[�m������$SNPX_AS�G 1�������� P� 0 '%�R[1]@1.1,����?���%֟� �&�	��\�?�f��� u��������ϯ��"� �F�)�;�|�_����� ��ֿ��˿���B� %�f�I�[Ϝ�Ϧ��� ��������,��6�b� E߆�i�{߼ߟ����� ������L�/�V�� e���������� ��6��+�l�O�v��� ������������2 V9K�o�� �����&R 5vYk���� �/��<//F/r/ U/�/y/�/�/�/�/? �/&?	??\???f?�? u?�?�?�?�?�?�?"O OFO)O;O|O_O�O�O �O�O�O�O_�O_B_ %_f_I_[_�__�_�_ �_�_�_�_,oo6obo Eo�oio{o�o�o�o�o �o�oL/V� e������� �6��+�l�O�v��������PARAM ������ W�	��P�����OFT_KB_CFG  ������PIN_SI/M  ���C��U�g�����RVQS�TP_DSB,��򂣟����SR ��/�� &  �ULTIROBO�TTASK������TOP_ON_�ERR  ����PTN z/�@�A	��RING_PRM�� ��VDT_?GRP 1�ˉ�  	�������� ����Я�����*� Q�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߣߠ߲��������� ��0�B�i�f�x�� ������������/� ,�>�P�b�t������� ��������(: L^p����� �� $6HZ �~������ �/ /G/D/V/h/z/ �/�/�/�/�/�/?
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8___�\_��VPRG_CoOUNT��@����RENBU��UM��S��__UPD �1�/�8  
 s_�oo*oSoNo`o ro�o�o�o�o�o�o�o +&8Jsn� �������� "�K�F�X�j������� ��ۏ֏���#��0� B�k�f�x��������� ҟ������C�>�P� b���������ӯί������UYSDE�BUG�P�P�)�d��YH�SP_PAS�S�UB?Z�LOoG ��U�S�)�#�0�  ���Q)�
MC:\x��6���_MPC����U���Qñ8� ��Q�SAV �b����ǲ&�η�SV;�TEM_T�IME 1��[k (m�4&�1:��}YT1SVGUNYS�P�U'�U����ASK_OPTICON�P�U�Q�Q���BCCFG Ì�[u� n�A�a�`a�gZo��߃ߕ� �߹�������:�%� ^�p�[������� �� �����6�!�Z�E��~�i���������&� ������&8��n Y�}�?��ԫ  ��(L:p ^������� / /6/$/F/l/Z/�/ ~/�/�/�/�/�/�/�/ 2?8 F?X?v?�?�? ?�?�?�?�?�?O*O <O
O`ONO�OrO�O�O �O�O�O_�O&__J_ 8_n_\_~_�_�_�_�_ �_�_o�_ o"o4ojo Xo�oD?�o�o�o�o�o xo.TBx� �j������ ��,�b�P���t��� ��Ώ��ޏ��(�� L�:�p�^�������ʟ ��o��6�H�Z� ؟~�l�������د� ��ʯ ��D�2�h�V� x�z���¿���Կ
� ��.��>�d�Rψ�v� �Ϛ��Ͼ�������*� �N��f�xߖߨߺ� 8���������8�J� \�*��n������ ������"��F�4�j� X���|����������� ��0@BT� x�d���� �>,Ntb�� ����/�(// 8/:/L/�/p/�/�/�/ �/�/�/�/$??H?6? l?Z?�?~?�?�?�?�? �?O�&O8OVOhOzO �?�O�O�O�O�O�O
_ _�O@_._d_R_�_v_ �_�_�_�_�_o�_*o oNo<o^o�oro�o�o �o�o�o�o J 8n$O����� X���4�"�X�B��v��$TBCSG_GRP 2�B���  ��v� 
 ?�  ������׏���� ���1��U�g�z����ƈ�d, ����?v�	 HC�=�d�>����e�?CL  B���П�ܘ�����\})��Y  A�ܟf$�B�g�B�Bl��i�X�ɼ���X��  D	J���r�����AC����үܬ���D�@v�=�W�j�}�H� Z���ſ���������v�	V3�.00��	m6;1c�	*X�PĘu�g�p�>���v�(�:�� ��p͟� ; O����p������z�JCFG -�B��� ����+������=��=�c�q�K�q� �߂߻ߦ�������� '��$�]�H��l�� �����������#�� G�2�k�V���z����� ���������p* <N���l��� ����#5GY }h����v� b��>�// /V/D/ z/h/�/�/�/�/�/�/ �/?
?@?.?d?R?t? v?�?�?�?�?�?O�? *OO:O`ONO�OrO�O �O��O�O�O_&__ J_8_n_\_�_�_�_�_ �_�_�_�_�_oFo4o jo|o�o�oZo�o�o�o �o�o�oB0fT �x������ �,��P�>�`�b�t� ����Ώ������� &�L��Od�v���2��� ��ȟʟܟ� �6�$� Z�l�~���N�����د Ư�� �2��B�h� V���z�����Կ¿� ���.��R�@�v�d� �ψϪ��Ͼ������ �<�*�L�N�`ߖ߄� �ߨ����ߚ����� ��\�J��n���� �������"���2�X� F�|�j����������� ����.TBx f������� >,bP�t �����/�(/ /8/:/L/�/�ߚ/�/ �/h/�/�/�/$??H? 6?l?Z?�?�?�?�?�? �?�?O�?ODOVOhO "O4O�O�O�O�O�O�O 
_�O_@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<oro`o�o�o �o�o�o�o�o&�/ >P�/���� �����4�F�X� �(���|�����֏� ���Ə0��@�B�T� ��x�����ҟ����� �,��P�>�t�b��� ������������ :�(�^�L�n������� 2d�����̿�$� Z�H�~�lϢϐ����� ���Ϻ� ��0�2�D� zߌߞ߰�j������� ���
�,�.�@�v�d� ������������ �<�*�`�N���r��� ����������& J\�t��B� �����F4 j|��^���8�/�  2 6#� 6&J/6"�$�TBJOP_GR�P 2����  ?��X,i#�p,� ��xJ� �6$�  �<� �� �6$� @2 �"	 ��C�� �&b  �Cق'�!�!>��1�
559>�0+1��33=�C�L� fff?+0?�ffB� J1�%Y?�d7�.��/>���2\)?0�5����;��hCY�� �  @� �!B�  A�P?�?�3~EC�  D�!8�,�0*BOߦ?�3�JB��
:���Bl�0��0�$�1�?�O6!Aə�A�̔C�1D�G6�=qq�E6O0�p��B��Q�;�A}�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH�1�ts�A@33@?1� C�� �@�_x�_&_8_>��D�U�V_0�LP�Q30<{�zR� @�0�V�P !o3o�_<oRifoPo^o �o�o�oRo�o�o�o�o M(�ol�p~(��p4�6&�q5	V3.00�#�m61c�$*�(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I�R�CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;S@;Q��|8�`rz@/&�8�6&<��1�w�^$�ESTPARS c *({ _#HR��ABLE 1�p+IZ�6#|�Q� � 1�|�|�|�5'=!*|�	|�
|�|�˕�6!|�|�|�N��RDI��z!ʟ@ܟ� ��$���O�������¯ԯ�����S��x# V���˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� U-����ĜP�9�K�]� o��-�?�Q�c�u���~6�NUM  ��z!� >  �Ȑ����_CFG ������!@b IMEBF_TT��p��x#��a�VER���b�w�a�R 1Ξp+
 (3�6"1 ��  6!������ ���� �9�$�:�H�Z� l�~����������������^$��_��@�x�
b MI_CH�ANm� x� kDOBGLV;0o�x��a!n ETHERA�D ?�� ��y�$"�\&n R�OUT��!p*!�*�SNMA�SK�x#�25�5.h�fx^$O�OLOFS_DI�[ՠ	ORQC?TRL �p+;/ ���/+/=/O/a/ s/�/�/�/�/�/��/��/�/!?��PE_D�ETAI��PON_SVOFF��33P_MON ��H�v�2-9STRTCHK ����42VTCOM�PATa8�24:0FPROG %��%MULTIROBOTTO!O06��PLAY��L:_�INST_MP 2GL7YDUS���?��2LCK�LPKQUICKMEt �O�2oSCRE�@�
tps��2�A�@�I��@_Y���9��	SR_GRP �1�� ���\�l_zZg_�_�_�_�_�_�^�^�oj �Q'ODo/ohoSe��o o�o�o�o�o�o�o !WE{i�������	1234567��!�ڎ�X�E1�V[
 ��}ipnl/�a�gen.htm�no��������ȏ~��Panel s/etup̌}�?�`�0�B�T�f� �� 񏞟��ԟ���o� ���@�R�d�v����� �#�Я�����*� ��ϯůr��������� ̿C��g��&�8�J� \�n�����϶����� ����uϣϙ�F�X�j� |ߎߠ����;��������0�B��*NUA�LRMb@G ?�� [������ ������ ��%�C�I��z�m�������v�SEoV  �����t�ECFG �Ё=]/BaA$  w B�/D
 �� /C�Wi{��� ���� PRց; �To\o�eI�6?K0(%�� ��0�����/ /;/&/L/q/\/�/�/�/l�D �Q�/�I_�@HIST �1ׁ9  (�  ��(/S�OFTPART/�GENLINK?�current=�menupage,153,1 E�c0p?�?�?�?/C��9 >?P=962n?�?�
OO.O�?�?�136 c?|O�O�O�OAOSO�? �O__0_�O�O_Lu_ �_�_�_:_�/�_�_o o)o;o�__oqo�o�o �o�oHo�o�o%7I~��a81�ou� �����o��� )�;�M��q������� ��ˏZ�l���%�7� I�[���������ǟ ٟh����!�3�E�W� ���������ïկ� v���/�A�S�e�P b������ѿ����� �+�=�O�a�s�ϗ� �ϻ�������ߒ�'� 9�K�]�o߁�ߥ߷� �������ߎ�#�5�G� Y�k�}�������� �������1�C�U�g� y���v����������� 	�?Qcu� �(���� )�M_q��� 6���//%/� I/[/m//�/�/�/D/ �/�/�/?!?3?�/W? i?{?�?�?�?�����? �?OO/OAOD?eOwO �O�O�O�ONO`O�O_ _+_=_O_�Os_�_�_ �_�_�_\_�_oo'o 9oKo�_�_�o�o�o�o �o�ojo�o#5G Y�o}�������?��$UI_P�ANEDATA �1������  	�}�0�B�T�f�x��� )����mt�ۏ� ���#�5���Y�@�}� ��v�����ן����� ��1��U�g�N������ �1��Ïȯ گ����"�u�F��� X�|�������Ŀֿ=� �����0�T�;�x� _ϜϮϕ��Ϲ������,ߟ�M��j�o� �ߓߥ߷������`� �#�5�G�Y�k��ߏ� ������������� �C�*�g�y�`����� ����F�X�	-? Qc����߫�� ��~;"_ F��|���� �/�7/I/0/m/�� ���/�/�/�/�/�/P/ !?3?�W?i?{?�?�? �??�?�?�?O�?/O OSOeOLO�OpO�O�O �O�O�O_z/�/J?O_ a_s_�_�_�_�O�_@? �_oo'o9oKo�_oo �oho�o�o�o�o�o�o �o#
GY@}d ��&_8_���� 1�C��g��_������ ��ӏ���^���?� &�c�u�\�������ϟ ���ڟ�)��M�� ���������˯ݯ0� ����7�I�[�m�� ��������ٿ�ҿ� ��3�E�,�i�Pύϟ�����Ϫ���Z�l�}����1�C�U�g�yߋ�) ߰�#������� �� $�6��Z�A�~�e�w� �����������2� �V�h�O�����v�p���$UI_PAN�ELINK 1��v�  ��  ��}�1234567890����	-? G ���o���� �a��#5GD�	����p&���  R����� Z��$/6/H/Z/l/ ~//�/�/�/�/�/�/ �/
?2?D?V?h?z?? $?�?�?�?�?�?
O�? .O@OROdOvO�O O�O �O�O�O�O_�O�O<_�N_`_r_�_�_�0, ���_�X�_�_�_ o2o oVohoKo�ooo�o�o �o�o�o�o��, >r}������� �����/�A�S� e�w��������я� ��tv�z����=� O�a�s�������0S�� ӟ���	��-���Q� c�u�������:�ϯ� ���)���M�_�q� ��������H�ݿ�� �%�7�ƿ[�m�ϑ� �ϵ�D��������!� 3�Eߴ_i�{�
�߂� ���߸������/�� S�e�H���~��R~ '�'�a��:�L�^� p���������������  ��6HZl~ ���#�5���  2D��hz�� ���c�
//./ @/R/�v/�/�/�/�/ �/_/�/??*?<?N? `?�/�?�?�?�?�?�? m?OO&O8OJO\O�? �O�O�O�O�O�O�O[� _��4_F_)_j_|___ �_�_�_�_�_�_o�_ 0ooTofo��o��o ��o�o�o,> 1bt����K ����(�:��� �{O������ʏ܏� uO�$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v�������� п���ϕ�*�<�N� `�rτ��O�Ϻ�Io�� �������8�J�-�n� ��cߤ߇����߽��� �o1�oX��o|�� ������������ 0�B�T�f�������� ������S�e�w�,> Pbt��'�� ���:L^ p��#����  //$/�H/Z/l/~/ �/�/1/�/�/�/�/?  ?�/D?V?h?z?�?�? �???�?�?�?
OO.O ��ROdO�߈OkO�O�O �O�O�O�O_�O<_N_ 1_r_�_g_�_7O�M�m�$UI_Q�UICKMEN � ���_AobRESTO�RE 1��  � |��Rto�o�im�o�o �o�o�o:L^ p�%����� �o����Z�l�~� ����E�Ə؏����  �ÏD�V�h�z���7� ������/���
��.� @��d�v�������O� Я�����ßͯ7� I���m�������̿޿ ����&�8�J��n� �ϒϤ϶�a������� Y�"�4�F�X�j�ߎ� �߲������ߋ����0�B�T�gSCRE�`?#muw1sco`u2��U3��4��5��6���7��8��bUSE�Rq�v��Tp���k�s����4��5��6���7��8��`ND�O_CFG ܶ#k  n` `P�DATE ���Noneb�SEUFRAME�  �TA�n�R�TOL_ABRT8y�l��ENB����?GRP 1�ci/aCz  A��� ��Q�� $6H!Rd��`U����~��MSK  ��4���Nv�%�U��%���bVISCAND_MAX��I��FAI�L_IMG� �P��P#��IMRE/GNUM�
,[gSIZ�n`�A��,VONTMOiU��@����2��a��a�����FR:�\ � �MC:\�\LO�G�B@F� !��'/!+/O/�Uz? MCV�8#oUD1r&EX{+�S�PPO64�_��0'fn66PO��LIb�*��#V���,f@��'�/� =	�(S�ZV�.����'W�AI�/STAT' ����P@/�?��?�:$�?�?��2�DWP  ���P G@+b=���� H�O_JMPERR 1�#k�
  �2345?678901dF�� �O{O�O�O�O�O�O_ �O*__N_A_S_�_
� MLOWc>
 ��_TI�=�'�MPHASE � ��F��PSoHIFT�1 9�]@<�\�Do�U #oIo�oYoko�o�o�o �o�o�o�o6l CU�y���� � ��	�V�-�e2�����	VSFT]1�2	VM��� �5�1G� ���~%A�  B8̀̀�@ pكӁ˂1�у��z�ME@��?�{��!c>&%�JaM1��k�0�{ ��$`0TDINE#ND��\�O� �z����S��w��P����ϜRELE��Q��Y���\�_ACTIV��:�R�A ��e���e��:�RD� ���YBOX �9�د�6���02���190.0.��83��25�4��QF�	 ��X�j��1��robot��� ?  p�૿�5pc��̿������7�����-�f�ZWABC�����,]@ U��2ʿ�eϢωϛ� �Ͽ����� ���V�@=�z�a�s߰�E�Z��1�Ѧ