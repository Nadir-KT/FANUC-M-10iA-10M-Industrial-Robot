��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1��GPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|�(�ARG_S�TR1 � �$TITP$I��1�{������5�6�7*�8�9�0��@z�����1�U1�1 '1
'2"�GSBN_CFG�1  8 $�CNV_JNT_�* |$DATA�_CMNT�!$�FLAGS�*C�HECK�!�AT�_CELLSET�UP  P �$HOME_I�O,G�%�#MA�CRO�"REPR��(-DRUN� D�|3SM5H UTOBACKU0� � $EN�AB��!EVICv�TI � mD� DX!2ST� �?0B�#$INTE�RVAL!2DIS?P_UNIT!20w_DOn6ERR�9�FR_F!2IN^,GRES�!0�Q_;3!4C_WA��471�8���AW�+0�$Y $DB\� 6COMW!2�MO� 21H A.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3��B�2���AXD��#
 d $�CARD_EXI�ST4$FSS�B_TYP!AH�KBD_SNB�1A�GN Gn $�SLOT_NUM��APREV4D�EBU� g1G ;1_�EDIT1 �� 1G=� S<�0%$EP�O$OP�U0LETE_OK�B{US�P_CR�A�$;4AV� 0LACIw1�R�@k ܢ1$@MEN�@$D�V�Q`PvVA�{QL� OU&R� ,A�0�!� B�� LM_O�
eR��"CAM_;1� xr$AT�TR4�@� ANN�N@5IMG_HE�IGH�AXcWID�TH4VT� �U�U0F_ASPEC��A$M�0EXP��.@AX�f�CF��D X $GIR� � S�!.@B�P�NFLI�`�d� U�IRE 3T!GITSCH+C�`N� S�d�_LZ`AC�"�`E�Dp�dL� J�4S��0� <za�!p;G�0 � 
$WARNM�0f�!�@�� -s�pNST� C�ORN�"a1FLT�R{uTRAT� T�}p  $AC�Ca1�p��|{�rOcRI�P�C�kRT0�_S~B\qHG,I.1 [ T�`�"3I�pTY4D�@*
2 3`#@� �!�B*HDDcJ* Cd�U2_�3_�4_�5_�U6_�7_�8_�94v�ACO�$ <� ��o�o�hK3 1#`O_�Mc@AC t 2� E#6NGPvABA� �c1�Q8��`,��@nr1�� d�aP�0e���axnpUP&Pb26���p�"MJ�p_R�rPBC��1J�rĘߜJV�@U�� B��s}�g1�"YtP�_*0OFS&R @� RO_K8T��a�IT�3T�NOM_�0�1p�34 >��D� �� Ќ@��hPV��mEX�p� �0g0�ۤ�p�r
$TF��2C$MD3i�T�O�3�0U� F� K��Hw2tC1(�	Ez�g0#E{"F�"F�40CP@�a2 m�@$�PPU�3N)ύRև�AX�!DU��AI�3BUF�F=�@�1 |pp���pP�IT� PP�M��M�y��F�SIMQSI�"ܢVA�ڤT�Q=�w T��`(zM��P�B�qF�ACTb�@EW��P1�BTu$?�M]C� �$*1�JB`p�*1DEC���F��ŏ�� ��H0CHNS_E;MP1�$G��8�B�@_4�3�p|@P��3�TCc�(r/�0-s x��ܐ� MBi��!����JR� i�SEGKFR��Iv �aR��TpN�C��PVF�4S?�bx &��f{uJc!�Ja���� !28�ץ�AJ���SCIZ�3S�c�B�TM����g��JaRSINFȑb���q�۽�������L�3�B���gCRC�e�3CCp ����c��mcҞb�1@J�cѿ�.����D$ICb�Cq�5r�ե��@�v�'���EV���zF*��_��F,pN��ܫ��?�4�0A�! �r���h�Ϩ�� p�2�͕a�� �د�p�R�Dx @Ϗ��o"27�!ARV�:O`C�$LG�pV��B�1�P��@�t�aA�0'�|�+0Ro�� �MEp`"1 CRA 3 AZV�g6p�O �FCCb�`�`�F�`K������ADI��a�A�bA'�@.p��p�`�c�`S4P�Ƒ�a�AMP��-`Y$�3P�M�]pUR��Q�UA1  $@TITO1/S@S�!�����"0�DBPXWO���B0!5�$SK4���28@DBq�!�"�"�PR�� �
� =����!# lS q1$2�$z�/ �L�)$�/PA���� %�/�#P�C�!&?4ENE��q.'*?�#� R�E�p2(H z��O�0#$L|3$$�#�B[�;���F�O_D��RO�Sr�#������3R�IGGER�6PA�pS����ETURN��2�cMR_8�TUrw��0EWM�ҍM�GN�P���BL�AH�<E���P��'&$P� �'P@�Q"3�CkD{��DQ���4�11��FGO_A7WAY�BMO�ѱQ�#!�DCS_޾)  �PIS � I gb {s�C��A��[ �B$�S��A�bP�@�EW-�TNT	Vճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_�SV�bEXCLUt��nONL2�b�SY�*a&�OT�a'�HI_V�4��B<���_ *P0� �9�_z��p v�TSG�� +nr r�@6Acc*b��G�#@�E�V.iHb?fANNcUN$0.$fdID�	U�2�SC@�`�i�a@��j�f�z��@I$2,O�$FibW$}��OT9@�1 $DUMMYk��da���dn�� � �E- 7` ͑HE4(s�g�*b�SAB��SUF�FIW��@CA*=�c5�g6�a��DMSW�E. 8�̀KEYI5���T�M�10s�qA�vIN���#�b��/ Dބ�HOST_P! �rk��ta��tn��tsp��pEMӰV��C�ڪpLc ULI�0 � 8	=ȳ����DTk0�!1 � �$S��ESAMPL��j�۰f璱f����I�0��[ $SUB�k�#0�C��T�r#a�SAVʅ��c��`�C��P�fP$n0yE�w YN_B#72 0�`DI{dlp�O(��9#$�R�_I�� �EN�C2_S� 3 ! 5�C߰�f�-  �SpU����!4�"g��޲�1T���5@X�j`ȷg��0�0K�4x�AaŔAVER�q8ĕ9g�DSP�v��PC��r"��(����ƓVALUߗHE4�ԕM+�IPճ���OPP ��TH��֤��P�S� �۰	F��df�J� �q�#(T�ET+�6 H�bLL_DUs�~a3@{��3:���OTX"���so�~�0NOAUTO�!7�p$)�$�*��c�4�(�C�8�C�, �"�q&�L�� �8H *8�L H <6����c"�`,  `Ĭ�kª�q��q��Psq��~q��7��8���9��0����1��1�̺1ٺ1�1�1� �1�1�2(�2T����2̺2ٺ2�U2�2 �2�2ʕ3(�3��3��̺3�ٺ3�3�3 �3
�3�4(�ɢT�?��!9 <�9�&�z���I��1���M��QFqE@'@� : ,6���Q? �@P?Q9��5�9�E�@�A��q�A� ;p�$TP�$VA�RI:�Z���UP2f�P< ���TDe�@��K`Q�����wBAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�H  ��P�!�F@`�!>t ;E��sC�ST�D�  D���c�<� 	C�� {��_���l���R  ����FORCEUyP?b��FLUS�`�H�N>�F ���RD_CM�@E������� ��@vMP��REMr F�Q��1������7Q
K4	NJ�5EcFFۓ:�@IN2Q��OVO�OVA��	TROV���DyTՀ�DTMX�  ��@�
ے_PHX"p��CL��_Tp�E�@�pK	_(�Y_QT��v(��@A;Q	D� ������!0�tܑ0RQ���_��a����M�7�CL�dρRIV'�{���EARۑIOHP�C�@����B�B��C�M9@���R �GgCLF�e!DYk(�M�ap#5TuDGЫ�� �%!ʠFS9SD �s? P�a�!�1���P_�!�(�!�1��E�3�!3�+5��&�GRA��7�@ҕ�;�PW��ON<n��EBUG_SD2�H �{�_E� A �p�R _�TERM`5Bi5N��ORI#:e0C�9SM_�P��Ze0D�9TA�9E�9�UP\�F� -��A{�AdPw3S@B�$SEG�:� EL�{UUSE�@NFIJ�B$�;1젎4�4�C$UFlP=�!$,�|QR@��_G�90Tk�D�~SNST��PAT����AP'THJ3Q�E�p% B`�'EC���A�R$P�I�aSHFT�y�A�A�H_SHOQRР꣦6 �0$�7rPE��E�OVR=���aPI�@�U�b �QAYLOW����IE"��A��?���ERV��XQ�Y��mG�>@�BN��U���Rz2!P.uASYMH��.uAWJ0G�ѡE q�A�Y�R�Ud>@ ��EC���EP;�uP�;�6WOR>@M`�]0SMT6�G3�cGR��13�aPAL@��P��q�uH � u���TOCA��`P	P�`$OP@����p�ѡ�`0YO��RE�`R4Cb�AO�p낎Be�`�R�Eu�h�A��e$7PWR�IMu�R�R_�cN��q=B �I&2H���p_AD�DR��H_LENAG�B�q�q�q$�R��S�JڢSS��SKN��u���u̳�uٳ�SE�A�ʠHS���MN�!K��`���b����OLX���p����`ACRO3pJ�@��X�+��Q8��6�OUP3�bE_�IX��a�a1�� }򚃳���(��H���D��ٰ��氋�IO2S�D�����x�`�7�L $d�<�`Y!_OFFr���PRM_��x�H�TTP_+�H:�M; (|pOBJ]"�p���$��LE~C|d���N � ��.֑AB_�Tqᶔ�S�`H�LVh�K�R"uHITCOmU��BG�LO�q���h�����`���`SS� ���HW��#A:�Oڠ<`I�NCPU2VISIOW�͑��n��to���to�ٲ �IOL]N��P 8��R��^r�$SLob oPUT_n�$p¾�P& ¢��Y F_�AS�"Q��$L ������Q  U�0	P�4A��^���ZPHY���-��Ky��UOI �#R `�K���@�$�u�"pP�pk���$�����Y�UeJ5�S-���NE6W�JOGKG̲DISĖ��Kp���#T �(�uAVF�+`�CTyR�C
�FLAG2v�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w� m� _�{0a�^��cg���4� ����Ǝ���{0��� �SCH_���a�SLN�d�VW���AE�"����4��UM��Aљ`LJ�@�DAUf�EAU�p��d|�r��GH�bD���BOO>��WL ?�6 �IT��y0�REC��SCR ܓ��D
�\���MARG m�!��զ ��d%�����S����W���U�� �JGM[�MNC�HJ���FNKEY�\�K��PRG��UqF��7P��FWD��HL��STP��V`��=@��А�RS��HO`����C9T��b ��7�[�UL���6� (RD� ����Gt��@CPO��������MD��FOCU��RGE]X��TUI��I��4�@�L��� ��P����`��P��9NE��CANA��B�j�VAILI�CL� !�UDCS_HII4��s�O�(!��S���S���� ��BUFF�!Xj�?PTH$m�@��v`��a���AtrY�?P��j�3��`WOS1Z2Z3Z�q1�� � Z � ���[aEȤ��ȤIKDX�dPSRrO�X��zA�STL�R}��Y&�� Y$E�C���K�&&8y�� [ LQ�� +00�	P���`#qdt
��U�dw<���_ \ ?�4Г�\��Ѩ#� �MC4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#b�D���'B�LD�%�$�%ORGڰ5�2 �PVŇVY8�s�T�r�$}d^ ���$6��$
�%S�`T� �B0�4}�6RCLMC�4`]?o?�9세�MI�p�}d_ d=њRQz��DSTB�pƽ ;F�HHAX��R JHdLEXC#ESr1!BM!p�a%`ip/B�TE�j�`a�p=F_A7J�i��KbOtH� K�db� \Q���v$MB�C�LI|�)SREQUIR�R�a.\o�AXODEBUZ�ALt M��c�b�{P����2ANDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��XB� N&��aZ���UwPST� ezr7LOC�RIrp�EX<fA�p�9AA�ODAQ��f XfY�OND��"MF,� �Łf�s"��}%�e/�� ��AFX3@IGG>�� g ��t"���ܓs#N�s$R�a%��iL��hL�v�@��DATA#?pE��%�tR��Y�Nh t $MD`qI}�)nv� ytq�yt�HP`�Pxu��(�zsANSW)�yt@��yu�D+�)\b���0o�i[ �@CUw�V�p� 0XeRR2��j �Du�{Q��7Bd$C'ALIA@��G���2��RIN��"�<OS�INTE��Ck�r^�آXb]���_N�qlk���9�Dt���Bm��DIVF�DH�@���qnIc$V,��S�$��$Z�X�o�*�����oH ��$BELT�u!A/CCEL�.�~�=�IRC�� ���D�yT�8�$PS�@
�"L�@�r��#^��S�Eы T�PATH3���I���3x�p�A�_W��ڐ���2nC܍�4�_MG�$�DD��T���$FW�Rp9��I�4���DE7�PPABN���ROTSPEE�[g�� J��[��C@4��@$USE�_+�VPi��SYhY���1 �aYN!@9A�ǦOFF�qǡ7MOU��NG���sOL����INC�t�Ma6��HB��0HBENCS+�8q9Bp�4�,FDm�IN�Ix�]��B��VE��#�y��23_UP񕋳LOWL���p� B���Du�9B#P`�x 䳵�BCv�r�MOSI��BMOU��@�7PERCH  ȳOV��â
ǝ�� ��D�ScF�@MP������ Vݡ�@y�j�L`Uk��Gj�p�UP=�8����ĶTRK��AYLOA�Qe��A���x�����N`�F�RcTI�A$��MOU� ��HB�BS0�p7D5����ë�Z�DUM�2ԓS_BCKLSH_Cx�k��� �ϣ���=���ޡ �	ACLAL"q��18м@��CHK� �S�RTY��^��%E1Qq_�޴_U�M�@�C#��SC�L0�r�LMT_J'1_L��9@H�qU�EO�p�b�_�e�k�e�SPC��u���&N�PC�N�Hz \Pd��C�0~"XT�.�CN_:�N9��&I�SF!�?�V���@U�/���x�T���CB!�SH�:��E�E1 T�T����y���T��3PA ��_P��_� =������!�����J6 L�@��O�G�G�TORQU��ONֹ��E�R���H�E�g_W2���_@郅���I��I�I��Ff`xJ��1�~1�VC3�0BD�B�1�@SBJRKF9�0?DBL_SM��2�M�P_DL2GRV����f�H_��d���CO1S���LNH� �������!*�,�aZ���fM1Y�_(�TH��)�THET0��NK�23���"��CB�&CB�CAA�B�"`��!��!�&SB 2�%GTS�Ar�C IMa�����,4#97#$DU���H\1@� ��Bk62��AQ(rNSf$NE�D�`I���B+5��$̀�!A��%�5�7���LP!H�E�2���2SC %C%�2-&FC0JM&�̀V�8V�8߀LV�JV!KV/KV=KV*KKVYKVgIH�8F�RM��#X!KH/KH�=KHKKHYKHgIOJ�<O�8O�YNOJUO!KO/KO=KOKKOYKOM&F�2�!+i�%0d�7SPBAL�ANCE_o![cLmE0H_�%SPc�� &�b&�b&PFULC�h�b�g�b%p�{1k%�UTO_�ОT1T2�i/�2N��"�{�t#�Ѱ`P�0�*�.�T��OÀ|<�v INSEG"��ͱREV4vͰl�D3IF�ŕ�1lzw��1m�0OBpq�я�?�MI{���nLC�HWARY���AB���!�$MECH`�!o ��q�AX���P����7Ђ�`n �
�d(�U�ROB���CRr�H���(?�MSK_f`�_p P �`_��AR/�k�z�����1S�~�|�z�{���z��qI�NUq�MTCO�M_C� �q � ���pO�$N'OREn����pЂor 8p GRe��uSD�0AB�$XYZ_DA�1<a���DEBUUq�������s z`$��C;OD�� L����p�$BUF�INDX|�  �<�MORm�t $فUA��֐���Д�r�<��rG��u �� $SIMU�L  S�*�Y�̑a�O�BJE�`̖ADJ�US�ݐAY_I�S�D�3����_[FI�=��Tu  7�~�6�'��p} =�C��}p�@b�D��FRI4r��T��RO@ \��E}��y�OPW�OYq�v0Y�S�YSBU/@v�$SCOPġd���ϪUΫ�}pPRUN����P�A��D���rɡL�_�OUo顢q��$)�IMAG��4w��0P_qIM��L��INv�K�RGO�VRDt��X�(�P0*�J�|��0L_�`]񘘵�0�RB1�02��M��ED}��p� ��N�PMֲ��̮�x�SL�`q�w �x $OVSL�4vSDI��DEX�����#���-�V} *�N4�\#�B�2èG�B�_�M�r���q�E� x Hxw��p��ATUSWЅ��C�0o�s���BSTM�ǌ�I�k��4��x�԰q�y DBw�E&���@E�r���7��жЗ�EXE ��ἱ�����f q�gz @w���UP'�f�$�pQ�XN����������� �P�G΅{ h $GSUB����0_��|�!�MPWAIv�P7ã�LOR�٠F�\p˕$RCVF�AIL_C��٠B�WD΁�v�DEF�SP!p | L�w���Я�\���UCNI+�����H�R�,p}_L\pP��x�t���p�}H�> �*��j�(�s`~�N�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��Gc�PLI��p��  $ˀP_�SWI�p��y�J_�PL��AL_ )�����A��B��� uC��D�$E�[�.�C_�U�� � � ����*�J3K0����TWIA4��5��6��MOM�������4��ˀB��AD����؟�����PU� NR ��������m���� A$PI �6q��	����� K4�)6�U��w`��_SPEEDgPG� �������Ի�4T��� � @��SAMr`��\�]��MOV_�_$�npt5���5���1���2���������'�S�Hp�IN�'�@� +����4($4+T+�GAMMWf�1'��$GET`�p���D�a���

pLIBRt>�II2�$HI=�!_g�t��2�&E;��(1A�.� �&LW�-6 <�)56�&]��v�p���V��$PD#CK���q��_?�����q�&���7����4���9+� ��$IM_SR�pD`�s�rF��r�rLE��¹Om0H]��0��-�pq��PJqUR_SCRN�FA����S_SAVE_�D��dE@�NOa�C AA�b�d@�$q�Z�I ǡs	�I� �J�K� �� ��H�L��>�"hq ������ɢ��  bW^US�A�   �M4���a��)q`� �3�WW�I@v�_�q�.�MUAo�� � �$PY+�$W�P�vNG�{��P:���RA��RH��RO�PL������q� ��s'�X;�OI�&�Zxe ����m�� p��ˀ�3 s�O�O�O�O�O�aa�_т� |��q�d@ ��.v��.v��d@��[wdFv��E���% ���u;B�w�|�tPn���PMA�QUa ��Q8��1٠wQTH�HOLW�oQHYS��ES�F�qUE�pZB��Oτ�  ـPܐ(�AP����v�!�t�O`�q��u�"���FA��IGROG�����Q2����o�"��p��INFOҁ�׃V����R��H�OI��� (�0SLEQ����@��Y�3����Á��P�0Ow0���!E�0NU��AUT<�A�COPY�=�(/�'��@Mg�N��=��}1������ ��RG4��Á���X_�P�C$;ख�`��W���P��@�������E�XT_CYC b�HᝡRpÁ�r��_NAe!А����ROv`	�� �s ���POR_�1�E2�SRV �)l_�I�DI��T_� k�}�'���dЇ�����U5��6��7��8i��H�SdB���2�$R��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,�0FL`�o@SYN��K�M��Ck��PWR+�9ᘐ���DELA}�dY��pAD�a�'��QSKIP4�� �A�$�OB`NT2����P_$�M� ƷF@\bIpݷ�ݷ� ݷd����빸��Š��Ҡ�ߠ�9���J2R� ��� 46V�EX� TQQ�� ��TQ������ ��`��#�RDC�V� �`��X)�R�p������r��m$RGEA�R_� IOBT�2FcLG��fipER��DTC���Ԍ���2T�H2NS}� 1����G T\0 ����u�M\Ѫ`I��dG�REF�1�Á� l�h��ENsAB��cTPE�0 4�]����Y�]��ъQ n#��*��"�������2�Қ�߼���������3�қ'�9�K�P]�o���4�Ҝ��@�����������5���!�3�E�W�i�{��6�Ҟ�������������7�ҟ-?PQcu�8�Ҡ������ ^��SMSKÁ�l�i�a��EkA��oMOTE6������@�݂TQ�IO�}5�ISTP?��PsOW@��� �pJ���n �������E�"$DSB_SIGN�1UQ�x��C\�TP��S232���R�iDEVI�CEUS�XRSRP�ARIT��4!OP�BIT�QI�OWCONTR+�TQ���?SRCU� MpSU_XTASK�3N�p��0p$TATU�P�E#�0�����p_�XPC)�$FRE?EFROMS	pna��GET�0��UPeD�A�2�SP� �:��� !$USAN�na&�����ERI�0_�RpRIYq5*"_j@_�Pm1��!�6WRK9KD����6��QFRIE3ND�Q�RUFg�҃��0TOOL�6MY��t$LENGT�H_VT\�FIR��pC�@ˀE> +IU�FIN-RM��R�GI�1ÐAITI��$GXñ3IvFG2v7G1���p3�B�GcPR�p�1F�O_n 0��!RE��p�53҅U�TC��3A�A�FG�G(��":���e1n!��J�8�%���%]�U�%�� 74��X O0�L
��T�3H&��8���%�b453GE�W�0�WsR�TD����T��M�����Q�T]�$V �2����1�а91T�8�02�;2k3�;3�:ifa�9-i�aQ0��NS��ZR$V��2B%VwEV�2A Q�B
;�����&�S�`���F�"�k�@�2a�PS�E��$r1C���_$Aܠ6wPR��7vMU�cS�t '�/89�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx_�����BSOC����N��DUMMY�14�p@SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU""ƐS�P �M�)0NS��cM�"r�$HW_C��U��S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}��#!�_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�S�A�pC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EG� �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G��+ AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC  o�ER|f�5� � $�@�_ A��!�PO���à�0#�V�_�MRAt�� d �� T��ٔERR�����;TY&���I��V�0�cz�TOQ�d�PL[ �d�"�� �?�w�! � p�p`T)0���_V1�Vr�aӔ����2ٛ2�E����@�H�E���G$W�����V!��$�P��o�c�I��aΣ	 HEL�L_CFG!�� 5��B_BA�Sq�SR3���� a#Sb���1��%��2��3��4���5��6��7��8���RO����I0�03NL�\CAB+�����ACK4�����,���2@�&�?�_PUf�CO. U�OUG�P~ ����m�������{TPհ_KAR�Ll�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h�8�]�l0SEM�4Ĳ(�M4�6�TYN�SO���DIZ�~�AӸ����m_TM�MOANRQ��k0E�����$KEYSWITCH���m���{HE��BEAT��E- LE~����ȅU��F!Ĳ���B�O�_HOM=OGREFUPPR&��y!�� [�C��O��-E�COC��Ԯ0_IO�CMWD
�a��'qk��� � Dh1$���UX���M�β<gPgCFORC���� ��m�OM.  �� @�5(�U��#P, 1��, 3���45��NPX_�ASt�� 0��A�DD���$SI}Z��$VAR��.�TIP/�.��A�ҹM�ǐ��/�1�$+ U"S�U!Cz���OFRIF��J�S���5Ԓ�NF�Ѝ�n � xp`SI���TE�C���CSGL��TQ2�@&����<� ��STMT��,�P �&BWuP��S�HOW4���SV|�$�� �Q�A00�@Ma}����@������&���5��U6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G��0 G���0G���@G���PG��1	1	1�	1+	18	1E	2���2��2��2��2���2��2��2��2���2��2	2	2�	2+	28	2E	3���3��3��3��3���3��3��3��3���3��3	3	3�	3+	38	3E	4��4��4��4��4���4��4��4��4���4��4	4	4�	4+	48	4E	5��5��5��5��5���5��5��5��5���5��5	5	5�	5+	58	5E	6��6��6��6��6���6��6��6��6���6��6	6	6�	6+	68	6E	7��7��7��7��7���7��7��7��7���7��7	7	7�	7+	78	7E*v	�VP��UPDs��  �`NЦ��
A�SYSLO>t�� � L��0d���A�aTA�0d��|�ALU:ed�~��CUѰjgF!aID�_L�ÑeHI�jI~��$FILE_����d��$2�
�cS�A>�� hO��`E_BLCK��b$�>�hD_CPUyM� yA��c�o�d�b�����R �Đ
PWl��!� oqLA���S=�ts�q~tRUN �qst�q~t���q�st�q~t�T��A�CCs��X ;-$�qLEN;��t�H��ph�_�I��ǀL�OW_AXI�F)1�q�d2*�MZ���ă��W�Im�ւ�aR�GTOR��pg�D�<Y���LACEk�ւp�pV�ւ~�_MA2�pv�������TCV��؁��T��ي����� t�V����V�Jj�R��MA�i�J��m�u�b����q2j�#�U��{�t�K�JK��VK�;���H���3��J0l����JJ��JJ��AAL��ڐ��ڐԖe4Օ5���N1��P�ʋƀW�LP�_(��g�!���pr�� =`�`GROUw`����B��NFLIC���f�REQUIRE3�EBU��qB���w�2����p���q�5�p�� \��A�PPR��C}�Y�
vްEN٨CLO7��S_M��H���u�y
�qu�� ����MC�����9�_M	G��C�Co��`M��ܲ�N�BRKL�NO�L|�N�[�R��_L!INђ�|�=�J����Pܔ������������������6ɵ�̲8�k�D����� ��
��q)��7�PATH3�L�B�L���H�wࡠ�J�CN��CA�Ғ�ڢB�I�N�rUCV�4a��C!�UM��Y,�����aE�p����ʴ���PAYLOA��J{2L`R_AN�q�Lpp���$�M��R_F2LSHR��N�LOԡ�Rׯ�|`ׯ�ACRL_G� �ŒЛ� ��Hj`߂�$HM���FLE�XܣE�J�u� :��������������1�F1 �V�j�@�R�d�v�������E����ȏڏ� ���"�4�q���6�M� ��~��U�g�y�ယ	T��o�X��H����� �藕?�����ǟِ ݕ�ԕ����%�7���JJ�� � `V�h�z���`AT��l��@�EL�� Sj��J|�Ŝ�JEy�gCTR��~�TN���FQ��HAND_�VB-���v`�� $��F2M�����ebSW�q�'��?� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)F�QAW�Z`i�Aw�A��PX X�'pi�Dw�D��ePf�G�p�)STk�h�!x��!N��DY�p נM�9$`%Ц�H�� H�c�׎���0� ��Pѵڵ�������8����� ����1��R�6��QASYIMvř���v��J�8��cі�_SH>��� �Ĥ�ED����������J�İ%��C�ID�.��_VI�!X�>2PV_UNIX�FThP�J��_R�5_Rc� cTz�pT�V��@���İ�߷��U �����2��Hqpˢ��a3EN��`DI����O4d�'�p`J�S� x g"IJAAȱ z�aabp�coc�`aE��dq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a�i�T�@<� $D�UMMY9Q�$�PS_��RFC� 9 S�v E����Pa� XƠ����STE���SBR�Y�M21_VF�8�$SV_ERF�O���LsdsCLRJtA���Odb`O�p �� D $GgLOBj�_LO����u�q�cAp�r�@aS;YS�qADR``�`TCH  �� ,��ɩb�W_N�A���7��S�R���l  ���
*?�&Q�0"?� ;'?�I)?�Y)��X��� h���x������)��Ռ �Ӷ�;��Ív�?��O�O�O�DFaXSCR�E栘p����ST��s}y`���_   �/_H�A�q� TơgpTYP�b���G�a�G���Od0ISb_䓀e�UEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI� m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� d�� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1 �ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���}� VSHIF��Nc�P�`ג�E��ȐR����OSURz��Wk`RADIL����_�a��:�9a���`a�r��LULQ$�OUTPUT_BM����IM�AB ��@�rTILSCO��C7��� ����&��3�� A���q���m�I�A2G�pq�y@Md�}���yDJU��N�/WAIT֖�}���{�%! NE�u�Y�BO�� ��� $`�t�SB�@TPE��NEC�p�J^FY�nB_T��R�І�a$�[$YĭcB��dM����F� �p�$�pb�O�P?�MAS�_DUO�!QT�pD���ˑ#%��p!"DELcAY�:`7"JOY� @(�nCE$��3@ 0�xm��d�pY_[�!"��`�"��[���P?� �F`ZABC~%��  $�"�R��
p�$$C�LAS����i��!pp � �VIRT]��/ 0A�BS����1 5�� < �!F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ8i{0-�AXL�p2���!�63  �{tIqN��qztPRE�����v�p�uLAR�MRECOV �9�rwtNG�� �.;	 A  � �.�0PPLIMC��?5�p��HandlingToolϐ�o� 
V7.5�0P/23-�  o�Pz��
��w_SWt� UP�!7� x�F0��t��QzA� v�� 864�� ��it�y�2���" 7DA�5�� �� d�@��o�None�isͅ˰ ���T���!�AyWx>�_l�V�utT��s9�UTO�"�Њt�y��HGAPCON
0g�1��Uh�oD 1581����̟ޟry����/Q 1���p �,�蘦���;�@���q_��"�" g�c�.�H����D�HTTHKYX��"�-�?�Q��� ɯۯ5����#�A�G� Y�k�}�������ſ׿ 1�����=�C�U�g� yϋϝϯ�����-��� 	��9�?�Q�c�u߇� �߽߫���)����� 5�;�M�_�q���� ����%�����1�7� I�[�m���������� !����-3EW i{����� �)/ASew ����/��/ %/+/=/O/a/s/�/�/ �/�/?�/�/?!?'? 9?K?]?o?�?�?�?�? O�?�?�?O#O]����TO�E�W�DO_CLEAN�����C�NM  � �__/_A_S_�DSPDRYR�O&��HIc��M@�O�_ �_�_�_oo+o=oOo aoso�o�o���pB��v# �u���aX�t�������9�PLUGGp���G��U�PRCvPB�@��_�or�Or_��SEGF}�K[mwxq�O�O������?rqLAP�_�~q�[�m���� ����Ǐُ����!�|3�x�TOTAL�f| yx�USENU�p��� �H���B��R�G_STRING� 1u�
�kMn�S5�
ȑ�_ITEM1Җ  n5�� ��$�6� H�Z�l�~�������Ư�د���� �2�D��I/O SIG�NAL̕Tr�yout Mod�eӕInp��S�imulated�בOut���OVERR�P =� 100֒In� cycl��ב�Prog Abo�r��ב��Sta�tusՓ	Hea�rtbeatїMH Faul��Aler'�W�E� W�i�{ύϟϱ������� �CΛ�A�� ��8�J�\�n߀ߒߤ� �����������"�4��F�X�j�|���WOR {pΛ��(ߎ����� � �$�6�H�Z�l�~��� ������������ 2PƠ�X �� A{������ �/ASew������SDEV[�o�#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g?>y?PALTݠ1 ��z?�?�?�?�?O"O 4OFOXOjO|O�O�O�O��O�O�O�O_�?GRI�`ΛDQ�?_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|� ���������0�B�T��oPREG �>�� f���Ə؏� ��� �2�D�V�h�z� ������ԟ���Z���$ARG_��D ?	���;���  �	$Z�	[�O�]O��Z�p�.�S�BN_CONFIOG ;��������CII_SA_VE  Z������.�TCELLSETUP ;��%HOME_I�OZ�Z�%MOVq_��
�REP�l�U�(�UTOBAC�Kܠ���FRA:\z� �\�z�Ǡ'`��z���n�INI�0�z���n�MESSAG���ǡC���ODE_D�������%�O�4�n�PAU�SX!�;� ((O>��ϞˈϾ� �����������*� `�N߄�rߨ߶�g�l ?TSK  w�Կ<׿q�UPDT+���d!�A�WSM_kCF��;���|'�-�GRP 2:�V?� N�BŰA�߾%�XSCRD1�1�
7� �ĥĢ ����������*��� ����r����������� 7���[�&8J\�n��*�t�GRO�UN�UϩUP_kNA�:�	t�n�_ED�17��
 �%-BCKEDT-�2�'LK�`���-t��z�q�q�z���2t1������q�k�(/��ED3/��/�.a/8�/;/M/ED4�/t/�)?�/.?p?�/�/ED5`??�?<?.�?8O�?�?ED6O�?�qO�?.MO�O'O9OED7�O`O_�O.�O8\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o�_�	-9o�oo%oCR _ 9]�oF�o��k� � NO_DE�L��GE_UN�USE��LAL_OUT �����WD_ABO�Rﰨ~��pITR�_RTN��|N'ONSk���˥�CAM_PARA�M 1;�!�
 �8
SONY �XC-56 234567890� ਡ@����?��( АP\�
���{����^��HR5q�̹��ŏR�57ڏ�Aff���KOWA S_C310M
�x�}̆�d @<� 
���e�^��П\ ����*�<��`�r��g�CE_RIA_UI�!�=�F��}�z� ��_�LIU�]���ꋐ<��FB�GP ]1��Ǯ��M�_�q�0�C*  �����C1��9��@Ҩ�G���CR�C]���d��l��s��R������[Դm��vꨰ������� +C����(������=�HE�`ONFI�ǰ�B�G_PRI 1�{V���� �ϨϺ����������CHKPAUS��w 1K� ,!u D�V�@�z�dߞ߈ߚ� �߾������.��R��<�b���O��x������_MOR��� �6��� 	 �����*��N�<�������?��qI?;�;����K���9�P���ça�-:���	�

��M���pU�ð��d<��,~��DB����튒)
mc:cpmidbg��f�:��p��:�¥�p�/� g �0�)�a� �s>��p���p�U�?Y�� \Ug��/���p�Uf��M/w�O/�
DEFg l��s)��< buf.txt s/�t/��ާ�)��	`�����=L�m��*MC��1��a��?43��1����t�īCz  B�HH�Co�C|���CqD���C���C��{iY
K�D���F.��F���E⚵F,�E�ٟ�K�F�N��IU��I?O��I<#I6�I�Y	��H,�$w�1���s�U��.�p�����1�BDw�M@x8��1eҨ����g@D�p@�0EYK�EX��EQ�EJP� F�E�F�� G��>^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE d��C
Q��;�(PG  B_<_��R�����	op6C4P�Y
s@ ]AQ�2s@�C�0B3�MaC{@@�*cw��UT�pFP?ROG %�z�o�oigI�q���v��ld�KEY_TBL � �&S�#� �	
��� !"�#$%&'()*+,-./01i��:;<=>?@A�BC� GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������vq���͓���������������������������������耇����������������������p`LCK�l4�p`��`STAT ��S_AUTO_DO����5�INDT_'ENB!���R�Q?��1�T2}�^�STO�Pb���TRLr`L�ETE��Ċ_S�CREEN ~�Zkcsc���U��MMENU �1 �Y  <�l�oR�Y1�[��� v�m���̟�����ٟ �8��!�G���W�i� �������ïկ��4� ��j�A�S���w��� ��迿�ѿ����T� +�=�cϜ�sυ��ϩ� ��������P�'�9� ��]�o߼ߓߥ���� ����:��#�p�G�Y� ����������$� ���3�l�C�U���y� ���������� ��	�VY)�_MANU�AL��t�DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�mg�(&/~&lMZ�IdPx�@P@#ONTIM6ه� d�`&��
�e�MOTNE�ND�o�RECO_RD 1(�[g2�/{�O��!�/k y"?4?F?X?�(`?�? �/�??�?�?�?�?�? )O�?MO�?qO�O�O�O BO�O:O�O^O_%_7_ I_�Om_�O�_ _�_�_ �_�_Z_o~_3o�_Wo io{o�o�_�o o�oDo �o/�oS�oL �o����@�� �+�yV,�c�u�� ������Ϗ>�P��� ��;�&���q���򏧟 ��P�ȟ�^������ I�[����� ���$��6�������jTO�LERENCwB����L�͖ C�S_CFG )��/'dMC:�\U�L%04d.'CSV�� c��/#[A ��CH��z� �//.ɿ��(S�R�C_OUT *���1/V�SGN� +��"��#��19-FEB-�20 16:00�017l�9:09�+ PQ�8�ɞ�/.��f�pa��m��PJP�Ѳ��VERSI�ON Y��V2.0.84,E�FLOGIC 1�,� 	:�ޠ=�ޠL��PROG_ENB��"p�ULSk' ����_WRSTJNK ���"fEMO_O�PT_SL ?	��#
 	R575/#=������0�B����TO  a�ݵϗ��V_F �EX�d�%��P�ATH AY�A�\�����5+IC�T�Fu-�|j�#egS��,�STBF_TTS�(�	d���l#!w�� MAU��z�^"�MSWX�.�<�(4,#�Y�/�
!J� 6%ZI~m���$SBL_FAU�L(�0�9'TDI�A[�1<�<� ����1234567890
��P��HZl~�� �����/ /2/�D/V/h/�� P� ѩ�yƽ/��6 �/�/�/??/?A?S? e?w?�?�?�?�?�?�?8�?�,/�UMP����3 �ATR��Ӝ1OC@PMEl�OOY�_TEMP?�ÈÓ3F���G�|DUN�I��.�YN_BR�K 2_�/�EMGDI_STA���]��ENC2_SC/R 3�K7(_ :_L_^_l&_�_�_�_0�_)��C�A14_�/�oo/oAoԢ�B�T5�K�ϋo~ol� {_�o�o�o'9 K]o����� ����#�5��/V� h�z��л`~�����ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T���x� ��������ү���� �,�>�P�b�t����� ����ο����(� f�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����:� �2�D�V�h� z������������ 
��.�@�R�d�v��� ����������� *<N`r��� ����&8 J\n������� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?��?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__No�ETMODE 1�6�5�Q 
�d�X
X_j_|Q�P�RROR_PROoG %GZ%�@���_  �UTABL/E  G[�?o�o)oRjRRSEV_NUM  �`WP�QQY`�Q�_AUTO_EN�B  �eOS�T_;NOna 7G[�Q}Xb  *��`���`��`��`d`+�`�o�o�o�dHIS�Uc�QOP�k_ALMw 18G[ �A��l�P+�ok} �����o_Nb�`  G[�a�R
��:PTCP_VER� !GZ!�_�$�EXTLOG_R�EQv�i\�S�IZe�W�TOL � �QDzr�{A W�_BWD�pp��xf́t�_DI��7 9�5�d�Tx�QsRֆSTEP���:P�OP_DO�v�f�PFACTORY_TUNw�dM�EATURE� :�5̀rQ�HandlingTool ��� \sfmE�nglish D�ictionar�y��rodu�AA Vis�� ?Master�����
EN̐nal?og I/O�����g.fd̐uto� Softwar�e Update�  F OR�m�atic Bac�kup��H596�,�groun�d Editޒ � 1 H5C_amera�F���OPLGX�ell�𜩐II) X�o�mmՐshw���c�om��co���\�tp���pane���  opl��t�yle sele{ct��al C���nJ�Ցonito�r��RDE��t�r��Reliab�𠧒6U�Diag�nos(�푥�55�28�u��hec�k Safety� UIF��Enh�anced Ro�b Serv%�q� ) "S�r�User Fr[������a��xt. DI�O �fiG� s�Ţ��endx�Er5r�LF� pȐĳ�r됮� ����  �!��FCTN Menu`�v-�ݡ����TP Inېf�ac�  ER �JGC�pבk� Exct�g��H�558��igh-wSpex�Ski1�?  2
P��?�~��mmunic'��ons��&�l�ur8�ې��ST Ǡ�^�conn��2���TXPL��ncr��stru����"�FATKAR�EL Cmd. �LE�uaG�545�\��Run-TiEnv��d
Q!���ؠ++�s)��S/W��[�L?icenseZ���� 4T�0�ogBo�ok(Syڐm)H54O�MAC�ROs,\�/Ofwfse��Loa��MH������r, �k�MechSto?p Prot����o lic/�Miв�Shif����ɒM�ixx��)���,e��S�Mode S�witch�� RM5W�Mo�:�.�֏ 74 ���g���K�2h�ulti�-T=�M���LN �(Pos�Regiڑ������d�>ݐt Fun�ǩ�q.�����Num~�<���� lne���>�� Adjup��|����  - W��Otatuw᧒T��RDMz�ot���scove �U�9���3Ѓ�u?est 492�*��o�����62;�S�NPX b ���8� J7`���Libr��J�48���ӗ�� �Ԅ�
�6O�� �Parts in_ VCCMt�32����	�{Ѥ�J99�0��/I� 2 �P��TMILIB���H���P�AcycD�L�
TE$sTX�ۨ�ap1S��Te����pkey���wգ�d���Unexceptx�motnZ���������є�� O8���� 90J�єSP CSXC<�f��Ҟ� Py�W9e}���PRI�>svr�t�men�� ��iPɰa������vGrid�play��v���0�)�H1�M-1�0iA(B201� �2\� 0\k�/�Ascii�lp�Т�ɐ/�Col���ԑGuar� 
d�� /P-�ޠ"K��;st{Pat ��!S�Cyc�҂�gorie��IF8�7ata- quҐ��� ƶ��mH5746��RL��am����Pb�HMI Deb3�(b����PC�~��Passwo+!n��"PE? Sp$��[���tp��� ve�n��Tw�N�p�Y�ELLOW BO�E	k$Arc��vi�s��3*�n0We{ldW�cial�47�V#t�Op����Y1y� 2F�a듏portN�(�p�T�1�T� �� ��xYy]�&TX��tw��igj�1� b� c�t\�JPN A�RCPSU PR���oݲOL� Sup�2fil� &PA�ɰאcro�� "�PM(����O$SS�� eвtex�� �r���=�t�ss�agT��P��P`@�Ȱ�锱�rtW�p�H'>r�dpn���n1
t�!� �z ��ascbin�4psyn��+Aj��M HEL�N�CL VIS P�KGS PLOA�`�MB �,�4V�W�RIPE G�ET_VAR F�IE 3\t��F�L[�OOL: A�DD R729.�FD \j8'�C4sQ�QE��DVvQ��sQNO WTWT�E��}PD  Dpx��biRFOR ���ECTn�`��AL�SE ALAfPC�PMO-130 � M" #h�D:� HANG FRcOMmP�AQfr���R709 DRA�M AVAILCHECKSO!��sQVPCS SU�@LIMCHK Q �+P~dFF POS���F�Q R593�8-12 C�HARY�0�PRO�GRA W�SA�VEN`AME�P.�SV��7��$En�*��p?FU�{�TRC�|� SHADV0UPDAT KCJ�>�RSTATI�`�P� MUCH y�1���IMQ MOT�N-003��}�R�OBOGUIDE? DAUGH�a���*�tou����I�u Šhd�ATH�P>epMOVET�ǔ�VMXPACK �MAY ASSEsRT�D��YCLfq�TA�rBE CO�R vr*Q3rAN��pRC OPTI�ONSJ1vr̐P�SH-171Z@x�tcǠSU1�1Hp0^9R!�Q�`_T�P���'�j�d{tby� app wa 15I�~d�PHI���p�aTEL�MXS�PD TB5bLu d1��UB6@�qENJ`[CE2�61��p��}s	�may n�L0� R6{�R� �R�traff)�� k40*�p��fr���sysvar scr J7��cj`'DJU��bH V���Q/�PSET EsRR`J` 68����PNDANT S�CREEN UNGREA��'�J`D�p�PA���pR`IO� 1���PFI�pB��pGROUN�PD���G��R�P�QnRSV�IP !p�a�PDI�GIT VERSl�r}BLo�UEWϕ? P06  �!��MAGp�abZV��DI�`� SSU�E�ܰ�EPLA�N JOT` DEIL�pݡ#Z�@D͐�CALLOb�Q p�h��R�QIPNDIMG�R71�9��MNT/�PE�S �pVL�c��H�ol�0Cq���tPG�:�`C�M�can�Π��pg.v�S:� 3D mK�vi/ew d�` �p���ea7У�b� of� �Py���ANNO�T ACCESS� M��Ɓ*�t4s� a��lok��FWlex/:�Rw![mo?�PA?�-������`n�pa SN�BPJ AUTO-�06f����TB��P�IABLE1q 6�36��PLN: �RG$�pl;pNWF�MDB�VI���tWOIT 9x�0@o���Qui#0�ҺPN wRRS?pUSB���� t & rem�ov�@ )�_��&A�xEPFT_=� 7�<`�pP:�OS-�144 ��h s8�g��@OST� �� CRASH D�U 9��$PھpW� .$��LOGIN��8&�J���6b046 iss?ue 6 Jg��: Slow ��st��c (Ho�s`�c���`IL`I�MPRWtSPOT�:Wh:0�T�ST�YW ./�VMGR��h�T0CAT��hos��E�q���� �O�S:+pRT)U' k�-S� ����E:��pv@�2�� 't\hߐ��m ��gall��0�  $��H� WA͐��3 ?CNT0 T�� �WroU�alar1m���0s�d � �0�SE1���r R{�O�MEBp���K� 5�5��REàSEst���g     ��KANJI�n�o���INISITALIZ-p�dn1cweρ<��dr��� lx`�SCII� L�fails� w�� ��`�YS�TEa���o��Pv� �IIH���1W�Gr}o>Pm ol\wp�Sh@�P��Ϡn �cflxL@АWR=I �OF Lq��p�?�F�up��de�-rela�d �"APo SY�ch��Abetwe:0I�ND t0$gbD�O���r� `�G�igE�#operoabilf  PAb�Hi�H`��c�lea=d�\etf�Ps�r�OS 030�&�: fig��GLAA )P ��i��7Np_ tpswx�B��If�g�������5aE�a EXCE�#dU�_�tPCLOSޡ�"rob�NT
dpFaU�c�!����PNIO V75�0�Q1��Qa��DB ��P M�+P�Q;ED�DET��-�� \rk��ONLwINEhSBUGI`Q ߔĠi`Z�IB�S� apABC JOARKYFq� ��N�0MIL�`� R�p�NД �p0GAR���D*pR��P�"! jK�0cT�P�Hxl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P�`nWIBPK05�!�FȐB/��BUS�Y RUNN�� !"�򁐈��R-p�sLO�N�DIVY��CUL��fsfoaBW�p���`30	V��ˠIT`ެa505.�@OF�UNEX�P1b�a�f�@�E��SVE;MG� NMLq� �D0pCC_SAFQEX 0c�08"qD ��PET�`N@�#J87����RsP�A�'�M�K�`K�H GUNCHG۔/MECH�pMc� =T�  y, g@�$� ORY LEA�KA�;�ޢSPE�m�Ja��V�tGRI�ܱ�@�CTLN��TRk�FpepR�j�50�EN-`IN�����p �`�Ǒk!Ɯ�T3/dqo�ST�O�0A�#�L�p  �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`DU���aO�supk�t4 d� P�F� Bnf�Q~�PSVGN-1���V�SRSR)J�U�P�a2�Q�#D�q �l O��QBRKCTR5Ұ�|"-�rp�<pc�j!INVP�D ZO� ��T`h#x�Q�cHset,|D<��"DUAL� w��2*BRVO117 A]�TNѫt�+bTa2473��q.?���r�{1 009.�fd8�y`j604�.\P-�`hancZ�U� F��e8�'�  ��npJtPd!�q��`��� 5h596p�!5d�� "p �P�P�Q�0�P2�p�A�� \P��R(}\\PeJ� aʰI���E���1��p� j  �� ,e��Dp� �A�Ap\P�q 5 sig��a��"AC;a��p
�bCe\Pb_p���.pc]l<bHbcb_circ~h<n�`tl1�~`\P`o�d\PX�b]o2�� �cb�c��i\P�jupfrmp�d\P�o�`exe�ax�oFd\Ptped}o���u`�cptlibxz\P�lcr�xr\P�\�blsazEd\P_fm�}gc\P�x���o�|sp�o�mc(��ob_jzop�u6�wQf��t��wms�1q���sld�)��jmc�o\�n��nuhЕ��|cst�e��>�pl�q�p�iwck���uv�f0uߒ��lvisyn�CgaculwQ�
E `RFciV\Pq�iP��Data A�cquisi��n<ZU�SR631`��T}R�QDMCM ��2�P75H�1�P5k83\P1��71��k59`�5�P57<P \P�Q����(���Q̖�o p\P!da�q\�oA��@��y ge/�etdms�?"DMER"؟,�GpgdD���.�m��8�-��qaq.<᡾F\Pmo��h���f{��oR503��MACROs, SksaCff�@lR���03�SQR�Q(��Q6��1�Q9ӡ�R�ZSh��P\P�J643�@7ؠ6X�P�@�PRS�@����e �Q�UС PIK��Q52 PTLC��W��\P3 (��p/O��!�Pn ��\P5��03\sf�mnmc "MNCMCq�<��Q��\$AcX�FM���ci,� ��X����cdpq+�
�sk�SK�\P�SH560,P��,��y�refp "R#EFp�d�A�j\P	�of�OFc�<gy�to�TO_���������+je�u>��caxis2�\P�E�\�e�q"ISD�Tc��]�prax ��MN��u�b�isde܃h�\�iR�\P! isbaskic��B� P]�ޔQAxes�R6p������.�(Ba�Q�ess��\P����2�D�@�z�atis���(�{�����4~��m��FMc�u�x{�
ѩ�MNIS�� ݝ����x����ٺ��jW75��Dev�ic�� Inte�rfac�RȔQJ�754��� \P�Ne`��\P�ϐ2��б����dn� "�DNE���
tpodnui5UI��ݝ	bd�bP�q_rsofOb
?dv_aro��u�����stchkc��z	 �(}�onl��G!ff L+H�J(��"l"/��n�b��z�haSmp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!2���xpc_2pcch=m��CHMP_�|8бpevws��2�ΌpcsF��#C �Sen\Pacro0�U·�-�R6�Pd�@\Pk�����p��gT�L��1d M�2`��8��1c4ԡ�3 qem��GEM,\i(��Dgesnd�5���H0{�}Ha�@sy���c��Isu�xD��Fmd ��I��7�4���u���AccuCal�P��4t@��ɢ7ޠB0���6+6f�6��9!9\aFF q�S(�U��2�
X�p�!Bd�ѳcb_�SaUL�� � �t@?�ܖto���otplus\tsrnغ�qb�W�p��t���1��To�ol (N. A�.)�[K�7�Z�(P��m����bfcllst@k94�"K4p���qtpap� �"PS9H�stpswo��p�L7��t\�q����D�yt5� 4�q��w�q��t@�Mz�uk��rkey�����s��}t�sfe7atu6�EA��t@cf)t\Xq�����df�h5���LRC0�md�!�587���a�R�(����2V��8lc?u3l\�pa3}@H�&r-�Xu���t,�t@�q "�q�Ot��~ ,���{�/��1c�}����y�p�r��5����S�XAg�-�y���Wj�874�- iR�Vis���Queu�t@Ƒ�-�6�1$���(����u����tӑ����
�tpv�tsn "VTS�N�3C�+�t@v\pR�DV����*�prd�q\�Q�&�vst�k=P������nmx&_�դ�clrqν���get�TX��Bd���aoQϿ�0q�str�D[t@��t0�p'Z����npv��@�enlIP0��D!0x�'�|���sc ߸��tvo/��2�q���vb����q����!���h]��(� Control�PRAX�P5��5�56�A@59�P5-6.@56@5A��J69$@982 �J552 IDVR7�hqA���16�Hx���La�� ���Xe�frlparwm.f�FRL��am��C9�@(F �����w6{���A���QJ643�t@5}0�0LSE
_p�VAR $SGS�YSC��RS_UNITS �P�2�4�tA�TX.$VN�UM_OLD 5`�1�| {�50+��"�` Funct ���5tA� }��`#@�`E3�a0�cڂ��9����@H5נt@�P���(�A����۶}�����ֻ}��bPR�b�߶~ppr4�TP�SPI�3�}�r�10�#;A� t�
`���1���96�����%C�� Aف��J�bIncr�	����\�`��1o5qni4�MNINp	�t@����!��Hour_  � 2�21 �A�AVM���0 ���TUP ��?J545 ���6162�VC�AM  (��CLIO ���R6�N2�MSC� "P ��STYL�C�28�~ 13\�NRE� "FHRM S�CH^�DCS}U%ORSR {b��04 �E�IOC�1 j 5742 � os| �? egist��Ի��7�1�oMASK�934"�7 ��OCO ���"3�8��2���� 0 HB��ڢ 4�"39N� R�e�� �LCHK�
%OPLG%��3�"%MHCR.%MCd  ; 4? ��6 d�PI�54�s� D[SW%MD� pQ�K!637�0�0p"�Y1�Р"4 �6<2?7 CTN K � +5 ���"7��<2�5�%/�T�%FRD�M� �Sg!��9�30 FB( NBA��P� ( HLB  7Men�SM$@jB�( PVC ��290v��2HTC�C?TMIL��\@?PAC 16U�hA�J`SAI \@ELN���<29s�UE�CK �b�@FRM� �b�OR���I�PL��Rk0CSXsC ���VVFna}Tg@HTTP �N!26 ��G�@~obIGUI"%�IPGS�r� H863 qb�!�07r�!�34 �r�84 �\so`! Qx`CC3� Fb�21�!969 rb!51 ���!S53R% 1!s3!���~�.p"9js V{ATFUJ775"���pLR6^RP�WS�MjUCTO�@xT5�8 F!80���1X�Y ta3!770 ���885�UOL�  GTSo
�{` L�CM �r| TSS��EfP6 W�\@CPgE `��0VR� �l�QNL"��@00�1 imrb�c3� =�b�0���0�`6� w�b-P- R-��b8n@5EW�b9 �Ґa� ���b�`ׁ~�b2 2000���`3��`4*5�`5 !�c�#$�`7.%�`�8 h605? U�0�@B6E"aRp76� !Pr8 t�a�@�tr2 iB/d�1vp3�vp5 ȂRtr9Σ�a4@-pN�r3 F��r5&0�re`u��r7 ��r�8�U�p9 \h7�38�a�R2D7�"�1f��2&�7<� �3 7iC���4>w5Ip�Or60� C�L�1bEN�4 I�pyL�uP��@N�&-PJ8�N�8NeN�C9 H�r`�E�b7]�|���8�ВࠂG9 2��a`0�q�Ђ5�%U097 �0��@1�0���1� (�q�3 5R ���0���mpU���0�0�7*�H@(q��\P"RB6�q124�b;��@���@�06� x�3 pB�/x�u ��x�6 H606�a1� ��7 6 ���p��b155 ����7>jUU162 ��3 g��4*�65 2e "_��P�4#U1`���B1���`=0'�174 �q���P�E186 R L��P�7 ��P�8&��3 (�90 B�/�s191����@2s02��6 3���A�RU2� d��O2 b2h`��4��b��2�4���19v RQ�2��u2d�Tpt)2� ��H�a2hP�$2�5���!U2�p�p"
�2�p��@5�0-�@��8 @�9��T�X@�� �e5�`rb	26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0@�gqGA���a�52ѐ�Ḳ6�6�0ہ5� ׁ2��84�E��9�EU5@ٰE\�q5hQ`S�2ޖ5�p\w�۲�pJ �4-P��5�p1\t�H�-4��PCH�7j��phiw�@��P�x��?559 ldu� P �D���Q�@�������A �`.��P>��8�g581�"�q58�!�AM۲T�A iC�a589��@�x���F�5 �a��12׀ 0.�1���,�2�����,�!P\h8��Lp ���,�7��6�084�0\t� "T20C}A��p��{��sran��FRA�� �Д�е���A%�� �ѹ�Ҁ�����(�� ��Ѐ���З���������р����$�G��1��ը��������� ,e�`�q�  �����`6�4��M��iC/50T-H������*��)p46��� C��xN����m75s֐�� Sp�ѯb46���v����ГM-7�1?�7�З����4A2������C��-��F��70�r�E��/h����O$��rlD���c7c7C� q��Ѕ���L��/���2\imm7c7�g������`���(��e�����"� �������a r��&c�T,�Ѿ�"��,��� ��x�Ex�m7�7t���k���5������)�iC��-HS-� B
_� >���+�Т�7U�]P���Mh7�s��a7������-9?�?/260L_������Q�������]�9pA/@���q�S�х��^�h621��c��92������.�)92c0�g$�@������)$��5$���pcylH"O"
�21�8��t?�350� ���p��$�
�� F�350!���0�x�9�U/0\m9��M9A3��4%�� s�3M$��X%u<���"him98J3����� i d�"m4~��103p�� �Ӏ�h�794̂�&R���H �0����\���g�5A ���Ԝ��0���*2� �00��#06�а�Ճ�է!07{r  ��������kЙ@�����EP�#�������?��#!�;&0s7\;!�B1P��@�A��/ЁCBׂ2�!��:/��?�ҽCD25�L����0�"l�2BL
#��B��\20�2_�r�re� ��X��1��N����A@��z��`C�pU��`�04��Dy	A�\�`fQ��s�U���\�5  ��� p�Dp���<$85���+P=�ab1l�1LT��lA8�!uDnE(�.20T��J�1 e�bH85���b�Հ�5[�16Bs��������d2��x��m6t!`Q����b�ˀ���b#�(�6iB ;S�p�!��3� ���b�s��-`�_�W80�_����6I	$�X5�1�U85��R�p6S����/�/+q�!@�q��`�6o��5m[o)�m6sW��Q�|�?��set06p h��3%H�5��10p$@����g/�JrH��?  ��A��856����F�� ���p/2��� ��܅�✐)�5��̑v�𘜐(��m6��Y�H�ѝ̑m�6�Ҝ��ae6�DM����-S�+��H2�����Ҽ� � �r̑��✐��l���p1���F����2�\t6h T6H����Ҝ�'Vl ���ᜐ�V7ᜐ/�(���;3A7��p ~S��������4�`堜��V���!3��2��PM[��%ܖO�chn��vel5���8�Vq���_arp#���̑�.���2l_h�emq$�.�'�6415���5���?����F�����5g�L�ј�[���1��𙋹1<����M7NU�Р���eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h������ u���㜐��ZS0�!ܑ4���M-����S�$̑�ք �� 0���<�����07shJ�H�v�À�sF� �S*󜐳���̑���vl�3�A�T�#��Q�0��Te��q�pr����T@75j�5�dd�̑ 1�(UL�&�(�,���0��\�?���̑�a�� ,e����a�eD�w�2��(�	�2�C��A/���\�+p�<����21 (ܱ�CL S����B̺@��7F���?�<�lơ1L����c� ���u19�0����e/q���O���9�K��r9 (��,�Rs�ז�5�<G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O���M1!41w���2T@� _std��G�y�� �ң�H� jdgm����w0\� �1L� ��	�P�~�W*�b���t 5������3�,���E{���d���L��5\L��3�L�|#~���~!���4�#��O����h�L6A�������a2璥���44������[6\j4s ��·���#��ol�E"w�8Pk�����?0x j�H1�1Rr�>��]�2a�2Aw�P ��	2��|41�8��ˡ��@{� �%�A<��� +� ?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R�� ˑb�W���Fs���) �ѐ�!���a�1�����5��16�16C���C����0\imBQ��d����b��\Be5�-���DiL����O�_�<ѠPEtL �E�RH�ZǠPgω�am1l��u���̑�b@�<����<�$�T� ̑�F����Ȋ�DpbĜ�X"��hr��pĻ ��Dp���9��0\� j971\�kckrcfJ�F�s�����c��e "CTME�r���ɛ�|�a�`main.[�8�g�`run}�_vc�#0�w�1Oܕ�_u����bctme���Ӧ�`ܑ�j73�5�- KARE�L Use {�U���J��1���p� Ȗ�9�B@���L�9��7j[�atk208 "K��(Kя��\��9��a���̹����cKRC4�a�o ��kc�qJ� &s�����Grſ�fs�D��:y��s��A1X\�j|хrdtB�, L��`.v�q�� �spǑIf�Wfj52��TKQuto Seut��J� H5K7536(�932���-91�58(�9�BA��1(�74O,A$�(TCP Ak���/�)Y� �\tpqtool.v���v���! con�re;a#�Cont�rol Re�b{le��CNRE(� T�<�4�2���D�)���NS�552��q(g�� (򭂯4X�cOux~�\sfuts�UTS`�i�栜���At�棂��? 6�T�!�SA OO+D6���������,!��6c+� igt�t6i��I0�T�W8 ���la��vo58�o�bFå򬡯i��Xh��!Xk�0Y!8�\m6e�!6EC���v��6���������<16�A���A�6s����U�g�T|�,����r1�qR����Z4�T�����,#�eZp)g����<ONO0���uJ��tCR;��F<�a� ,e��f���prdsuchk� �1��2&&?���t��*D%$�r(�✑ �娟:r��'�s�qO��<scrc�C�\At�trldJ"o��\�V����Pay�lo�nfirm�l�!�87��7��A�3ad�! �?@ވI�?plQ��3���3"�q��x pl��`���d7��l�calC�uDu���;���mov�����initX�:s8O��a8�r4 ��r67A4|��e Genera#tiڲ���7g2q$g R� (S�h��c ,|�bE��$Ԓ\�:�"���4��4�4�. sg��5�F$d6"�e;Qp "SHA�P�TQ ngcr pGC�a(�&"� ���"GDA¶��r�6�"aW�/�$d�ataX:s�"tp�ad��[q�%tput;a__O7;a�o8�1�yl+s�r�?�:�#$�?�5x�?�:c O�:Ay O�:�IO�s`O%g�qǒ�?�@0\ۜ�"o�j92;!�Pp�l.Collis�QSkip#��@5� �@J��D��@\ވ�C(@X�7��7�|s}2��ptcls�#LS�DU�k?�\_� ets�`�< �\�Q��@���`dcKLqQ�FC;��J,όn��` (��4eN����T�{���' j(�c�����/IӸaȁ<��̠H������зa�e\mcc�lmt "CLM��/��� mate\v��lmpALM�?>p7qmc?�����2vm�q��%�3s��_�sv90�_x_msu�2L^v_� K�o��{in�8(3r<�c_logr��r�trcW� �v_3�~yc��d�<�ste��der$c;Ce� Fiρ��R��Q�?�l�enter߄|��(�Sd��1�TX�+fZK�r�a99sQ9+��5�r\tq\� _"FNDR����STDn$�LANG�Pgui��D⠓�S������csp�!ğ֙uf䟀ҝ�s����$�����e +�=����������������w�H�r\fn�_�ϣ��$`x�tcp�ma��- TCP������R638 aR�Ҡ��38��M7p,���Ӡ�$Ӡ��8p0Р�VS,�>�tk��99�a��B3���P�զԠ��D�2�����UI��t���hqB���8���������p���re8�ȿ��exe@4π��B���e38�ԡG�r�mpWXφ�var @�φ�3N�����v�x�!ҡ��q�R�BT $cOP�TN ask E�0��1�R MAS�0�H593/�96g H50�i�480ԅ5�H0��m�Q�K(��7�0�g�Pl�h�0ԧ�2Ҧ�DP���@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`am��b��7�.f���u�d��r��splayD�E���1wПUPDT Ub��8o87 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60�q��B����qs�can��B���aAd@�������q`� �䗣�#��К�`2�� vlv��Ù�$�0>�b���! S���Easy/К�Ut�il��룙�511# J�����R7 ���Nor֠��inc�),<6Q�� �`c��"4�[���986(FVRx So����q�nd6����P��4� a\ (��
  ������"�d��K�bdZ����men7���- Me`tyFњ�Fb��0�TUa�577?i3R��\�5�au?��!� n����f������l\m�h�Ц�űE|h#mn�	��<\O�$��e�1�� l!���y��Ù�\|p�����B���Ћmh �@��:.aG!�� �/�t�55�6�!X��l�.us��Y/k)eOnsubL���eK�h�� �B\1;5g?�y?�?�?D��?*rmx�p�?Ktbox O�2K|?�G��C?A%d�s���?�P"�!�  �TR��/��P�T6@�`��U�P�V�P�Ue�P0�U�PO��\3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q�� �R?Ă�Q3t.�P׀#al��P+OP7517��IN0a��Q(}g��PESTf3ua�PB�l�ig��h�6�aq��P �� ,e��` y n�0mbumpPn�Q969g�69�Qq��P0�baAp�@Q� BOX��,>v�che�s�>vet�u㒣=wffse�3���]�;u`aW��:zol�sm<ub`�a-��]D�K�ibQ��c����Q<twaǂ t�p�Q҄Taror? Recov�b�9O�P�642�����a�q��a⁠QErǃ�Qry��`�P'�T�`�aar������	{~'�pak971��71��m���>��`jot��PXc��C�1�madb -�ail���nag���b�QR6�29�a�Q��b�P�  �
  |�P��$$CL[q? ����������$�PS_�DIGIT���"�!�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ��������*璬1:PR�ODUCT�Q0\_PGSTK�bV,�n�99�����$FEAT?_INDEX��~�������ILECOMPW ;��)���"��SETUP2� <����  N !�_�AP2BCK 1�=�  �)�}6/E+%,/i/� �W/�/~+/�/O/�/ s/�/?�/>?�/b?t? ?�?'?�?�?]?�?�? O(O�?LO�?pO�?}O �O5O�OYO�O _�O$_ �OH_Z_�O~__�_�_ C_�_g_�_�_	o2o�_ Vo�_zo�oo�o?o�o �ouo
�o.@�od �o���M�q ���<��`�r�� ��%���̏[����� ��!�J�ُn������� 3�ȟW������"��� F�X��|����/��� ֯e������0���T� �x������=�ҿ� s�ϗ�,ϻ�9�b��� P/ 2) �*.VRiϳ�!�*�����������PC�7�!�FR6:"�c��χ��T��߽�Lը��ܮxx���*.F��D>� �	N�,�k���<���STM ������Qа���!�i�Pendant �Panel���H ��F���4������GIF�������u�8���JPG&P���<����	P�ANEL1.DT��������2�Y�G��
3w�����//�
4�a/�O/�//�/�
TPEINS.XML�/����\�/�/�!C�ustom To�olbar?��PASSWORD�/�FRS:\�R?? %Pas�sword Config�?��?k? �?OH�6O�?ZOlO�? �OO�O�OUO�OyO_ �O�OD_�Oh_�Oa_�_ -_�_Q_�_�_�_o�_ @oRo�_voo�o)o;o �o_o�o�o�o*�oN �or��7�� m��&���\�� ���y���E�ڏi��� ���4�ÏX�j����� ���A�S��w���� �B�џf�������+� ��O���������>� ͯ߯t����'���ο ]�򿁿�(Ϸ�L�ۿ pς�Ϧ�5���Y�k�  ߏ�$߳��Z���~� ߢߴ�C���g���� ��2���V����ߌ�� ��?����u�
���.� @���d������)��� M���q�����<�� 5r�%��[ �&�J�n ��3�W�� �"/�F/X/�|// �/�/A/�/e/�/�/�/ 0?�/T?�/M?�??�? =?�?�?s?O�?,O>O �?bO�?�OO'O�OKO �OoO�O_�O:_�O^_ p_�O�_#_�_�_Y_�_�}_o�_�_Ho)f�$�FILE_DGB�CK 1=���5`��� ( �)
SU�MMARY.DG<Ro�\MD:�o�o�
`Diag Summary�o��Z
CONSLO�G�o�o�a
J�a�Console �logK�[�`MEMCHECK@�'�o�^qMem�ory Data|��W�)�qHADOW����P��sShado�w Change�sS�-c-��)	FTP=��9�����w`qmment� TBD׏�W0<��)ETHERNET̏�^�q�Z���aEthern�et bpfigu?ration[��P~��DCSVRFˏp��Ïܟ�q%��� verify �allߟ-c1PY=���DIFFԟ���̟a��p%��d�iffc���q��1pX�?�Q�� �����X��CHGAD��¯ԯi��px��� ���2`�G�Y��� ��� �GD ��ʿܿq��p������FY3h�O�a���� ��(�GD ������y��p�ϡ��0�UPDATE�S.�Ц��[FR�S:\�����aU�pdates L�ist���kPSRBWLD.CM.���\��B��_pPS�_ROBOWEL ���_����o��,o!� 3���W���{�
�t��� @���d�����/�� Se�����N �r� =�a �r�&�J�� �/�9/K/�o/� �/"/�/�/X/�/|/�/ #?�/G?�/k?}??�? 0?�?�?f?�?�?O�? OUO�?yOO�O�O>O �ObO�O	_�O-_�OQ_ c_�O�__�_:_�_�_ p_o�_o;o�__o�_ �o�o$o�oHo�o�o~o �o7�o0m�o�  ��V�z�!� �E��i�{�
���.� ÏR����������.� S��w������<�џ `������+���O�ޟ H������8���߯n�����$FILE�_��PR����������� �MDONLY� 1=4�� 
 ���w�į��� ��ѿ�������+Ϻ� O�޿sυ�ϩ�8��� ��n�ߒ�'߶�4�]� �ρ�ߥ߷�F���j� ����5���Y�k��� ����B�����x�� ��1�C���g������ ,���P����������?��Lu�VIS�BCKR�<�a�*�.VD|�4 F�R:\��4 �Vision V?D file�  :LbpZ�#� �Y�}/$/�H/ �l/�/�/1/�/�/ �/�/�/ ?�/1?V?�/ z?	?�?�???�?c?�? �?�?.O�?ROdOO�O O�O;O�O�OqO_�O *_<_�O`_�O�__%_��_�MR_GRPw 1>4�L�U�C4  B�P	� ]�ol`��*u���R�HB ��2 ���� ��� ���He�Y�Q`orkb Ih�oJd�o�Sc�o�o�L�SJe�I���F�5U�aQ��0��o��oD�	�G��aE�9��o9cݨ>���F}@M$G@Q���lr?@N��@O�K}E�� F@ �r��d�a}J��NJ�k�H9�H�u��F!��IP�s}?�`�.�9�<9��896C'�6<,6\b��}A+~�BS/��B� JA���?B#�VA�4�. �"7�A��_B|EDA����A�a�A������,.��PA� ����|�ݏx���%������4,AX4�P@#x�@ICm4���j�����ǟ ���֟��!��E�`�r�UBH�P p�a`�M�H��o"K�豯ï�T
6�PS@�PS�`˯�o�o�B��P5���@�33@���4�m�T��UUU��U�~w�>u.�?!x��^��ֿ���3��=�[z�=�̽=�V6<�=�=�=$q��~���@8�i7�G��8�D�8@9!�7���@Ϣ���:t�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p���������.��� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__>���  DE_�Hly_�\@@m_B�=��vR/��I�O�SMT
�G�SUoo&o�RHOSTC�19H�I� ��zM�SM�l[�bo�	127.�0�`1�o  e �o�o�o#z�oF�Xj|�l60s	a�nonymous��������(ao�&�&��o� x��o������ҏ�3 ��,�>�a�O���� ������Ο�U%�7�I� �]����f�x����� ���ү����+�i� {�P�b�t�������� ����S�(�:�L� ^ϭ�oϔϦϸ���� ��=��$�6�H�Zߩ� ��Ϳs���������� � �2���V�h�z�� �߰���������
�� k�}ߏߡߣ���߬� ��������C�*< Nq�_����� �-�?�Q�c�eJ�� n������ �/"/E�X/j/|/ �/�/�%'/? [0?B?T?f?x?��? �?�?�?�??E/W/,O�>OPObO�KDaENT� 1I�K P!�?�O   ��O�O �O�O�O#_�OG_
_S_ ._|_�_d_�_�_�_�_ o�_1o�_ogo*o�o No�oro�o�o�o	�o -�oQu8n� �������#� �L�q�4���X���|� ݏ���ď֏7���[����B�QUIC�C0��h�z�۟��1 ܟ��ʟ+���2,����{�!ROUT�ER|�X�j�˯!�PCJOG̯���!192.16?8.0.10��}GNAME !�J!ROBOT��vNS_CFG 1�H�I ��Auto-st�arted�$FTP�/���/�?޿ #?��&�8�JϏ?n� �ϒϤ�ǿ��[����� �"�4ߵ&�������� ��濜���������� '�9�K�]�o���� ����������/�/�/ G���k��ߏ������� ������1T��� Py�����"� 4�	H-|�Qcu �VD���� /�;/M/_/q/�/� ���/
/�/>?%? 7?I?[?*/?�?�?�? �/�?l?�?O!O3OEO �/�/�/�/�?�O ?�O �O�O__�?A_S_e_ w_�O4_._�_�_�_�_ oVOhOzO�O�_so�O �o�o�o�o�o�_ '9Kno�o��� ��o*o<oNoP5� �oY�k�}�����pŏ ׏����0���C�U��g�y���_�T_ER�R J;�����P�DUSIZ  j��^P����>ٕ?WRD ?z����  guest���+�=��O�a�s�*�SCDMNGRP 2Kz�wÐ���۠\��K�� 	�P01.14 8~�q   y���B   � ;����{ ������������������?�����~ �ǟ�I�4�m�X�|���  i  ��  
���� �����+�������
���l��.x����"�l�ڲ۰s�d����|���_GROU��]L�� ��	���۠07K�QUPD'  ���PČ��TYg�����T�TP_AUTH �1M�� <!iPendan����<�_�!K?AREL:*�����KC%�5�G���VISION �SETZ���|�� Ҽߪ��������� 
�W�.�@��d�v���CTRL N��軡���
�F�FF9E3����FRS:DEFA�ULT�FA�NUC Web �Server�
 ������q��������������WR_CONFIG O��� ���IDL_CPU_PC"���B��= �BH#MIN.�B?GNR_IO���� ���% NPT_S_IM_DOs}�TPMODNTO�Ls �_PRT�Y�=!OLNK 1P����'9K]o�MA�STEr �����O�_CFG��UO�����CYCLE����_ASG s1Q���
 q 2/D/V/h/z/�/�/�/ �/�/�/�/
??y"NUM���Q��IPCH��£R?TRY_CN"�u<���SCRN��擊��� ����R����?��$J�23_DSP_E�N�����0OB�PROC�3��J[OGV�1S_�@��?8�?�';ZO�'??0CPOSRE�O�KANJI_@�Ϡu�A#��3T ����E�O�ECL_�LM B2e?�@EYL_OGGIN��������LANGU�AGE _�=e� }Q��LG�2YU����� �x������PC � �'�0�����M�C:\RSCH\�00\˝LN_D?ISP V���0����TOC�4�Dz\A�SOGB?OOK W+��`o���o�o���Xi��o�o�o�o�o~}	x(y��	ne�i��ekElG_BUF/F 1X���}2����Ӣ��� ���'�T�K�]��� ��������ɏۏ����#�P��ËqDCS� Zxm =���%|d1h`���ʟܟ|�g�IO 1[+G �?'����'� 7�I�[�o�������� ǯٯ����!�3�G� W�i�{�������ÿ׿z�El TM  ��d��#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝߜ�t�SEV�0m.�TYP�� �0�$�}�ARS"�(_|�s�2FL 1\��0���������0�����5�TP<P����DmNGNA�M�4�U�f�UPSF`GI�5�A�5s��_LOAD@G �%j%@_M�OV�u����MAXUALRMB7�P8 ��y���3�0]&q
��Ca]s�3�~��� 8@=@^+ �Z�v	��V0+�P1�A5d�r���U����� �E(iTy� ������/ / A/,/Q/w/b/�/~/�/ �/�/�/�/??)?O? :?s?V?�?�?�?�?�? �?�?O'OOKO.OoO ZOlO�O�O�O�O�O�O �O#__G_2_D_}_`_ �_�_�_�_�_�_�_o 
ooUo8oyodo�o�o �o�o�o�o�o�o-���D_LDXDIS�A^�� �MEMO�_APX�E ?��
 �0y� ���������ISC 1_�� �O����W�i� ����Ə�����}� �ߏD�/�h�z�a��� ����������� @���O�a�5������� �����u��ׯ<�'� `�r�Y������y�޿ �ۿ���8Ϲ�G�Y� -ϒ�}϶ϝ�����mπ����4��X�j�#�_MSTR `��~}�SCD 1as}�R���N�������� 8�#�5�n�Y��}�� �����������4�� X�C�|�g��������� ������	B-R xc������ �>)bM� q�����/� (//L/7/p/[/m/�/ �/�/�/�/�/?�/"? H?3?l?W?�?{?�?�?��?n�MKCFG �b���?��LT�ARM_�2cRu;B �3Wp|TNBpMETPUOp��2����NDS?P_CMNTnE@8F�E�� d���N��2A�O�D�EPO�SCF�G�NPS�TOL 1e-�4=@�<#�
;Q�1 ;UK_YW7_Y_[_m_�_ �_�_�_�_�_o�_o Qo3oEo�oio{o�o�a��ASING_CH�K  �MAqODAQ2CfO�7J�e�DEV 	Rz	�MC:'|HSI�ZEn@����eTA�SK %<z%$�12345678�9 ��u�gTRI�G 1g�� l<u%���3����>svvYPaq��kE�M_INF 1h�9G `�)AT&FV0�E0(���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ���ڄH�� ����G�ֈAO�w� 2�������џ ���� ����͏ߏP��t��� ����]�ί����� (�۟�^��#�5��� ��k�ܿ� ϻ�ů6� �Z�A�~ϐ�C���g� y��������2�i�C� h�ό�G߰��ߩ��� �ϫ��������d�v� )ߚ��߾�y����� ���<�N��r�%�7� I�[������9�& ��J[�g��>�ONITOR�@G� ?;{   	?EXEC1�3�U2�3�4�5�T�p�7�8�9�3�n�R�R�R RRR(R@4R@RLR2YU2e2q2}2�U2�2�2�2�U2�3Y3e3���aR_GRP_SOV 1it��q(�a���C?BPR��A4�>%���gYw>rﳌ"}~q_DCd~�1P�L_NAME �!<u� �!D�efault P�ersonali�ty (from� FD) �4RR�2k! 1j)TE�X)TH��!�AX d�?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�Ox2-?�O�O�O__@0_B_T_f_x_�b<�O �_�_�_�_�_�_o o�2oDoVoho&xRj" �1o�)&0\�b,� �9��b�a �@D�  �a?�ľc�a?�`�a�aA'�6�ew;�	�l�b	 ��xJp���`�`	p �<w �(p� �.r�� K�K ���K=*�J����J���JV�`�kq`q�P�x��|� @j�@T;;f�r�f�q�a�crs�I�����p���p�r�p�h}�3��´  � �>��ph��`z��ꜞ�a��Jm�q� H�N��ac���dw���  �  �P� Q� �� |  а�m�Əi}	'� � ��I� �  �����:�È~�È=���(��ts�a	���I  ?�n @H�i~�ab�Ӌ�b�w���urN0��  '�Ж�q�p@2��@Ǔ���r�q5�C��pC0C�@ C�����`
��A1q) " � @B�V~X�
nwB0h�A��p�ӊa�p�`���aDz����֏���Я	�pv��( �� -��I��-�=��A&�a�we_q�`�p� �?�ff ���m��� �����Ƽuq@ݿ�>N1�  P�apv(�` ţ� �=�qst��/?���`x`�� �<
6b<߈�;܍�<�ê�<� <�&P�ό�AO��c1��ƾ��?fff?O�?y&��qt@�.���J<?�`�� wi4����dly�e߾g ;ߪ�t��p�[ߔ�� �ߣ����� ����6�wh�F0%�r�!�߷�1ى����E��� E�O�G+� F�!���/���?�e�P���t���lyBL�cB��Enw4��� ����+��R��s���������h�Ô�>��I�mXj�F��A�y�weC�p�������#/�*/c/N/wi�����fv/C�`� CHs/�`
=$�p�<!�!������'�3A�A��AR1AO�^?�$�?���5p±
=ç>�����3�W
�=�#�]�;e��׬a@����{�����<��>(�B�u���=B0��?����	R��z�H�F�G����G��H�U`�E���C�+���}I#�I���HD�F���E��RC�j�=�>
I���@H�!H�(� E<YD0 w/O*OONO9OrO]O �O�O�O�O�O�O�O_ �O8_#_\_G_�_�_}_ �_�_�_�_�_�_"oo oXoCo|ogo�o�o�o �o�o�o�o	B- fQ�u���� ���,��P�b�M� ��q�����Ώ���ݏ �(��L�7�p�[��� ���ʟ���ٟ����6�!�Z�E�W���#1(�$1��9�K���<ĥ%����Ư!3�8���!�4Mgs��,�I�B+8�J��a���{�d�d������ȿ���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ��ϰ�������  %��  ��h�Vߌ�z߰�&ڀg�/9�$������� 7����A�S�e�w�  ��������������2 F��$�&Gb��������!C���@����$����F�� DzN�� F?�P D�������)#B�'9K]�o#?���@@*v
��8�8��u8�.
 v ���!3EW i{����:�� ��ۨ�1���$MSKCFM�AP  ��� ����(.�ONREL  �!9��EXCFENBE'q
#7%^!FNCe/�W$JOGOVLI�ME'dO S"d�K�EYE'�%�R�UN�,�%�S?FSPDTY0g&<P%9#SIGNE/W$�T1MOT�/T!��_CE_GRP� 1p��#\ x��?p��?�?�?�? �?O�?OBO�?fOO [O�OSO�O�O�O�O�O _,_�OP__I_�_=_ �_�_�_�_�_oo�_�:o�TCOM_�CFG 1q	-оvo�o�o
Va_A�RC_b"�p)U?AP_CPL�ot$�NOCHECK {?	+ � x�%7I[m ���������!�.+NO_WAI�T_L 7%S2NT�^ar	+�s�_7ERR_12s	)9�� ,ȍޏ��x����&��dT_M�O��t��, 	i�*oq�9�PARAuM��u	+��`a�ß'g{�� =?��345678901��,��K�]�9� i�������ɯۯ��&g������C��cU�M_RSPACE�/�|����$OD�RDSP�c#6p(O�FFSET_CAsRT�o��DISƿ���PEN_FIL�E尨!�ai��`OPTION_IO�/���PWORK 5ve7s# ��V���8� "�ep�4�p��	 ���p��<����RG_DSBL'  ��P#������RIENTTOD ?�C�� !l����UT_SIM_ED$�"���V��?LCT w}���6��a[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ���� ��ڐH(���H3k7HS�M5G�22G�?��Gp
͜��'f�/-,ڐCR�>�D!�M#{Z/���3�����4y H "�c/u/�/�0B_����=jc��t�!�/ �/�"t32���~�/6  ��UP%�Q%��%�|T���S62�q?'e	'�� � �2I�� �  ��+==��ͳ?�;	��h	�0�I  �n @�2�.���Ov;��ٟ?&gN�]O  ''�uD@!:� C�C�@F#H!��/�O�O sb
�T��@�@��@$�e0@B�QA�0Y�v: �13Uwz $oV_�/z_e_�_�_	���( �� -�2�1�1ta�UDa�c���:A-���~.  �?�ff���[o"o�_U�`oXâ0A8���o�j>�1  Po�V(���eF0��f�Y���L�?˙���xb0@<
�6b<߈;����<�ê<�? <�&�,�/aA�;r�@Ov0P?offf?�0?&ipޘT@�.{r�J<?�`�u#	�B dqt�Yc�a�Mw �Bo��7�"�[�F� �j�������ُ� ���3����,���~(�E�� E��3?G+� F��a�� ҟ�����,��P�(;���B�pAZ�>� �B��6�<OίD���P� �t�=���a�s������6j�h��7o��>�S��O�����Fϑ�A�a�_���C3Ϙ�/�%?��?Ƀ��������#	���P �N||CH����Ŀ������@�I�_�'�3A��A�AR1A�O�^?�$�?������±
=�ç>����3�W
=�#� U���e���B��@���{����<����(�B��u��=B0�������	��b�H�F�G����G��H��U`E���C��+��I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻�������� � �9�$�]�H�Z��� ~�������������# 5 YD}h�� �����
C .gR����� ��	/�-//*/c/ N/�/r/�/�/�/�/�/ ?�/)??M?8?q?\? �?�?�?�?�?�?�?O �?7O"O[OmOXO�O|O �O�O�O�O�O�O�O3_:Q(������b���gUU��xW_i_2�3�8��_<�_2�4Mgs�_�_��RIB+�_�_�a?���{�mi�Go5okoYo�o}l��P'rP�nܡݯ�o=_`�o�_�[R?�Q�u���  �p���o��/�� S��z
uүܠ�������ڱ�����������  /�M�w��e��������l2 wF�$��Gb���t��a�`�p�S�C��y�@p�5�G�Y�۠F�� Dz��� F�P D��]����پ��ʯܯ�� ��~�?��ͫ@@�?�K��K���K���
 �|�������Ŀֿ �����0�B�T�f�ܽ�V� ���{���1��$PARA�M_MENU ?�3�� � DEF�PULSEr�	�WAITTMOU�T��RCV�� �SHELL_�WRK.$CUR�_STYL���	�OPT��PT�B4�.�C�R_DECSN���e��� �ߣ����������� !�3�\�W�i�{����USE_PROG %��%�����CCR���e�����_HOST !F��!��:���T�`�V��/�X����_TIME��^���  ��GDEB�UG\�˴�GINP_FLMSK�����Tfp����PGA�  ����)CH�����TYPE���������� � -?hcu �������/ /@/;/M/_/�/�/�/ �/�/�/�/�/??%?�7?`?��WORD �?	=	RS�fu	PNSU�Ԝ2JOK�DRT�Ey�]TRACE�CTL 1x3���� �`� &�`�`�>�6_DT Qy3�%@~�0D � �co�a:@V�@BR�2ODOVOhOzO�B�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofox`|d�b�h�o�g �m�a�o�o�o�ouJ� }�`M �b5GY~�`F��b�J�tr� ��O�ol���t� #�5��xZ�l�~�P���D\vR��d��N�qf 
��.�@�R�d�v��� ������П����� *�<�N�`�.Iv����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p��j��� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o��o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*���$PGTRACELEN  )��  ���(��>�_UP �z���m��u�Y�n�>�_C�FG {m�W�(�n���PК����DEFSPD �|��'�P���>�IN��TRL +}��(�8�����PE_CONFI���~m���mњ��ղ�LID����=�GRP� 1��W���)�A ���&f�f(�A+33D��� D]� C�O� A@1��Ѭ(��d�Ԭ��0�0�� 	 1�ح֚Ҏ�� ´�����B �9����O�9�s��(�>�T?�
�5�������� =?��=#�
�� ��P;t_�������  Dz (�
H� X~i����� �/�/D///h/S/��/��
V7.1�0beta1���  A�E>�"ӻ�A (�� �?!G��!>���"����!����!BQ��!A\�� �!���!2p����Ț/8?J?\?n?};!� ���/��/�? }/�?�?OO:O%O7O pO[O�OO�O�O�O�O �O_�O6_!_Z_E_~_ i_�_�_�_�_�_�_' o2o�_VoAoSo�owo �o�o�o�o�o�o.�R=v1�/�#F@ �y�}��{m� �y=��1�'�O�a� �?�?�?������ߏʏ ��'��K�6�H��� l�����ɟ���؟� #��G�2�k�V���z� �������o��ί C�.�g�R�d������� ���п	���-�?�*� cώ���Ϯ��� ���B�;�f�x��� ����DϹ��߶����� ���7�"�[�F�X�� |�����������!� 3��W�B�{�f����� ���� �����/ S>wbt��� ���=Oz� �Ͼψ����ϼ�  /.�'/R�d�v߈߁/ 0�/�/�/�/�/�/�/ #??G?2?k?V?h?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O ���O�O�O__?_*_ c_N_�_r_�_�_�_�_ �_o�_)oTfx� to���/�o/ >/P/b/t/mo� |������� 3��W�B�{�f�x��� ��Տ�������A� S�>�w�b����O��џ ������+��O�:� s�^�������ͯ��� ܯ�@oRodo�o`��o �o�o��ƿ�o���* <N�Y��}�hϡ� ���ϰ��������
� C�.�g�Rߋ�v߈��� ������	���-��Q� c�N�ﲟ���l��� �����;�&�_�J� ��n����������� ,�>�P�:L������ ������(�:� 3��0iT�x� ����/�/// S/>/w/b/�/�/�/�/ �/�/�/??=?(?a? s?��?�?X?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O* \&_8_r���_�_���$PLID_�KNOW_M  ���| Q�TSV ����P� �?o"o4o�OXoCoUo��o R�SM_GROP 1��Z'0{`��@�`uf�e�`
�5� �gpk 'Pe]o� ��������V�SMR�c��mT�EyQ}? yR������ ����폯���ӏ�G� !��-����������� 韫���ϟ�C��� )�����������寧����QST�a1 1Ն�)���P0� A 4��E2�D� V�h�������߿¿Կ ���9��.�o�R�dπvψ��ϬϾ����2r�0� Q�<3߂�3�/�A�S��4 l�~ߐߢ��5���������6
��.�@��7Y�k�}���8��������MAD  )���PARNUM  �!�}o+��SCHE� S�
��f���S��UPDf�x���_CMP_0�`H�� �'�U�ER_CHK-����ZE*<RS8r��_�Q_MOG���_�X�_RES_G��!���D� >1bU�y� ����/�	/����+/�k�H/ g/l/��Ї/�/�/� 	��/�/�/�X�?$? )?���D?c?h?�����?�?�?�V 1�x�U�ax�@c]�@}t@(@c\�@}�@D@c[�*@���THR_IN�Rr�J�b�Ud2FM�ASS?O ZSGM�N>OqCMON_QUEUE ��UX�V P~P X�N$ �UhN�FV�@ENqD�A��IEXE�O��E��BE�@�O�CO�PTIO�G��@P�ROGRAM %�J%�@�?���B?TASK_IG�6^OCFG ��Oxz��_�PDATA�c]��[@Ц2=� DoVohozo�j2o�o�o �o�o�o);M^ jINFO[��m��D����� ���1�C�U�g�y� ��������ӏ���	�4dwpt�l )�Q~E DIT ��_|i��^WERFLX�	C�RGADJ ��tZA�����?�נʕFA��IORI�TY�GW���MPGDSPNQ����U�GyD��OTOE@�1�X� (!�AF:@E� c�Ч�!tcpn����!ud����!�icm���?<�XYm_�Q�X���Q)� *�1�5��P��]�@�L���p� �������ʿ��+�@=�$�a�Hυϗ�*��OPORT)QH��P��E��_CAR�TREPPX��S�KSTA�H�
SS�AV�@�tZ	2500H863��P�_x�
�'��X�@�swPtS�ߕߧ�^��URGE�@B��6x	WF��DO�F"�[W\�������WR�UP_DELAY� �X���R_HOTqX	B%�c����R_NORMAL�q^R��v�SEMI������9�QSKI�P'��tUr�x 	7�1�1��X�j� |�?�tU���������� ����$J\n 4������� �4FX|j �������/ 0/B//R/x/f/�/�/��/tU�$RCVT�M$��D�� DC�R'���Ў!?��1�C�k�>��>5F=��� �0r�������A����i�:�o?2? �<
6b<���;܍�>u.��?!<�&�?h?�?�?�@>��? O O2ODOVOhOzO�O �O�O�O�O�?�O�O_ _@_+_=_v_Y_�_�_ �?�_�_�_oo*o<o No`oro�o�o�o�_�o �o�o�o�o8J- n��_����� ��"�4�F�X�j�U ������ď���ӏ� ��B�T��x����� ����ҟ�����,� >�)�b�M��������� ���ïկ�Y�:�L� ^�p���������ʿܿ � ����6�!�Z�E� ~ϐ�{ϴϗ�����-� � �2�D�V�h�zߌ� �߰���������
��� .��R�=�v��k�� ���������*�<� N�`�r���������� ������&J\ ?������� �"4FXj|���!GN_ATC� 1�	; �AT&FV0E�0�ATDP�/6/9/2/9��ATA�,�AT%G1%�B960�+�++�,�H/,��!IO_TYPE'  �%�#t��REFPOS1 �1�V+ x�u/�n�/j�/
= �/�/�/Q?<?u??�?�4?�?X?�?�?�+2 1�V+�/�?�?\O��?�O�?�!3 1� O*O<OvO�O�O_�OS4 1��O�O�O�_�_t_�_+_S5 1�B_T_f_�_o	o|Bo�_S6 1��_��_�_5o�o�o�oUoS7 1�lo~o�o�o�H3l�oS8 1�%_����SMASK 1�V/  
?�M��'XNOS/�r�������!MOTE  �n��$��_CFG �����q���"PL_RANG������POWER �����SM_D�RYPRG %�o�%�P��TAR�T ��^�UME_PRO-�?�����$_EXEC_E�NB  ���GSPD��Րݘ��gTDB��
�RM�.
�MT_'�T�����OBOT_N�AME o�����OB_ORD_NUM ?��b!H863  �կ�����PC_TI�MEOUT�� xޚS232Ă1��� LTE�ACH PENDcAN��w��-���Maint�enance CGons���s�"��~�KCL/Cm�Ț

���t�ҿ No Use-p��Ϝ�0�NPO�\򁋁��.�oCH_L�������q	��s�MAVGAIL�����糅���SPACE1 ;2��, j�߂ �D��s�߂� �{~S�8�?�k� v�k�Z߬��ߤ��ߚ � �2�D���hߊ�|� ��`��������� � �2�D��h��|� ��`���������y���2����0�B��� f�����{���3);M_ ������/� /44FXj |*/���/�/�/?(??=?5Q/c/u/ �/�/G?�/�/�?O�? $OEO,OZO6n?�? �?�?�?dO�?�?_,_@�OA_b_I_w_7�O �O�O�O�O�_�O_(o�Ioo^oofo�o8 �_�_�_�_�_�oo6o Ef){����G �o� t���
M� � ��*�<�N�`�r����� ��w���o�収���d.��%�S�e�w� ����������Ǐَ�� �Θ8�+�=�k�}��� ����ůׯ͟���� %�'�X�K�]������� ��ӿ������#��E�W� `� @�������x�����\�e���������� �R�d߂�8�j߬߾� �ߒߤ���������� 0�r���X�����������8����
��ύ�_MODE�  �{��S E��{|�2�0�����3�	S|)�CWORK_AD޳���+R  �{�`� �� _INTVAL����d���R_OPT�ION� ���H VAT_GRPw 2��upG(N�k |��_���� �/0/B/��h�u/T�  }/�/�/�/�/�/�/ ?!?�/E?W?i?{?�? �?5?�?�?�?�?�?O /OAOOeOwO�O�O�O �OUO�O�O__�O=_ O_a_s_5_�_�_�_�_ �_�_�_o'o9o�_Io oo�o�oUo�o�o�o�o �o�o5GYk- ���u���� �1�C��g�y���M� ����ӏ叧�	��-� ?�Q�c����������� ����ǟ�;�M��_����$SCAN�_TIM��_%�}�R �(�#�((�<04Wd d 
�!D�ʣ��u��/�����U�"�25���@�d5�P�g��]	����������dd�x�  P~���� ��  8� ҿ�!���D��$�M�_�q� �ϕϧϹ��������8ƿv��F��X��/� ;�o�b��pm��t�_DiQ̡  � l�|�̡ ĥ�������!�3�E� W�i�{�������� ������/�A�S�e� ]�Ӈ����������� ��);M_q ������� r���j�Tfx� ������// ,/>/P/b/t/�/�/�/p�/�/�%�/  0�� 6��!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O *�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo �O�OJ�o�o�o�o�o �o�o 2DVh z�������
�7?  ;�>�P� b�t���������Ǐُ ����!�3�E�W�i��{�������ß � ş3�ܟ��&�8�J��\�n�������������ɯ����,�� �+�	12�345678��W 	� =5���@f�x���������� ���
��.�@�R�d� vψϚ�៾������� ��*�<�N�`�r߄� �Ϩߺ��������� &�8�J�\�n�ߒ�� �����������"�4� F�u�j�|��������� ������0_�T fx������ �I>Pbt �������! /(/:/L/^/p/�/�/ �/�/�/�/�2�/�?�#/9?K?]?�i�Cz  Bp˚ /  ��h2��*��$SCR_GR�P 1�(�U8�(�\x�d�@ � ��'�	 ?�3�1 �2�4(1*�&�I3�Fp1OOXO}m��CD�@�0ʛ)���H�UK�LM-10�iA 890?�9�0;��F;�M61�C D�:�CP��1

\&V�1	�6F� �CW�9)A7Y	(R�_��_�_�_�_�\���0i^�oOUO>o Po#G�/���o'o�o��o�o�oB�0ƐrtAA�0* C @�Bu&Xw?���ju�bH0{UzAF?@ F�`�r� �o�����+�� O�:�s��mBqrr����������B�͏b�� ��7�"�[�F�X���|� ����ٟğ���N��� AO�0�B�CU
L���xE�jqBq>7�����$G@�@pϯ BȆ��G�I
E�0E�L_DEFAUL�T  �T���E��MI�POWERFL � 
E*��7�WF�DO� *��1E�RVENT 1����`(�� L�!DUM_EI�P��>��j!AF_INE�¿C�O!FT�����r�!o:� ���a�!RPC_M'AINb�DȺPϭ�Nt�VIS}�Cɻ�����!TP��PU��ϫ�d��E�!
P�MON_PROX	YF߮�e4ߑ��_��f����!RD�M_SRV�߫�g��)�!R�IﰴYh�u�!
v�M���id���!RL�SYNC��>�8|���!ROS��4��4��Y�(�}��� J�\����������� ��7��["4F� j|����!��Eio�ICE_�KL ?%� �(%SVCPRG1n>���3��3���4//�5./3/�6V/[/��7~/�/��D�/�9�/�+�@��/�� #?��K?��s?�  /�?�H/�?�p/�? ��/O��/;O��/ cO�?�O�9?�O� a?�O��?_��?+_ ��?S_�O{_�)O �_�QO�_�yO�_� �Os����>o�o }1�o�o�o�o�o�o�o ;M8q\� �������� 7�"�[�F��j����� ��ُď���!��E� 0�W�{�f�����ß�� �ҟ���A�,�e� P���t��������ί��y_DEV ���MC:����_!�OU�T��2��RE�C 1�`e�j�� � 	��  �������Fg �������̿��Ge��������
 �PSD#6 r�����O��������`D�����`e�����堆�0�  +T^�3���I3��3�!3����^Ͽ�_�^`ePSJ;:��U��?��(�ϋ �������RZ������E3�����
�k���Cl:̠��̒���
^��&�2�D�Vߜ�T�ߌ�":���=��*����؆����Y����-�����
��"3����b���*� �������(��L�:� p���d�����������  ��$ZH~ l�������  VDz�n ������/./ /R/@/b/�/v/�/�/�/}�2��/�/�/? :?(?^?L?�?�?v?�? �?�?�?�?�? O6OO FOlOZO�O~O�O�O�O �O�O_�O2_ _B_h_ V_�_n_�_�_�_�_�_ 
o�_.o@o"odoRoto vo�o�o�o�o�o�o <*`Np�x �������8� J�,�n�\��������� Ə�Ώ�����F�4��j�X���`�p�V 1�}� P����ɿ��$ 
�_ �y���TYPE\���HELL_CF�G �.�є��8��}��RS-Ѡ� ����֯������	� B�-�f�Q�c���������������ؐ�%�3�E��Q�)�a��M�o�p�����2��d]�K�:�H�K 1�H�  u�������A�<�N� `߉߄ߖߨ������߀����&�8��=�OMM �H���9��FTOV_ENB�&�1�OW_RE�G_UI��8�IM/WAIT��a���OUT������T�IM�����V�AL����_UNI�T��K�1�MON_�ALIAS ?e~w� ( he�� ����������ж�� );M��q��� �d��%� I[m�<�� ����!/3/E/W/ /{/�/�/�/�/n/�/ �/??/?�/S?e?w? �?�?F?�?�?�?�?�? O+O=OOOaOO�O�O �O�O�OxO�O__'_ 9_�O]_o_�_�_>_�_ �_�_�_�_�_#o5oGo Yokoo�o�o�o�o�o �o�o1C�og y��H���� 	��-�?�Q�c�u� � ������ϏᏌ��� )�;��L�q������� R�˟ݟ�����7� I�[�m��*�����ǯ ٯ믖��!�3�E�� i�{�������\�տ� ����ȿA�S�e�w� ��4ϭϿ����ώ��� �+�=�O���s߅ߗ� �߻�f�������'� ��K�]�o���>�� ��������#�5�G� Y��}���������n���$SMON_D�EFPRO ������� *SYS�TEM*  d=���RECALL� ?}�� ( ��}3copy �frs:orde�rfil.dat� virt:\t�mpback\=�>inspiro?n:3648��r؄�n�}*.mdb:*.*CU
Y����	.x.:\�8R�n��
�/.a6H_^ �//�-?Qb/ t/�/�/�F/��/�/ ??)�M�/p?�? �?�8?J?��? OO��%
xyzrate 61 �?�?�?�nO�O�O�%.GR(6044 HOZO�O�O _"/4/�/�Ga_s_�_ �_�/E_�HY_�_�_o !?3?FO�C�_no�o�o �?6oHo�@^o�o &_8_�_�_m��_ �_�_Z���"o4o �oXoi�{����o�oC� �o����0BT e�w�����I��� ����,���P�a�s� ������;�Ώ`��� �(�:�ßޯo����� ����ʟ\�����$� ��ɯZ�k�}ϏϢ��� E�د����� O2O�����g�yߋߞO�O:5076�OY������ !�3�����a�s��� ��E��Y������!� 3�F�����n������� 6�H���^���&� 8�����m���� ��Z��"�4��� X�i{�����C�� ��/�0���e/�w/�/�߮�� 4060��Y/�/�/?!3 ��(a?s?�?�?�E?��(Y?�?�?O!8�$�SNPX_ASG 1����9A�� P �0 '%R[1]@1.1O 9?�#3%dO�OsO �O�O�O�O�O�O __ D_'_9_z_]_�_�_�_ �_�_�_
o�_o@o#o doGoYo�o}o�o�o�o �o�o�o*4`C �gy����� ��	�J�-�T���c� ������ڏ����� 4��)�j�M�t����� ğ������ݟ�0�� T�7�I���m������� �ǯٯ���$�P�3� t�W�i��������ÿ ����:��D�p�S� ��wω��ϭ��� ��� $���Z�=�dߐ�s� �ߗߩ������� �� D�'�9�z�]���� �����
����@�#� d�G�Y���}������� ������*4`C �gy����� �	J-T�c ������/� 4//)/j/M/t/�/�/ �/�/�/�/�/?0?4�,DPARAM �9ECA ��	��:P�4�0�$HOFT_KB_?CFG  p3?E��4PIN_SIM  9K�6�?�?��?�0,@RVQST_P_DSB�>�2�1On8J0SR ���:� & C�AR=O~N�6T�OP_ON_ER�l@�F�8�APTN� �5�@�A�BRING_�PRM�O J0V�DT_GRP 1y�Y9�@  	�7 n8_(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 Dkhz���� ���
�1�.�@�R� d�v���������Џ�� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\������� ����ȯگ����"� I�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� tߛߘߪ߼������� ��(�:�a�^�p�� ���������� �'� $�6�H�Z�l�~��������������3VPRG_COUNT�6���A�5ENB��OM=�4J_U�PD 1��;8  
p2��� ��� )$6H ql~����� /�/ /I/D/V/h/ �/�/�/�/�/�/�/�/ !??.?@?i?d?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_�_�_Y?SDEBUG" � ��Pdk	�PSP_�PASS"B?~�[LOG ��+m�P�X�_�  �g�Q
M�C:\d�_b_M�PCm��o�o��Qa�o �vfSAV �m:dUb�U�\gSV�\TE�M_TIME 1]�� (�PճT�ԱXfoT1SV�GUNS} #'�k�spASK_OPTION" �g�ospBCCFGg ��| �b�{�}`����a &��#�\�G���k��� ��ȏ������"�� F�1�j�U���y���ğ ���ӟ���0��T�f��UR���S���Ư A������ ��D��n d��t9�l��������� ڿȿ�����"�X� F�|�jϠώ��ϲ��� ������B�0�f�T� v�xߊ��ߦؑ����� ��(��L�:�\�� p�����������  �6�$�F�H�Z���~� ������������2  VDzh��� ������4F dv����� �//*/�N/</r/ `/�/�/�/�/�/�/�/ ??8?&?\?J?l?�? �?�?�?�?�?�?�?O O"OXOFO|O2�O�O �O�O�OfO_�O_B_ 0_f_x_�_X_�_�_�_ �_�_�_oooPo>o tobo�o�o�o�o�o�o �o:(^Ln p�����O�� $�6�H��l�Z�|��� ��Ə؏ꏸ����2�  �V�D�f�h�z����� ԟ����
�,�R� @�v�d���������ί Я���<��T�f� ������&�̿��ܿ� �&�8�J��n�\ϒ� �϶Ϥ���������� 4�"�X�F�|�jߌ߲� ������������.� 0�B�x�f��R����� �������,��<�b� P�������x������� ��&(:p^ �������  6$ZH~l� �������/&/ D/V/h/��/z/�/�/�/�/�&0�$TB�CSG_GRP �2��%��  �1 
 ?�  /?A?+? e?O?�?s?�?�?�?�?��;23�<d�, �$A?1	 �HC���6>���@E�5CL  B�'2^OjH4J��B\)LFY  3A�jO�MB��?�I#Bl�O�O�@�JG_>�@�  D	�15_ __$YC-P{_F_`_j\��_�]@0�>�X �Uo�_�_6oSoo0o�~o�o�k�h�0	�V3.00'2	�m61c�c	�*�`�d2�o�e>�dJC0(�a�i ,p��m-  �0�����omvu1JCFoG ��% 1Y #0vz��rBr�|�|����z � �%��I�4�m�X� ��|��������֏� ��3��W�B�g���x� ����՟������� �S�>�w�b�����'2 A ��ʯܯ������ E�0�i�T���x���ÿ տ翢����/��?� e�1�/���/�ϜϮ� �������,��P�>� `߆�tߪߘ��߼��� �����L�:�p�^� ������������  �6�H�>/`�r���� ������������  0Vhz8��� ���
.�R @vd����� ��//</*/L/r/ `/�/�/�/�/�/�/�/ �/?8?&?\?J?�?n? �?�?�?�?���?OO �?FO4OVOXOjO�O�O �O�O�O�O__�OB_ 0_f_T_v_�_�_�_z_ �_�_�_oo>o,obo Poroto�o�o�o�o�o �o(8^L� p������� $��H�6�l�~�(O�� ��f�d��؏���2�  �B�D�V�������n� ���ԟ
���.�@�R� d����v�������� Я���*��N�<�^� `�r�����̿���޿ ��$�J�8�n�\ϒ� �϶Ϥ�������ߊ� (�:�L���|�jߌ߲� �����������0�B� T��x�f������ �������,��P�>� t�b������������� ��:(JL^ ������ � 6$ZH~l� �^���dߚ // D/2/h/V/x/�/�/�/ �/�/�/�/?
?@?.? d?v?�?�?T?�?�?�? �?�?OO<O*O`ONO �OrO�O�O�O�O�O_ �O&__6_8_J_�_n_ �_�_�_�_�_�_�_"o oFo��po�o,oZo �o�o�o�o�o0 Tfx�H��� ����,�>��b� P���t���������Ώ ��(��L�:�p�^� ������ʟ���ܟ�  �"�$�6�l�Z���~� ����دꯔo��&� ЯV�D�z�h������� Կ¿��
��.��R��@�v�dϚτ�  ���� ��������$TBJOP_�GRP 2ǌ���  �?�������������x�JBЌ��9� �< �X�ƞ�� @���	� �C�� t�b�  C����>ǌ�͘Րդ�>���йѳ33=��CLj�fff?>��?�ffBG���Ќ�����t�ц�>;�(�\)�ߖ��E噙�;��h{CYj��  @h�~�B�  A�����f��C�  D�hъ�1��O��4�N����
:�/��Bl^��j�i��l�l����Aə�3A�"��D���Ǌ=qH���нp��h�Q�;��A�j�ٙ�@L��D	2�������<$�6�>B�\��T����Q�tsx�@g33@���C����y�1����>��Dh����������O<{�h�@i�  ��t��	� ��K&�j� n|���p�/��/:/k/�ԇ����!��	V3.0}0J�m61cIԃ*� IԿ��/�'� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�I�!CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;��;Q�UT,8�4` *���?�2���3\�X/�O��ESTPAR�S  ��	���H�R@ABLE 1%����0��
H�7Q 8��9
G
H
H�����
G	
H

H�
HYE��
H
H:
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_t_�^:BS _� �JGoYo ko}o�o�o�o�o�o�o �o1CUgy ����`#oRL�y�_ �_�_�_�O�O�O�O�O�X:B�rNUM  ����P���� V@P:B_CF�G ˭�Z�h�@���IMEBF_T�T%AU��2@�VE�RS�q��R {1���
 (�/����b� ����J� \���j�|���ǟ��ȟ ֟�����0�B�T�@��x�������2�_����@�
��MI_�CHAN�� � >��DBGLV����������ETHE�RAD ?��
O�������h������ROUT�!���!������SN�MASKD��U�255.���#������OOLOFS_�DI%@�u.�OR�QCTRL � ����}ϛ3rϧϹ��� ������%�7�I�[��:���h�z߯�APE?_DETAI"�G��PON_SVOF�F=���P_MON� �֍�2��S�TRTCHK ��^�����VTCOMPAT��O������FPROG =%^�%CA����~��ISPLAY&H���_INST_M�ް ������US8�q��LCK���QUICKME��=���SCREZ�}G�tps� @���u�z����_���@@n�.�SR_GR�P 1�^� �O����
��@+O=sa�� ��
m������ L/C1gU� y�����	/��-//Q/?/a/�/	1234567�0h�/�/@Xt�1����
 �}ipn�l/� gen.htm�? ?2?D?V?�`Panel� setupZ<}�P�?�?�?�?�?�? �??,O>OPObOtO �O�?�O!O�O�O�O_ _(_�O�O^_p_�_�_ �_�_/_]_S_ oo$o 6oHoZo�_~o�_�o�o �o�o�o�oso�o2D Vhz�1'� ��
��.��R�� v���������ЏG����UALRM��G ?9� �1�#� 5�f�Y���}������� џן���,��P���SEV  �����ECFG C��롽�A���   BȽ�
 Q���^����	�� -�?�Q�c�u�������4������ ������I��?���(%D�6� �$�]�Hρ� lϥϐ��ϴ�������`#��G���� ��߿U�I_Y�HIS�T 1��  �(� ��(�/SOFTPAR�T/GENLIN�K?curren�t=editpa7ge,��,1����(�:�'����m7enu��71�߅� ����J�=������ �+�=���a�s����� ����J�����' 9����o���� �X��#5G �k}������f��f//'/9/ K/]/`�/�/�/�/�/ �/j/�/?#?5?G?Y? �/�/�?�?�?�?�?�? x?OO1OCOUOgO�? �O�O�O�O�O�OtO�O _-_?_Q_c_u__�_ �_�_�_�_�_��)o ;oMo_oqo�o�_�o�o �o�o�o�o%7I [m� ��� ����3�E�W�i� {������ÏՏ��� ����A�S�e�w��� ��*���џ����� ooO�a�s������� ��ͯ߯���'��� K�]�o���������F� ۿ����#�5�ĿY� k�}Ϗϡϳ�B����� ����1�C���g�y� �ߝ߯���P�����	� �-�?�*�<�u��� �����������)� ;�M������������ ����l�%7I [������� hz!3EWi �������v�////A/S/e/P����$UI_PAN�EDATA 1������!  	�}w/��/�/�/�/?? ) ?>?V�/i?{?�?�? �?�?*?�?�?OOO AO(OeOLO�O�O�O�O��O�O�O�O_&Y� b�>RQ?V_h_z_ �_�_�__�_G?�_
o o.o@oRodo�_�ooo �o�o�o�o�o�o* <#`G��}�-\�v�#�_��!� 3�E�W��{��_���� ÏՏ���`��/�� S�:�w���p�����џ ������+��O�a� ��������ͯ߯� D����9�K�]�o��� �����ɿ���Կ� #�
�G�.�k�}�dϡ� �����Ͼ���n���1� C�U�g�yߋ��ϯ��� 4�����	��-�?�� c�J�������� �������;�M�4�q� X����������� %7��[��� ����@�� 3WiP�t� ����/�//A/ ����w/�/�/�/�/�/ $/�/h?+?=?O?a? s?�?�/�?�?�?�?�? O�?'OOKO]ODO�O hO�O�O�O�ON/`/_ #_5_G_Y_k_�O�_�_ ?�_�_�_�_oo�_ Co*ogoyo`o�o�o�o �o�o�o�o-Q08u�O�O}��� �����)�>� �U-�j�|�������ď +��Ϗ���B�)� f�M���������������ݟ��XS�K�$�UI_PANEL�INK 1�U�  ��  ��}12�34567890 s���������ͯդ�R q����!�3�E�W�� {�������ÿտm�m��&����Qo�   �0�B�T�f�x��v� &ϲ���������ߤ� 0�B�T�f�xߊ�"ߘ� ���������߲�>� P�b�t���0���� ��������$�L�^� p�����,�>�������0 $�0,&�[ �XI�m���� ���>P3t �i��Ϻ� - n��'/9/K/]/o/�/ t�/�/�/�/�/�/? �/)?;?M?_?q?�?� UQ�=�2"��?�?�? OO%O7O��OOaOsO �O�O�O�OJO�O�O_ _'_9_�O]_o_�_�_ �_�_F_�_�_�_o#o 5oGo�_ko}o�o�o�o �oTo�o�o1C �ogy����� B�	��-��Q�c� F�����|������� ֏�)��M���=�? ��?/ȟڟ���� "�?F�X�j�|����� /�į֯�����0� �?�?�?x��������� ҿY����,�>�P� b��ϘϪϼ����� o���(�:�L�^��� �ߔߦ߸�������}� �$�6�H�Z�l��ߐ� ���������y�� � 2�D�V�h�z����-� ��������
��. RdG��}�� ��c���<��` r�������� //&/8/J/�n/�/ �/�/�/�/7�I�[�	� "?4?F?X?j?|?��? �?�?�?�?�?�?O0O BOTOfOxO�OO�O�O �O�O�O_�O,_>_P_ b_t_�__�_�_�_�_ �_oo�_:oLo^opo �o�o#o�o�o�o�o  ��6H�l~a �������� 2��V�h�K����� ��1�U
��.�@� R�d�W/��������П ������*�<�N�`� r��/�/?��̯ޯ� ��&���J�\�n��� ����3�ȿڿ���� "ϱ�F�X�j�|ώϠ� ��A���������0� ��T�f�xߊߜ߮�=� ��������,�>��� b�t�����+�� ����:�L�/�p� ��e�����������  ��6���ۏ���$UI_QUI�CKMEN  >���}���RESTORE� 1٩�?  �
�8m3\n� ��G����/ �4/F/X/j/|/'�/ �/�//�/�/??0? �/T?f?x?�?�?�?Q? �?�?�?OO�/'O9O KO�?�O�O�O�O�OqO �O__(_:_�O^_p_ �_�_�_QO[_�_�_I_ �_$o6oHoZoloo�o �o�o�o�o{o�o  2D�_Qcu�o� ������.�@� R�d�v��������Џ�⏜SCRE� ?��u1s]c� u2�3�U4�5�6�7�y8��USER��d��T���ks'����4��5��6��7�8��� NDO_�CFG ڱ � �  � PDA�TE h���None�SE�UFRAME  �ϖ��RTO?L_ABRT�����ENB(��GR�P 1��	�Cz  A�~�|�%@|�������į֦ை�X�� UH�X�7�MSK  K�S�7�MN�%uT�%������VISCAN�D_MAXI�I��3���FAIL_�IMGI�z �% #�S���IMREGN�UMI�
���SI�ZI�� �ϔ,~�ONTMOU'��K�Ε�&�����(��(��~s�FR:\��� � MC{:\(�\LOGh�7B@Ԕ !{���������z �MCV����U�D1 �EX	�|z ��PO64_úQ��n6��PO!�LI�Oڞ�e�9V�N�f@`�I��� =	_�SZV�mޘ��`�WAI�mߠ�STAT 	�k�% @��4�F�T��$#�x �2DW�P  ��P yG��=��͎����_JMPE�RR 1ޱ
 � �p2345678901���	� :�-�?�]�c������������������$�M�LOW�ޘ�����_�TI/�˘'��M�PHASE  �k�ԓ� ��SHI[FT%�1 Ǚ��<z��_�� ��F/|S e������� 0///?/x/O/a/�/@�/�/�/�/����k�	VSFT1[��	V��M+3 ��5�Ք p����A_�  B8[0[0E�Πpg3a1Y2�_3�Y�7ME��K�͗�	6e���&%��Mҿ��b��	��$���TDINEND3�4��4OH�+�G1��OS2OIV I��=�]LRELEvI���4.�@��1_ACT�IV�IT��B��A ��m��/_��BR�DBГOZ�YBOX� �ǝf_[���b�2�TI1�90.0.�P83vp\�V254p^:�Ԓ	 �S�_��[b��ro�bot84q_  � p�9o[�pc�PZoMh�]Hm��_Jk@1�o�ZABCd��k�,���P[� Xo}�o0);M �q���������>��aZ�b�� _V