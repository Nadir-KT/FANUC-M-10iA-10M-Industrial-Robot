��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|(�ARG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"GSB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�:�OFF_ N�3D;ELHLOGn25Aa2?i1@N�?�� -M��W�+0�$Y $DB\� 6COMW!2�MO� 21H _A.�	 \rVE�1�$F��A{$O��D�B�CTMP1k_F�E2�G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYPuAHK�BD_S�B�1AG�N Gn $SLOT_NUM�JQPREV,DBU�� g1G ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�AETE�_OKRUS�P7_CRQ$;4�V�� 0LACIw�1�RAPk �1x@ME>@$D�V�Q��Pv�A{�BLv� OUzR ,mAЧ0�!� B� LM�_O�^eR�"CAsM_;1 xr~$ATTR4�NP� ANN�@5I�MG_HEIGH|Q�cWIDTH4�VT� �UU0F_�ASPECQ$�M�0EXP��@A�X�f�CFT ?X $GR� � �S�!�@B@NFL�I�`t� UIREx 3dTuGITCHCj�`N� S�d_L�`2�C�"�`EDlpE
� J�4S�0� �zsa�!ip;G0 �� 
$WARNM��0f�!,P� �s�pN{ST� CORN�"�a1FLTR�uTRkAT� T�p H0ACCa1���{��ORI
`"S={R�T0_S�B�CHuG,I1 [ �Tp�"3I9�TYP�D,P*2 �`w@�� �!R*HD�cJ�* C��2��3��4���5��6��7��8���94�ACO�$ <� $6xK3 1�w`O_M�@�C �t � E#6NGP�ABA� �c��@ZQ���`���@nrH��� ��P�0��E^��w�p�PzPb2�6����"J�_R��BC�J��3�JVP��tBS��}Aw؅�"\�P_*0OF�SzR @� RO1_K8���aIT�3��ONOM_�0�1ĥ�3��pPT Ԑ� $���AxP��K}EX�� �0g0I01��p��
$TFa��C$7MD3��TO�3�0yU� �� �)Hw2�C1|�EΡg0wE{vF�vF�40�CPp@�a2 
P�$A`PU�3Nc)#�dR*�AX�!�sDETAI�3BU�FV�p@1 |X�p۶�pPIdT� +PP[�MZ�Mg�Ͱ�j�F[�SIMQS I�"0��A.�����Nlw Tp|zM�x�P�B�FACTrbHPEW7�P1Ӡ��v��MCd� �$*1JB�p<�*1DECHښ�H��a�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF4��� &k�Bv�u�cu��a E�� !2��+�MQ��EчSIZ�3����T��P�����aRSINF�����kq��������LX������F�CRCMu�3CC lpG��p���O}���b��1�������2�V�D
xIC��C���r����0P��{� EV �zUF_��F�pNB
0�?������A�! �r�Rx���� V�lp�2��aR�t�,��g�RTx �#�5�5"2��uARt���`CX�$LG�p��B�1 `s�P�t�a!A�0{�У+0R���tME�`!BupCr3RA 3tAZ�л4�pc�OT�FC�b�`��`FNp���1��ADI+�a%��b��{��p$�pSp�c�`S0�P��a,QMP6�`IY�3��M'�pU���aU  $>�TITO1�S�S�!���$�"0�DBPXW�O��!��$S9K��2SPC� ��"�"@�PR8� 
G�D���g# >�q1$��S$��+�L9$?H(�V�%@?R4C9&_?R4ENE���'~?�AI�!RE|�pY2(H ��OS��#$L�3$�$3R��;3�MVO�k_D@!V�ROS�crr�w�S���CRIoGGER2FPA�S|��7�ETURN0Bn�cMR_��TUܐ�[��0EWM%�ơ�GN>`��RLAȜ��Eݡ�P�&$P�t�'�@����C�DϣV�DXQ��4��1��MVGO_AWAYRMO#�aw!�DCS_o)  `IS# � �� �s3S�AQ�� 4Rx�ZSW�AQ�p��@1UW��cTNTV)�5RV
a���|c���Wƃ��JB��x0���SAFEۥ�V_S}V�bEXCLUU�:;��ONL��c1Yg�~az�OT�a{�HI_V? ��R, M�_ *�0� ��9_z�2� �Q;SGO  +�rƐ m@�A�c~b���w@���V�i�b�fANNU�Nx0�$�dIDY�UABc�@Sp�i�a+ D�j�f	_�ΰAPIx2,��$F�b�$ѐ�OT�@A $DUMMY��Ft���Ft±D`6U- 7` !�HE�|s��~bc�B@ SUF�FI��4PCA*�Gs5Cw6Cq�DMSWU. 8�!�KEYI��5�T�M�1�s�qoA�vIN�ޱ�D, / D���HOST�P! 4���<���<�°<��p�<�EM'���Z�D`S�BL� UL��0  �	��E�D`�T�01 � �$��9USAMPL�о�/���決�$ I�@갯 $SUB ӄ��w0QS�����#��SAV�����c�S�< 9�`�fP$�0E�!� YN_B�#2� 0�`DI�d�pO�|�m��#$F�R_�IC� �ENC�2_Sd3  ��< 3�9���� cgp����4�"��2�rA��ޖ5�� �`ǻ�@Q@K&D-!<�a�AVER�q�����DSP
���PC_�q��"�|�ܣ�oVALU3�HE��(�M�IP)���OkPPm �THЈ*��S" T�/�F�b�;�d����d �xp�16 H(rLL_DUǀ�a�@`��k���֠OT�"�U�/���@@NOA�UTO70�$�}�x�~�@s��|�C�����C� 2�w�L�� 8H *��L� ���Բ @sv��`� �� ÿ��� Xq��cq���q���q��U7��8��9��0����1�1 �1-�1�:�1G�1T�1a�1Jn�2|�2��2 �U2-�2:�2G�2T�U2a�2n�3|�3ʩ3� �3-�3:�3�G�3T�3a�3n�4�|������9 < ���z�ΓKI����H硵BaFEq@{@�: ,��&a? P_P?��>���E��E�@�ᶰ�QQ���;fp$TP~�$VARI��ܮ�,�UP2Q`< W�߃TD��g���`�������_BAC��"= T2����$)�,+r³�p IFI@��p�� q M�P"��l@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� Fa@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(��a�#5T�DG���� �%��FSS� )�? �P(q1�1�`_(1"811�EC1�3D;5D6�GRA����@�����PW��ON2EBU�G�S�2�C`gϐ_?E A �@a �TERM�5�B�5$Z �OR�Iw�0C�5����SM_-`���0D��9TA�9E�9UP>��F� -Qϒ�A�P�3�@B$S�EGGJ� EL�UU�SEPNFI���pBx��1@��4>DC$sUF�P��$����Q�@C���G�0T������SNSTj�P�ATۡg��APTH	J�A�E*�Z%qB\`@F�{E��F�q�pARxP<Y�aSHFT͢qA|�AX_SHOR$��>��6 @$GqPE���OVR���aZP�I@P@$U?r *aAGYLO���j�I�"���Aؠ��ؠERV ��Qi�[Y)��G�@R���i�e��i�R�!P�uASYM���uqA#WJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P���WkOR�@M��k0�SMT��G��GR��3�aPA�@���p|5�'�H � j��A�TOCjA7pP<]Pp$OPd�O�P�C�%�p�O!���RE.pR�C�AOX�?��Be5pR�E�ruIx'QG�e$PW�R) IMdu�RR_�$s �5��B �Iz2H8�=�_AD�DRH�H_LENAG�B�q�q:�x�R��So�J.�SS��SK������ ��-�cSE*����HSN�[MN1K	�j�05�@r�֣OL��\��WpW�Q�>pACRO �p���@H ����Q�� ��OUPW3�b_">�I��!q�a1���� ����|���������-���:���iIO
X2S=�D�e���p<`���L $��p��!_OFF[r_�P�RM_���HT�TP_�H��M (�pOBJ�"�pG�[$H�LE�C��>ٰN � 9�*��AB_�T��
�S��`�S��LV��KR�W"duHITCOU�?BGi�LO�q ����d� Fpk�GpsSS� ���HWh��wA��O.��`IN�CPUX2VISIO��!��¢.�á<��á-� �IOLN.)�P 87�R'�[p�$SL�bd P7UT_��$dp��Pz �� F_AuS2Q/�$LD���D�aQT U�0]P�Aa������PHYG�܁�Z� �
4�UO� 3R `F���H�@Yq�Yx�ɱvpP�S�dp���x��ٶ��UeJ��S����NE�W�JOG�G �DIS���r�KĠ��3T �|��AV��`_�CTyR!S^�FLAGf2vr�LG�dU �n��:��3LG_SIZ��ň��=���FD��I����Z �� ���0�Ʋ�@s��-ֈ� -�=�-���-��0-�I�SCH_��Dq��NT?���V��EE!2�C��n�U�����`�L�Ӕ�DAU��E�A��Ġt����GH�r��OGBOO>)�WL ?`�� �ITV���0\�REC�SCRf 0�a��D^�����MARG ��`!P�)�T�/ty�?I�S�H�WW�I����T�JGM��MNC�H��I�FNKEY���K��PRG��UqF��P��FWD��HL�STP��V`��@�����RSS�H�` �Q�C�T1�ZbT�R ���U����� |R��t�i���G��8PCPO��6�F�1�M���FOCU��RGE]XP�TUI��I���c��n��n�� ��ePf���!p6�eP7�9N���CANAI�jB޾�VAIL��CL�t!;eDCS_HI�4�.��O�|!��S Sn��0I�BUFF1XjY��PT�$��@ �v��fĵ�1�A�rYY��P �����pWOS1�2�3����0Z � � ��aiE�*��ID%X�dP�RhrO�+��A&ST��R��Y�z�<! Y$E�K&CK+���Z&m&8�5�0[ L��o� 0��]PL�6pwq�t^�𩐸t�7�_ \ ����瀰�7��#��0C��] ��C�LDP��;eTRQ�LI�jd.�094F�LGz�0r1R3�DM�R7��LDR5<4R5ORG.���e2(`�ŀ�V�8.��T<�4�d^� �q�<4��-4R5SB�`T00m��0DFRCLMC!D�?�?�3I@��pMIC��d_� d���RQm��q�DSTB	�  ��Fg�HAX;b ��H�LEXCESHZr��rBMup�a`�A�B;d�F`��`a��F_A�J��$[�Ot�H0K�db \���ӂS�$MB��LI�Б}SREQUIR��R>q�\Á�XDEB}U��DI�ML� MP�c�ba��P؃ӂ!B�AND���`�`ad�҆�c�cDC1��IN�����`@�(hB?Nz�@q��o��UwPST8� e�r7LOC�RI�p�EX�fA�p��A�A�ODAQP�f Xf��ON��[rMF�� ���f)�"I��%�e���T� �FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y�[�Eѭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?
�uD�)�b�	@Ð�i �@CU��V��T0�eRR2�j� Dɐ�Qނ�Bd$OCALI�@F�G�:s�2�RIN��v�=<�INTE����kE���,��b����_Nl��ڂ��o���tځRm�DIV�DH�@ـn�c$V��'c!$��$Z�����~��p@R�oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS�@#2L�q�Ɣ83ಀ����� ��PAT!H��������3̒Vp�A_�Q�.�4�B��Cᐈ�_MGh��$DDQ���G�$FWh��p��m������b�DE��PPAB�NԗROTSPE!ED����00J�Я�8��@���$US�E_��P��s�S�Y��c�A >qYNru@Ag��OFF�qn�MOUN�NGg��K�OL�H�INC *��a��q��Bj�L@�BENCS��q�BđX���D��IN#"I̒0��4�\BݠVEO�w�>Ͳ23_UPE�߳/LOWL���00����D���BwP���� �1RCʀƶMO3SIV�JRMO���@�GPERCH  �OV��^��i� <!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸUPp������TRKr�>"AYLOA'a��  Q-�̒<�1Ӣ`0 ���RTI$Qx�0 MO ���МB R�0J��D���s�H����b�DU�M2(�S_BCKLSH_C̒��>� =�q�#�U��ԑ���2�<t�]ACLALvŲp�1n�P�CHK00:'%SD�RTY4�k���y�1�q_6#2�_�UM$Pj�Cw�_�S�CL��ƠLMT_OJ1_LO��@���q��E�����๕�幘SPC��7���L���PCo���H� ȰPU�m�C/@�"XT\_�c�CN_��N��Le���SFu���V��&#����9�̒��=�C�u�SH6#��c��� �1�Ѩ�o�0�͑
��f_�PAt�h�_Ps�W�_10��4�R�01D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�sR0Hљ��_W��-ԁ_=��C��I��I*�I�II�F�`�aJLA.�1[�VC��0�D�BO1U�@i�B\JRKU��~	@DBL_SMd�:BM%`_DLC�BGRV��C��I���H_� �*CcOS+\�(LN� 7+X>$C�9)I�9)u*c,)�Z2 HƺcMY@!�( "TH&-��)THET0�N�K23I��"=�A C-B6CB=�C�A�B�(261C�616SB8C�T25GTS QơC��aS$" �4c#<�7r#$DUD�EX��1s�t��B�6���AQ�|r�f$NE�DpI B U�\B5��$!��!�A�%E(G%(!LCPH$U�2׵�2SX pCc%pCr%�2�&�C�J�&!�VAHV6H3�YLUVhJVuKV�KV�KUV�KV�KV�IHAH@ZF`RXM��wXuKH�KUH�KH�KH�KH�I�O2LOAHO�YWNO�hJOuKO�KO�KO*�KO�KO�&F�2#1�ic%�d4GSPBA?LANCE_�!�c�LEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%�Ċ1ky�UTO_<?�jT1T2Cy��2N&�v�ϰctw�gѠp�0Ӓ~���T��O����� INSEGv�!�REV�v!���gDIF��1l�w6�1m�0OB�q
����MIϰ1��L�CHWAR����A�B&u�$MEC�H,1� :�@�U�AX�:�P��Y�G$�8pn� 
Z��|���RO�BR�CR��N���'`�SK_�`f�p� P Np_��R ����΄ݡ�1��Ұ�Т΀ϳ��΀"�IN��q�MTCOM�_C@j�q  �L��p��$NO�RE³5���$�7r 8� GR�E��SD�0ABF�$?XYZ_DA5A���DEBU�qI���Q�s �`$�COD�� ��k�F��f�$BUFIwNDXР  ���MOR��t $-�U��)��r�B���������Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��E����͐OPWOܭŀv0��SY�SBU�@ʐ$SO!P����#�U"��p�PRUN�I�PA��DH�D����_O�U�=��qn�$^}�IMAG��ˀ��0P�qIM����I�N�q���RGOVCRDȡ:���|�P~���Р�0L_6p���Li��RB���0��M���EDѐF� J��N`M*���ⷀ�˱SL�`ŀw x $OVSL�vwSDI��DEXm�@g�e�9w�����V� ~�N���w����Û�d�ȳ�M�̐ ��q|<��� x Hˁ�E�F�ATUS����C�0àǒ��BT�M����If���4p����(�ŀy Dˀ!Ez�g���PE�r��p���
���EXE���V��E�Y�$Ժ ŀz3 @ˁ��UP{�h�3$�p��XN����9�H� �PG�"�{ h $S#UB��c�@_��01�\�MPWAI��PL����LO��<�F�p��$RCVFA�IL_C�f�BW�D"�F���DEFS}Pup | Lˀ�`�D�� U�UN!I��S���R`��V�_L�pP����P�ā}��� B��~���|��`ҲN�`KSET��y���P� �$�~���0SIZAE�ଠ{���S<��OR��FORMA�T/p � F���rEeMR��y�UX����@�PLI7�ā�  $�P_�SWI��Ş_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W �U����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�!O�0\H��6@�Q� ��ŀ�P�qUR_�SCR�ӚAZ��S_SAVE_D�,�E��NO��CgA�� ���@�$����I��	 �I� %Z[� ��RX " ��m���"�q�' "�8�Hӱt�W��UpS��рM�� O㵐.'}q��Cg�� �@ʣ���тM�AÂ�� � $PY���$WH`'�NGp���H`��Fb��Fb��Fb��PLM���	�P 0h�H�{�X��O���z�Z�eT�M���� pS��C��O_�_0_B_�a��_%�� |S����@	�v��v �@���w�v��EM��% �fr�B��ː��ftP���PM��QU� ŉU�Q��Af�QT�H=�HOL��QH�YS�ES�,�U�E��B��O#��  -�P0�|�gAQ����ʠu���O��ŀ��ɂv�-�A;ӝROG��a2D�E�Â�v�_�ĀZ�INFOB&��+����bȁ�OI킍 ((@SLEQ/�#�������o���S`c0O��0�01EZ0N9Ue�_�AUT�Ab�COPY��Ѓ�{�
�@M��N�����1�4P�
� ��RGI��͏��X_�Pl�$P�����`�W��P���j@�G���EXT/_CYCtb���p����h�_NAƹ!$�\�<�RO��`]�� � m��POR�ㅣ�.��SRVt�)����DI �T_l���Ѥ@{�ۧ��ۧ �ۧ5٩�6٩7٩8��R�S��B쐒��$�F6���PL�A�A^�TAR��@E `�Z�����<��d� ,�(@FLq`h��@YN�L���M�C���P�WRЍ�쐔e�D�ELAѰ�Y�pA�D#q�RQSKIPN�� ĕ�x�O�`�NT!���P_ x���ǚ@�b�p1� 1�1Ǹ�?� �?���>��>�&�>�3�>�9��J2R;쐖� 4��EX� TQ ����ށ�Q���[�K�Fд���RDCIf�S �U`�X}�R��#%M!*�0�)��$RGoEAR_0IO�T�JBFLG�igpE	Ra��TC݃�����ӟ2TH2N��� �1�b��Gq TN�0 ����M����`Ib���QREF:�1�� l�h���ENAB��lcTPE?@���!(ᭀ�� ��Q�#�~�+2 H�W S��2�Қ�߀�"�4�F�X�W���3�қ{��������
��4�Ҝ��
��.�(@�R���5�ҝu��������������6�Ҟ���(:L��7�ҟo�����
��8�Ҡ��"x4F��SMSK������a��E�A�����MOTE������@ "1��Q�IO�5"%I��P��POWi@쐣 8 �����NA��h��쐤��Y"$DSB_SIGN4A�Qi��̰C��>%S232�%�Sb�iDEVI�CEUS#�R�RP�ARIT�!OP�BIT�Q��OWCONTR��Qⱬ��RCU� M�SU_XTASK�3NB���0�$TATU�P%��S@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�UKPDl�ARB73P%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG �G|�.2���F��1�!d�9Z�8+5K��+5��E�y�L0�4��X �0m�LN�T�3Hz��89��%�4�3%G��W�0�W�RdD�Z��Tܳ��K�a�3d��$cV 2!���1��I1H�0U2K2sk3K3J ci�aI�i�a�L��SLL��R$Vؠ�BV�E�Vk�]V*R��� � ,6Lc���9V2F{/P�:B��PS_�E���$rr�C�ѳ$A0��wPR���v�U�c�Sk�� {��8��� 0���VX`�!�tX`A��0P�Ё�
�5�SK!� �-qRH��!0���z�NJ SAX�!h�A�@LlA���A�THIC�1p�������1TFE��|�q>�IF_CH�3�A�I0�����G1@�x������9�Ɇ7_JF҇PR(����RVAT��� �-p��7@����D9O�E��COU(���AXIg��OFF{SE+�TRIG�S K��c���Ѽ�e�[�K��Hk���8�IGMA�o0�A-��ҙ�OR?G_UNEV���� �S�쐮d� �$������GgROU��ݓTO2���!ݓDSP��JO1G'��#	�_P'�2�OR���>P6KE�Pl�IR�0�PML�RQ�AP�Q��E�08q�e���SYSG��"v��PG��BRK*Rd�r�3�-��������ߒ<pAD��ݓJ�B�SOC� N�D?UMMY14�p\@�SV�PDE_OP�3SFSPD_O+VR��ٰCO��&"�OR-��N�0.��Fr�.��OV�S!Fc�2�f��F��!�4�S��RA�"LCH�DL�RECOV(��0�W�@M�յF�RO3��_��0� @�ҹ@VE}RE�$OFS�@3CV� 0BWDG�Ѵ`C��2j�
�TR�!���E_FDO>j�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�<#�8$CA�{�|����8$HBK|1,c��IO��.�:!aPPA"�N�3�^��F���:"�DVC_DB�C��d�w"���D�!��1���ç�3��^��ATIO� �q�0�UC�&CAB�BS�PⳍP��䖁�_0c�SUB'CPUv"�S�Pa  aá�}0�Sb��c��V"~ơ$HW_C�����:c��IcA�A-�l_$UNIT��l���ATN�f����CY{CLųNECA���[�FLTR_2_�FI���(��}&��L�P&�����_SCT@SF_��F����G����FS|!�¹�CH�AA/����2��RSD�x"ѡb�w!: ;_T��PRO��OÖ� EM�_��8u�q u�q���DI�0e�RAIL�AC��C�MƐLOԠdC��:anq��wq�����PR��SLQ��pfC�ѷ 	��F�UNCŢ�rRIN�kP+a�0 ��!RA� >R 
Я��ίWAR�BLFQ��A������DA�����L�Dm0�aB9��nqBTIvrbؑ��μPRIAQ1�"AFS�P�!�����`(%b���M�I1UÇDF_j@��y1°L�ME�FA�@HRDiY�4��Pn@RS@Q��0"�MULSE�j@f�b�q �hX��ȑ���$.A[$�1$c1Ó~���� x~��EG� ݓ�q!AR����09>B�%AXE��ROB���W�A4�_�-֣S�Y���!6��&S�'W�R���-1���ST�R��5�9�E��C 	5B��=QB90`�@6������OT�0�o 	$�ARY�8�w20���	%�F�I��;�$LINQK�H��1�a_63��5�q�2XY�Z"��;�q�3@��1��2�8{0B�{`D��� CFI���6G��
�{�_J���6��3aOP_dO4Y;5�QTBmAd"�BC
�z�DU"�z66CTURN3��vr�E�1�9�ҍGFL�`���~ �@�5<:y7�� 1�?0%K�Mc�68Cb�8vrb�4�ORQ��X �>8�#op������wq�Uf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W�� �Tυ� ;����QH� !`�ҽ��U�Q�WkeK#�kecXER��	BGE	0��S�dAWa Ǣ:D���7!�!AX�rB!{q��1 uy-!y�pz�@ z�@z6Pz\Pz�  z1v�y�y� +y�;y�Ky�[y��ky�{y��y�q�yD7EBU��$�����L�!º2WG`  A!B!�,��SV���� 
w���m���w� ���1���1���A���A ��6Q��\Q���!�m@���2CLAB3B��U�����S � ÐER���� �� $�@� Aؑ!p�PO��Z�q0�w�^�_MRAȑ�/ d  T�-��ERR��TYz�B�I�V3@�cΑ'TOQ�d:`L� �d�2�]�X�C[! /� p�`T}0i��_V1�r�a'�
4�2-�2<����@Pq�����F�$W���g��V_!�l�$��P����c��q"�	��SFZN_C;FG_!� 4��?� ��|�ų����@�ȲW� p ��\$� � n���Ѵ��9c�Q��(��FA�He�,�XE�DM�(�����!s��Q�g�P{RV HEL}Lĥ� 56��B_BAS!�RSQR��ԣo �#S��T[��1r�%��2ݺU3ݺ4ݺ5ݺ6ݺ�7ݺ8ݷ��ROO0I䰝0�0NLK!�C�AB� ��ACK��IN��T:�1�! p�@ z�m�_PU!�CO� ��OU��P�� Ҧ) ��޶��T�PFWD_KAR�ӑ��RE~��P8��(��QUE������P
��CSTOPI_AL�����0B�p���㰑�0SEMl�db�|�M��d�TY|�3SOK�}�DI����p�(���_TM\�MANRQ�ֿ0E�+�|�$KEYSWITCHB�	����HE
�BEAT4����E� LEҒ��
�U��FO�����_O_HOM�O�7REF�PPRz�(�!&0��C+�OA��ECO��B�rI�OCM�D8׵�p]���8�` � D�1$����U��&�MH��<�P�CFORC���� �'����OM>�  � @V��*|�U,3P� 1-�`ʀ 3-�4��NP�X_ASǢ� 0�ȰADD����$�SIZ��$VA�Rݷ TIP]�\�2�A򻡐��Ȑ]�_� �"S꣩!C<ΐ��FRIF⢞�aS�"�c���NF�ҸV ��` � x�`S�I�TES�R6SSKGL(T�2P&���AU�� ) STMTdQZPm 6BW�P�*SHOWb���SV�\$�� ���A00P�a� 6�@�J�T�U5�	6�	7�	8�	9�	A�	� �!�'��C@�F�0u �	f0u�	�0u�	�@�u[Pu%121�?1L1Y1f1�s2�	2�	2�	2��	2�	2�	2�	2�22%222�?2L2Y2f2�s3P)3�	3�	3��	3�	3�	3�	3�33%323�?3L3Y3f3�s4P)4�	4�	4��	4�	4�	4�	4�44%424�?4L4Y4f4�s5P)5�	5�	5��	5�	5�	5�	5�55%525�?5L5Y5f5�s6P)6�	6�	6��	6�	6�	6�	6�66%626�?6L6Y6f6�s7P)7�	7�	7��	7�	7�	7�	7�77%727�?7,i7Y7Fi7�s�VP�UPD>��  ��|�԰��YSLOǢ� � z��и����o�E��`>�^t��АAcLUץ����CU��z�wFOqID_L��ֿuHI�zI�$F�ILE_���t���$`�JvSA��� �h���E_BLC�K�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� ��LA��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ���TBCu�C� ��X -$�LENi��v�������I��G�LOW_A�XI�F1��t2�X�M����D�
 ��I�� ��}�TOR�����Dh��� L�=��⇒�s���#�_�MA`�ޕ��ޑT#CV����T��� &��ݡ����J�����IJ����Mo���J�Ǥ� �������2���� v�����F�JK���VKi�Ρv�Ρ3f��J0�ңJJڣ;JJ�AALң�(ڣ��4�5z�&��N1-�9���␅�L~�_Vj�������� ` �GRO�U�pD��B�NF�LIC��REQ�UIREa�EBU`A��p����2¯������c�� �\��APPR��C����
�EN�CsLOe��S_M �v�,ɣ�
���� ���MC�&���Ng�_MG�q�C� ��{�9���|�BRK�z�NOL��|ĉ R��_LI|��Ǫ�k�	J����P
���ڣ��@���&���/���6�Ŕ6��8��r��Ə� ��8�%�xW�2�e�PATHa׀z�p�z�=�vӥ�ϰ�6x�CN=�CA����l�p�IN�UC���bq��CO�UM��YZ������qE%���2�������PAYLO�A��J2L3pR_AN��<�L��F�B��6�R�{�R_F2LgSHR��|�LOG���р��ӎ���ACRL_u�������.���9H�p�$H{���FLEX
��J>�� :�/� ���6�2�����;�M�_�F16����n��� ������ȟ��Eҟ� ����,�>�P�b�� �d�{����������H��5�T��X�� v���EťmFѯ �������&�/��A�S�e�+p�x�� � ������j�4pcAT����n�EL S �%øJ���ʰ;JE��CTR�Ѭ��TN��F&��HA_ND_VB[
�ܤpK�� $F2�{�6� �rSWi���("U��� $$	Mt�h�R��08��@<b 35��^6A�p3�kƈ�q{9t�A�̈p��A���A�ˆ0��U���D*��D��P��G��ICST��$A��$AN��DYˀ�{�g4�5D� ��v�6�v��5缧�^�@��P������#�,�5�>�(#�� &0�_�ER!V9�SQOASYM��] ��¤��x��ݑ���_SHl�������sT�(����(�:�JA���S�pcir��_VI�#�Oh9�``V_UN!I��td�~�J���b �E�b��d��d�f��n���������uN$���(!�H����3��"CqEN� a�SDI��>�Obt DќDpx�� ��2IxQA�q��q��-��s� �� s����� �^�OMME�h�rr/�TVpPT�P  ���qe�i����P��x ��yT�Pj� �$DUMMY9��$PS_��R�Fq�sp$:� �s���!~q� XX����K�STs�ʰ�SBR��M21_�Vt�8$SV_E�Rt�O��z���CLRx�A  O�r?p? �Oր � D ?$GLOB���#LO��Յ$�o���P�!SYSADqR�!?p�pTCHM0 � ,����oW_NA��/��e�os�TSR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T>D�XSCRE�ƀ5�� ��STF���#}�pТ6�sq] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��tC�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$sqVSHIF��|s�P�p�6��s���R���OSU�RW�pRADIz��2�_�q�h�g!� �q)�LUza�$OUTPUT_3BM��IML�oRp6(`)�@TIL<'SCO�@Ce�; ��9��F��T��a ��o�>�3�����w�2u�b�V�zu✫�%�DJU��|#_�WAIT������%ONE���YBOư ��� $@p%�C�S�Bn)TPE��NE�C��x"�$t$���*B_T��R��%�qRH� ���sB�%�tM�+ ��t�.�F�R!݀���OPm�MAS�_�DOG�OaT	�D�����C3S�	�O2DE�LAY���e2JO ��n8E��Ss4'#J�aP`6%�����Y_��O2$��2���5��`?� b�ZABC~S��  $�2��J�
sp�$$C�LAS������Aspb�'@@VI�RT��O.@ABS��$�1 <E�� < *AtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v�����M@�[�AXLր�&A�ndC  ���IN��ā��PRE������LARMRECOV <Il䂥�NG�� \K	 A   J�|\�M@PPLIC��?<E�E��Handlin�gTool �� �
V7.50P�/28[�  �Xۭ��
�_S�W�� UP*A�� ��F0ڑ����A��0�� 20���*A���:���(��FB �7DA5�� ~'@Y�@�����None������� ��T���*A4I�x�l�_��V����g�UTOB�ค��~��HGAPON8@蕮LA��U��D 1-<EfA����������� Q 1EשI Ԁ�� Ԑ�:�i�n����#B�)B ����\�HE�Z�r�?HTTHKY��$B I�[�m�����	�c� -�?�Q�o�uχϙϫ� ���������_�)�;� M�k�q߃ߕߧ߹��� �����[�%�7�I�g� m����������� ��W�!�3�E�c�i�{� ��������������S /A_ew�� �����O+ =[as���� ���K//'/9/W/ ]/o/�/�/�/�/�/�/ �/G??#?5?S?Y?k? }?�?�?�?�?�?�?CO OO1OOOUOgOyO�O �O�O�O�O�O?_	__`-_K_Q_��(�TO4��s���DO_CLE�AN��e��SNM ; 9� �9o�Ko]ooo�o�DSP�DRYR�_%�HI��m@&o�o�o# 5GYk}���`�"���p�Ն �ǣ�qXՄ��ߢ��g�PLUGGҠ�Wߣ���PRC�`B`"9��o�=�OB��o^e�SEGF��K�� ����o%o����#�85�m���LAP�oݎ ����������џ������+�=�O�a���T�OTAL�.���U�SENUʀ׫ �X���R(�RG_S�TRING 1~��
�M���Sc�
��_ITwEM1 �  nc� �.�@�R�d�v����� ����п�����*��<�N�`�r�I/�O SIGNAL���Tryou�t Mode��Inp��Simu�lated�O�ut��OVE�RR�` = 10�0�In cy�cl���Pro?g Abor������Status��	Heartb�eat��MH �FaulB�K�AlerUم�s߅ߗߩ������������ �S���Q��f�x� ������������� �,�>�P�b�t�������,�WOR������ V��
.@Rd v��������*<N`PO��6ц��o�� ���//'/9/K/ ]/o/�/�/�/�/�/�/8�/�/�DEV�*0 �?Q?c?u?�?�?�? �?�?�?�?OO)O;O�MO_OqO�O�O�OPALTB��A���O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo8(o:o�OGRI�p�� ra�OLo�o�o�o�o�o �o*<N`r ������`o��RB���o�>�P�b� t���������Ώ��� ��(�:�L�^�p����PREG�N��.� �������*�<�N� `�r���������̯ޯ����&����$A�RG_��D ?	����i���  	]$��	[}�]}����Ǟ�\�SBN_�CONFIG �i�������C�II_SAVE � ��۱Ҳ\�T�CELLSETU�P i�%H?OME_IO�͈�?%MOV_�2ώ8�REP���V�U�TOBACK
��ƽFRA;:\�� �Ϩ���'`!��������� ����$��6�c�Z�lߙ��Ĉ�������������!� ����M�_�q���� 2���������%�7� ��[�m��������@� ������!3E$���Jo����\���INI�@���ε��MESS�AG����q��ODE_D$����O,0.��PAUS��!�i� ((Ol������ �� /�//$/Z/�H/~/l/�/�'akTSK  q������UPDT%�d�0;WSM_C5F°i�еU�>'1GRP 2h�93+ |�B��A�/S��XSCRD+11
N1; ����/ �?�?�? OO$O��� �?lO~O�O�O�O�O1O �OUO_ _2_D_V_h_��O	_X���GROU�N0O�SUP_N5AL�h�	�ĠV�_ED� 11;
� �%-BCKEDT-�_`�!oEo%���a��o��e���ߨ���eA2no_˔o�o�b����ee�o"�o�oED3 �o�o ~[�5GED4�n#��� ~�j���ED5 Z��Ǐ6� ~���}���ED6����k�ڏ� ~G���!�3�ED7 ��Z��~� ~�V�şןED8F�&o��Ů�}����i�{�ECD9ꯢ�W�Ư
}03�����CRo�� ���3�տ@ϯ����P~�PNO_DEL�_��RGE_UNUS�E�_�TLAL_OUT q�c�QWD_ABOR� ��΢Q��ITR_R�TN����NON�Se���CA�M_PARAM �1�U3
 8�
SONY XC�-56 2345�67890�H �� @���?}���( АVڪ|[r؀~�X�H�R5k�|U�Q�߿�R�57����Aff���KOWA S_C310M|[r�}̀�d @6� |V��_�Xϸ���V� �� ���$�6��Z�l���CE_RIA_UI857�F�1���R|]��_�LIO4W=� ��P<~�F<�GP ]1�,���_�GYk*C*  ���C1� 9� @Ң G� �CLC]�� d� l� s�R�� ��[�m� v� � �� �� +C�� �"�|W���7�HEӰONFI�� ��<G_PRI 1�+P�m®/ ��������'CHKPAUS� w 1E� ,� >/P/:/t/^/�/�/�/ �/�/�/�/?(??L?�6?\?�?"O��x���H�1_MOR��� �0�5 	 �9 O�?$OOHO6K�2	���=9"�QI?55��C�PK�D�3P������a�-4�O__|Z
�OG_�7�PO�� ��d6_��,xV�ADB����='�)
mc:cpmidbg�_|`��S:�  � +���Up�_)o�S�  �  	A���R�P�_mo8j�"�Koo�o9i+�)�Փog�o�o
�m��of�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`)ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCo��C|��Cq�D��C����C�{iSZE@D���F.��F���E⚵F?,E�ٙ�E@�F�N�IU���I?O�I<#�I6�I洤SY���vqG��T�Em�)�.��)��)��<�q�G�x�2��Ң �� a�D��j���ES\E@E�X�EQ�E�JP F�E�F� G�ǎ�^F E�� F�B� H,- Ge��H3Y����  >�33 ����xV  n42xQ@��5Y��8B� A�AST<#�
�� �_'�%��wR_SMOFS���~�2�yT1�0DE 3�O@b 
�(�;;�"�  <�6��z�R���?�j�C�4��SZm� W�(�{�m�C��B-G��Cu�@$�q��T�{�FPROG !%i����c�I��� ��Ɯ�f�KEY_TOBL  �vM�u�� �	
��� !"#$%&'�()*+,-./�01c�:;<=>�?@ABC�pGH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������p���͓���������������������������������耇����������������������!j�LCK�.�j���STAT����_AUTO_�DO���W/�IN?DT_ENB߿21R��9�+�T2w�X�STOP\߿2TR�Ll�LETE�����_SCREEN� ikc�sc��U��MME�NU 1 i  <g\��L�SU +�U��p3g����� ��������2�	��A� z�Q�c����������� ����.d;M �q����� �N%7]�m ���/��/ J/!/3/�/W/i/�/�/ �/�/�/�/�/4??? j?A?S?y?�?�?�?�? �?�?O�?O-OfO=O OO�OsO�O�O�O�O�O�_�O_P_Sy�_M�ANUAL��n�DwBCOU�RIG��>�DBNUM�p���<���
�QPXW�ORK 1!R� ү�_oO.o@oRk�Q__AWAY�S��/GCP ��=��df�_AL�P�db�RYв������X_�p 1}"�� , 
�^@���o xvf`MT��I^�rl@�:sON�TIM�����ɼZv�i
õ�cMO�TNEND���dR�ECORD 1(�R�a��ua�O� �q��sb�.�@�R� �xZ�������ɏۏ 폄���#���G���k� }�����<�ş4��X� ��1�C���g�֟�� ������ӯ�T�	�x� -���Q�c�u������� ���>����)Ϙ� Mϼ�F�࿕ϧϹ��� :�������%�s`Pn&� ]�o��ϓ�~ߌ���8� J�����5� ��k� ���ߡ��J�����X� �|��C�U������ ����0�����	���dbTOLEREN�CqdBȺb`L��͐PCS_CFG� )�k)wd�MC:\O L%0?4d.CSV
�p�c�)sA �CH
� z�p)~����hMRC_OUT *�[�`+P ?SGN +�e�r���#�10-M�AY-20 10�:59*V17-F;EBj9:0rv PQ�8��)~�`pa��m��PJP���VERSIO�N SV�2.0.8.|EF�LOGIC 1,^�[ 	DX�P�7)�PF."PROG�_ENB�o�rj U�LSew �T�"_?WRSTJNEp�V��r`dEMO_OPT_SL ?	�e�s
 	R575)s7)�/??*?�<?'�$TO  ��-��?&V_@pE�X�Wd�u�3PA�TH ASA�\�?�?O/{ICTZ�aFo`-�gd>segM%&A�STBF_TTS��x�Y^C��SqqF��PMAU� t/XrMKSWR.�i6.|S/�Z!D_N�O 0__T_C_x_g_�_�t�SBL_FAUL�"0�[3wTDIAbU 16M6p�A�123456�7890gFP ?BoTofoxo�o�o�o �o�o�o�o,>�Pb�S�pP�_ ���_s�� 0`� ����)�;�M�_� q���������ˏݏ�|)UMP�!� �^�TR�B�#+��=�PMEfEI�Y_�TEMP9 È��3@�3A v�UNI��.(YN_BRK� 2Y)EMG?DI_STA�%W�!bՐNC2_SC/R 3��1o"� 4�F�X�fv�������0��#��ޑ14�����)�;�����ݤ5�����x�f	 u�ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/߭P� b�t�� ��xߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N���r� �������������� &8J\n�� ������" `�FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/4?,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O?�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�O�O �o�o�o
.@R dv������ ���*�<�N�`�r� ���o����̏ޏ��� �&�8�J�\�n����� ����ȟڟ����H��ETMODE 1�6��� 
��ƨ
R�d�v�נ�RROR_PROoG %A�%�:����  ��TABL/E  A�������#�L�RRSEV_NUM  ��Q��K�S����_AUTO_EN�B  ��I�Ϥ_;NOh� 7A�{�}R�  *�������������^�+રĿֿ迄�HIS�O���I�}�_ALMw 18A� �;�����+�e�w� �ϛϭϿ��_H���  A���|���4�TCP_VER� !A�!����$�EXTLOG_R�EQ��{�V�S�IZ_�Q�TOL � ��Dz��{A Q�_BWD��p��r���n�_DI��7 9��}�z�x��m���STEP�����4��OP_DO����ѠFACTORY_TUN��dG�EATURE� :����l��HandlingTool ���  - CE�nglish D�ictionar�y��ORDE�AA Vis�� ?Master����96 H��nal?og I/O����H551��uto� Softwar�e Update�  ��J��mat�ic Backu�p��Part�&�ground �Edit��  8�\apCam�era��F��t\;j6R�ell����LOADR�omm���shq��TI"� ��co��
!� o���pane��� 
!��t�yle sele�ct��H59��n�D���onitorf��48����tr��?Reliab����adinDiagnos"�����2�2 ual Ch�eck Safe�ty UIF l�g\a��hanc�ed Rob S�erv q ct�\��lUser sFrU��DIF���Ext. DIOm ��fiA d���endr Err� L@��IF�rd��  �П�90���FCTN MeneuZ v'��74� �TP In��fa�c  SU (�G=�p��k Excn g�3���High-Spe�r Ski+�  s�O�H9 � mmun�ic!�onsg�tFeur� ����V�����conn���2��EN��In{crstru�����5.fdK�AREL Cmd7. L?uaA� �O�Run-TiN� Env����K� ���+%�s#�S/W���74��Lice�nseT�  (�Au* ogBoook(Sy��m)���"
MAC�ROs,V/Of�fse��ap��MqH� ����pfa5��MechStop� Prot��� �d�b i�Shiyf���j545�!�xr ��#��,[��b ode Sw�itch��m\eҙ!o4.�& p#ro�4��g��Multi-T7�G��net.�Pos Regi���z�P��t Fsun���3 Rz1��Numx ������9m�1�  Adjyuj��1 J7�7�* ����6tat�uq1EIKR�DMtot��scove�� ��@Bxy- }uest1��$Go� � U5\?SNPX b"��x�YA�"Libr�����#�� �$~@h��pd]0�Jts in VCCM�����0�  �u!��23 R�0�/I�0�8��TMILIB^�M J92�@P�gAcc>�F�97��TPTX�+�BRS�QelZ0�M8 Rpm��q%��692���Unexcept�r motnT  �CVV�P���KC�����+-��~K  �II)�VSP C7SXC�&.c�� e��"�� t�@W9ew�AD Q�8bsvr nmen�@��iP� a0y�0��pfGridAplay !� nh�@�*�3R�1M-10iA(B201 �`�2V"  F���sc{ii�load��/83 M��l�����Guar�d J8	5�0�mP'�L`���;stuaPat�&]$�Cyc���|0oryi_ x%Data'P3qu���ch�1�h�g`� j� RLJ�am�5���IMI� De-B(\A�cP�" #^0C  �etkc^0assswo%q�)650�A1pU�Xnt��P�ven�CTqH�5��0YELLO�W BO?Y��� A;rc�0vis��Ch�WeldQc�ial4Izt�Oap� ��gs�` 2@�ma��poG yR�jT1 NE�#HT�� xyWb��! �p�`gd`���p\�� =P��JPN A7RCP*PR�A��� OL�pSup̂fil�p��J��� ��cro�670`�1C~E�d��SS�p]e�tex�$ �P�� So7 t� ssKagN5 <Q�BP:d� �9 "0�QrtQ�C��P�l0dpn��笔�rpf�q�e�pp�mascbi�n4psyn�' �ptx]08�HEL�NCL VIS? PKGS �Z@�MB &��B J�8@IPE GE�T_VAR FI�?S (Uni� L�U�OOL: AD}D�@29.FD�TiCm���E�@DVp���`A�ТNO WTWTEST ��� f�!��c�FOR� ��ECT �a!�� ALSE AL�A`�CPMO-1�30��� b D: �HANG FRO�Mg��2��R70�9 DRAM A�VAILCHEC?KS 549��m�VPCS SU֐�LIMCHK��P��0x�FF POS� F�� q8�-12 CHAR�S�ER6�OGRA� ��Z@AVEH�A;ME��.SV��В�אn$��9�m "�y�TRCv� SH�ADP�UPDAT� k�0��STAT�I��� MUCH� ���TIMQ �MOTN-003���@OBOGU�IDE DAUG�H���b��@$to�u� �@C� �0��P�ATH�_�MOV{ET�� R64���VMXPACK �MAY ASSE�RTjS��CYCL�`�TA��BE C�OR 71�1-�A�N��RC OPT?IONS  �`���APSH-1�`fix��2�SO��B�0�XO򝡞�_T��	��i��0j��du�byz p wa��y�٠#HI������U�pb XSPD TB/��F� \hchΤBl0���END�CE�0�6\Q�p{ smOay n@�pk���L ��traff�#�	� ��~1fr�om sysva_r scr�0R� ���d�DJU���H��!A��/��SET� ERR�D�P7�����NDANT �SCREEN U�NREA VM 4�PD�D��PA����R�IO JNN��0�FI��B��G�ROUNנD Y��Т٠�h�SVI�P 53 QS��D�IGIT VERqS��ká�NEW�� P06�@C�1I�MAG�ͱ���8�� DI`���pSS�UE�5��EPLA�N JON� DE�L���157QאD��CALLI���Qx��m���IPND}��IMG N9 P�Z�19��MNT/Υ�ES ���`LocR Hol߀=��2:�Pn� PG:��=�M��can����~С: 3D mE2�view d XL��ea1 �0b�pwof Ǡ"HCɰ��ANNOT A�CCESS M �cpie$Et.Qs� a� loMdFl�ex)a:��w$qmWo G�sA9�-'p�~0��h0pa��eJ? AUTO-�0���!ipu@Т<ᡠI/ABLE+� 7�a ?FPLN: L�gpl m� MD<��VI�и�WIT �HOC�Jo~1Q�ui��"��N��U�SB�@�Pt & remov���D�v�Axis FT_t7�PGɰCP:�OS-144 � ?h s 268QՐ�OST�p  CR�ASH DU��$�P��WORD.$>�LOGIN�P���P:	�0�046 issueE�H�: Slow +st�c�`6����໰IF�IMPR���SPOT:Wh84���N1STY��0�VMGR�b�N�CkAT��4oRRE��9 � 58�1���:%�RTU!Pe -\M a�SE:�@pp�H��AGpL��m�@all��*0a�O�CB WA���"3 CNT0 T9D�WroO0alarqm�ˀm0d t�0M�"0�2|� o�Z@�OME<�� ��E% w #1-�SRE���M�st}0g   �  5KANJ�I5no MNS�@�INISIToALIZ'� E��f�we��6@� dr��@ fp "��S�CII L�afa�ils w��SYSTE[�i���  � Mq�1QG;ro8�m n�@vA����&��n�0q���RWRI OF �Lk��� \ref�"�
�up� de-�rela�Qd 0k3.�0SSchő�betwe4�IN�D ex ɰTPFa�DO� l� ��ɰGigE�sop�erabil`p l,��HcB��@]��le�Q0cflxpz�Ð���OS {�����v4pfigi GCLA�$�c2�7H�� lap�0ASBֻ If��g�2 lC\c�0�/�E��? EXCE 㰁�!P���i�� o0��Gd`]Ц�fq�l �lxt��EFal���#0�i�O�Y�n�CwLOS��SRNq1+NT^�F�U��Fq�KP�ANIO V7�/ॠ1�{����D�B �0��ᴥ�EDN��DET|�'� �}bF�NLINEb�GBUG�T���C"R�LIB��A��ABC JARKY@���� rkey�`I)L���PR��N��ITWGAR� D$�R  �Er *�T��a��U�0��h�[�ZE �V� TASK op.vr�P2" 8.�XfJ�srn�S谎�dIBP	c���B�/��BUS��UNN� j0-�{��c�R'���LOE�DIVS�CULs$cb����BW!��R~�0W`P�����IT(঱�tʠ�OF��UN#EXڠ+���p�Ft}E��SVEMG3`NML 505� �D*�CC_SAF�E�P*� �ꐺ� P�ET��'P�`�F  !���IR����c� i S>� K��K��H GUNCH�G��S�MECH���M��T*�%p6�u��tPORY L�EAK�J���S�PEgD��2V 74\GRI��Q�gޙ�CTLN��TR�e @�_�p ���EN'�IN������$��̸r��T3)�i�ST%O�A�s�L��͐!X	���q��Y� ���TO2�J m��0F0<�K����DU�S��%O��3 9�J �F�&���SSVG�N-1#I���RS	RwQDAU�Cޱ� �T�6�g��� 3�]���BRKCTR/"� �q\j5��_�Q�S�q�INVJ0D ZO �Pݲ���s��г�Ui �ɰ̒�a�DUAL�� J50e�x�RVO117 AW��TH!Hr%�N�24�7%�52��|�&aol ���R���at�S�d�cU���P,�LE�R��iԗQ0�ؖ  CST���Md�Rǰ�t� \fosB�A��0Np�c����{�U>��ROP 2�b�p}B��ITP4M��b !AUt c0< >� plete�N@�� z1^qR63�5 (AccuC�al2kA���I)C "�ǰ�1a\�Ps��ǐ� bЧ0P��������ig\cbacul "A3p�_ �1��ն���et�aca��AT���PaC�`�����_p��.pc!Ɗ��:�c�ircB���5�tl0��Bɵ�:�fm+��Ċ�V�b�ɦ�r�upfrm.����ⴊ��xed��Ί�~�pe�dA�D �}b�pt�libB�� �_�r!t��	Ċ�_\׊���6�fm�݊�oޢ� e��̆Ϙ���c�Ӳ�b5�j>�����tcȐD��	�r����mm 1��T�sl^0��T�1mѡ�#�rm3��qub Y�q�std}�f�pl;�&�ckv�=�r�vf�䊰��9�cvi����ul�`h�0fp�q �.f���� daq; i D�ata AcquWisi��n�
�h�T`��1�89����22 DMCM� RRS2Z�75���9 3 R71Y0�o59p5\�?��T "��1 #(D�T� nk@�� ������E Ƒȵ��Ӹ��etdmm ��ER����gE��1�q\mo?۳�= (G���[(

�2��` ! �@JMA�CRO��Skip?/Offse:�a���V�4o9� &qR�662���s�H�
 6Bq8�����9Z�43 J77z� 6�J783��o ��n�"v�R5�IKCBq2 PgTLC�Zg R�w3 (�s, �0������03�	з�JԷ\sfmnmc "MNMC�����ҹ�%mnf�F�MC"Ѻ0ª et�mcr� �8����� ,[��Df�   �874\prdq�>,jF0���ax�isHProce�ss Axes �e�rol^PRA�
�Dp� 56 J8m1j�59� 56oa6� ���0w�690 s98� [!IDV�1Ĵ�2(x2��2ont�0�
����m2���?C��etis "ISD��9��^ FpraxRAM�Pp� D��defB��,�G�isbasicHB�@޲{6��� 708�6��(�Acw:������D
��/,��AMOX�� ��D@vE��?;T��>Pi� �RAFM';�]�!PAM �V�W�Ee�U�Q'
�bU�75�.�ce�Ne� nterfGace^�1' 5&!�54�K��b(Devam±�/�#���/<��Tane`"DNE�WE���btpdnu�i �AI�_s2�d_rsono���b�AsfjN��bdv_arFvf�xhpz�}w抰hkH9xstc8��gAponlGzv{�ff��r����z�3{q'Td>p�champr;e�p� ^5977��	܀�4}0��mɁ�/������lf�!�pcchmp]aMP&B�� �mpev������pcs��YeS�� _Macro�OD��16Q!)*�:$�2U"�_,��Y�(PC  ��$_;������o��J��gegemQ@GE�MSW�~ZG�ges�ndy��OD�ndd1a��S��syT�KɆ��su^Ҋ���n�mx���L��  ����9:p'ѳ޲��sp?otplusp����`-�W�l�J�s��t8[�׷p�key�ɰ��$��s�-Ѩ�m���\�featu 0FEqAWD�oolo�srn'!2 p����a�As3��tT.� (N. A.)�@�!e!�J# (j��,��oBIB�oD �-�.�n��k9�"AK��u[-�_���p� "PSEqW��~��wop "sE� ��&�:�J������y� |��O8��5��Rɺ�� ��ɰ[��X������ �%�(
ҭ�q HL�0k�
�z�a!�B�Q�"(g�Q��� ��]�'�.�����&���`<�!ҝ_�#��tpJ� H�~Z��j�����y�� ����2��e������Z ����V��!%���=��]�͂��^2�@iRV�� on�QYq͋J�F0� 8ހ�`�	(|^�dQueue����X\1�ʖ`�+F1tp/vtsn��N&��f�tpJ0v �RDV �	f��J1 Q����v�en��kvs�tk��mp��btkclrq���get����r<��`kack�XZ��strŬ�%�satl��~Z�np:! �`���q/�ڡ6!!l�/Yr�mc�N+v3�_� �����.v�/\jF��� �`Q�΋ܒ�N5?0 (FRA��+���͢frapar�m��Ҁ�} 6�J�643p:V�ELS�E
#�VAR �$SGSYSCF�G.$�`_UNITS 2�DG~°@��4Jgfr��4A�@FRL-��0ͅ�3ې�� �L�0NE�:�=�?@@�8�v�9~Qx304�8�;�BPRSM~Q�A�5TX.$VNUM_OL��5��D�J507��l� Functʂ"qwAP8��琉�3 H�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6N�k�AP����S��"T�PPR���QA�prnaSV�ZS��AS^8Dj510U�-�`�cr�`8 ��ʇ�DJ�R`jYȑH  k�Q �PJ6�a�21��48A�AVM 5�Q�b0y lB�`TUP xbJ545 `b��`616���0�VCAM 9��CLIO b1��5 ���`MSC�8�
rP R`\s�STYL MN{IN�`J628Q;  �`NREd�;@��`SCH ��9pD�CSU Mete>�`ORSR Ԃ�a�04 kREI�OC �a5�`542�b9vpP<�nP�a��`�R�`7�`�MASK Ho��.r7 �2�`OCO	 :��r3��p�b�p����r0X��a�`13�\mn�a39 H�RM"�q�q���LCHK�uOPLsG B��a03 �q=.�pHCR Ob�p=CpPosi�`fP�6 is[rJ5594�òpDSW�bM�qD�pqR�a37 }Rfjr0 �1�s4 �R�6�7��52�r5 \�2�r7 1� P6�~��Regi�@�T�uFRDM�uStaq%�4�`930�u�SNBA�uSHL]B̀\sf"pM��NPI�SPVC��J520��TC��`"MNрTMI�L�IFV�PACy W�pTPTXp�6.%�TELN oN Me�09m3?UECK�b�`�UFR�`��VCO�R��VIPLpq8�9qSXC�S�`VV9F�J�TP �q���R626l�u S��`Gސ�2IGsUI�C��PGSt�=\ŀH863�S�qX�����q34sŁ684���a�@b>�33 :B��1 T���96 .�+E�51� y�q53�3�b1� ���b1 n�jr9y ���`VAT ߲�q75 s�F��`�s�AWSM��`TO3P u�ŀR52p����a80 
�ށXY� q���0 ,b�`8k85�QXрOLp�}�"pE࠱tp�`L�CMD��ETSS����6 �V�CP�E oZ1�VRC�d3
�NLH�h��0c01m2Ep��3 f���p��4 /165�C��6l���7PR���008 tB��9� -200�`U02�pF�1޲1 ��޲A2L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�~J�7 rbcfA��L�8\PC����"�3!2m0u�n�K�Rٰn�5 5EW
n�s9 z��40 kB���3 ��6ݲ�`0/0iB/��6�u��	7�u��8 µ�������sU0�`�t �1 �05\rb��2 �E���K���j���5˰��60��a�HУ`:�63�jAF�_���F�#7 ڱ݀H�8�eH�L���cU0��7�p���1u��8u��9� 73������D7�� ��5t�97 ���8U�1��2��1R�1:���h��1np��"��8(�U1��\pyl��,࿱v ��.B�854��1V���ZD�4��im��1� <���>br�3pr�q4@pGPr�6 B��H�цp��1����1�`�͵155ض157 �2��62�S�����1b��2����1dΠ"�2���B6`2�1<c�4 7B��5 DR��8_�B/���187 uJ�8w 06�90 rB�n�1 (��202_ 0EW,ѱ2^�4�2��90�U2�p�2���2 b��4��2N�a"RB����9\��U2�`w�l���4 60Mp��7������Xb�s
5 ��3��x��pB"9 3 ��؆�`ڰR,:7  �2��V�2��5���2�^��a^9���qr����n�5����5�D��"�8a�Ɂ}�5B�"��5����`UA���d� ��86 �6 S��0��5�p�2�#�529 �2^�b1P�5~�2`���T&P5��8��5���u�!�5��ٵ544J��5��R�ąP nBX^z�c (�4�������U5J�V�5��1�1^��%����:��5 b21��lgA��58W82� �rb��5N�E�58�90r� 1�95 �"������c8"a�@�|�L ���!J"5|6��^!�6��B�"�8�`#��+�8%�6�B�AME�"1 i�C��622�Bu�6hV��d� 4��84�`�ANRSP�e/S� C�5� �6� ��� \� �6� �V� �3t��� T20CA�R��8� Hf� �1DH�� AOE� ��� ,[|��� �0\�� �!64�K��ԓrA� �1 (�M-7�!/50T@�[PM��P�Th:1 �C�#Pe� �3�0� }5`M75T"� �D8p� �0Gc� u��4��i1-710i��1� Skd�7j�?6�:-HS,� �RN��@�UB�f�X�=m�75sA*A6an����!/CB�B2.6A  �0;A�CIB�A�2�QF1ԣUB2�21� /7!0�S� �4����Aj1�3p���r#0 B'2\m*A@C��;bi"i1K�u"A~AAU� ?imm7c7��ZA�@I�@�Df�A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A�EA��5B�4>\77
B7@=Q�D�2�Q$B�E7�CJ�D/qAHEE�W7�_ |`jz@� 2�0�EBjc7�`�E"l7�@�7�A
1�E�V~`�W2�%Q�R9ї@0L_�#����"A���b��9H3s=rA/2�R5 nR4�74rNUQ1ZU�A�s\m9
1M92�L2�!F!^Y�ps� 2cci��-?�qhimQ �t  w043�C�p2�mQ0�r�H_ �H20�Evr0�QHsXBSt62�q`s������ ��Pxq3g50_*A3I)�2��d�u0�@� '4TX��0�pa3i1A3`sQ25�c��st�r"�VR1%e�q0
�� j1��O2 �A�UEi�y�.�‐ �0Ch20$CXB79#A�ᓄM 8Q1]�~�� 9�Q�� ?PQ��qA!Pvs� 5 	15aU���?PŅ�8��ဝQ9A6�zS*�7�qb5�1����QN��00P(��V7]u �aitE1���ïp?7�� !?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ���y00\ry�"�R2BL�tN  ���� �1D�f��2�qeR�5����_b�3�X]1m1lcqP1�a�E�Q� �5F����!5���@M-16Q�� f���r� �Q�e� ��� PN�LT_�1��i1��94�53��@�e�|�b1l>F1u*AY2�
��R8�Q����RJ�cJ3�D}T� 85
Q g�/0��*A!P�*A��Ȑ𫿽�2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt ]1^u�ajrI�B�����~�|I�b��yI�\m�Qb�I�uz�A�c3A�pa9q� B6S��S0��m���}�85`N�>N�  �(M ���f1���6����16�1��5�s`�SC��U��A����5\s�et06c����10�y�h8��a6���6��9r�2HS @���Er���W@}�a�� I�lB���Y�ٖ�m�u�C����5�B��B��h`�F���X0��@�A:���C�M��AZ��@��4�6i����� e�O�-	���f1�� �F �ᱦ�1F�Y	���T6HL3��U66�~`���U�dU�9D20Lf0��Qv� ��f jq��N������0v
�� ��i	�	��72lqQ2������� �\chngmove.V��d���@2l_arf	�f ~��6������9C��Z���~���kr4�1 S���0��V��t������U�p7n�uqQ%�A]��V�1E\�Qn�BJ�2 W�EM!5���)�#�:�64��F�e50S�\��0�=�PV ���e������E��x���m7shqQSH"U��)��9�!A��(����� ,[��ॲTcR1!��,�60e"=�4F�����2��	 R-��������Ӏ��Ж��4���LS`R�)"�!lOA��Q�) %!� 16�
 U/��2�"2�E�9p��|�2X� SA/i��'�
7F�H�@!B�0 ��D���5V��@2c@VE��p��T��pt���1L~E�#�F�Q��9E�#De/��RT��59���	�A�EiR��������9\m20�20��+�-u�19r4�`�E1�=`O9`@�1"ae��O�2���_$W}am41�4��3�/d1c_stAd��1)�!�`_T���r�_ 4\jdg �a�q�PJ%!~`-�r��+bgB��#c30�0�Y�5j�QpQb1��bq��vB��v25��U�����qm43 � �Q<W�"PsA�� e����t�i�P �W.��c�FX.�he�kE14�44��~6\j4�44�3sj��r�j4up@���\E19�h�PA�T �=:o�APf��coW�o!\�2a��2A;_2��QW2�bF�(�V11�23�`��X,5�Ra21�J*9$�a:88J9X�l5�m1a첚��*���(85�&������ �P6���R,52&AĀ���,fA9IfI50	\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP1���vB)e�m�����1pw� �1Df��2�7�F�KAREL� Use S��F�CTN��� J9a7�FA+�� (�Q`޵�p%�)?�Vj9F?�(�j�Rtk208� "Km�6Q�y�j��iæPr�9�s#���v�krcfp�RC�Ft3���Q��kcc7tme�!ME�g�����6�main�dV�� ��ru��kD��c���o����J�d�t�F �»�.v!rT�f�����E%�!���5�FRj73B�K����UER�HJ�O  J�� (ڳF���F�q�Y�&T��p�F�z��19�tkvBr��ĄV�h�9p�E�y�<�k�������;�v���"CT��f����)�
� ���)�V	�6���! ��qFF��1q���=� ����O�?�$"���$���je��TCP �Aut�r�<520w H5�J53E1k93��9��96�!�8��9��	 �B57�4��52�Je�(�� Se%!Y������u��ma�Pqtoo�l�ԕ������c�onrel�Ftr�ol Relia'ble�RmvCU!��H51����� a�551e"�CNRE¹I�c��&��it�l\sfutst "UTա��"X�\u��g@��i�6Q]V0�B,Eѝ6A� �Q�)C���X@��Yf�I�1|6s@;6i��T6IU��vR�d�
$e%1��2�C#58�E6��8�Pv�iV4OFH58SOeJ� �mvBM6E~O58 �I�0�E�#+@�&�F �0���F�P6a���)/�++�</N)0\tr�1�����P ,[��ɶ�rmaski�m#sk�aA���ky'd��h	A	�P�sDis�playIm�`v�����J887 (�"A��+HeůצprCds��Iϩǅ�h�0pl�2�R2��:�G9t�@��PRD�TɈ �r�C�@Fm��D�Q�A'scaҦ� V<Q0&��bVvbrl�eۀ�@��^S��&5Uf�j38710�yl	��Uq���7�&�p�p���P^@�P�firm Q����Pp�2�=bk�6��r�3��6��tppl��PL���O�p<b�ac�q	��g1J�U�`�d�J��gait_ 9e��Y�&��Q���	��Shap��era�tion�0��RG67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G���q.F�205p�5S��ɜՁ�retsap�BP��O�\s� "G�CR�ö? �qngda�G��V��s"t2axU��Aa]�Ɔbad�_�btp�utl/�&�e���t�plibB_��=�2�.����5���cir�d�v�slp��x�h3ex��v�re?�Ɵ�x�key�v�pm���x�us$�6�gcr��F������[�q�27j92�v�ol7lismqSk�9O|�ݝ� (pl.��$�t��p!o��29$Fo�8��cg7no@�tp�tcls` CLS0�o�b�\�km�ai_B
�s>�v�o	�t�b���ӿ�E�H���6�1enu501:�[m��utia|$�calmaUR��C�alMateT;R51%�i=1]@-��/ V� ��Z�� �fq1�9 "K9E�L����2m�CLMT�q�S#��et �L�M3!} �F�c�n�spQ�c���c_mioq��� ��c_e������su��ޏ �_� �@�5�G�join��i�j��oX���&c`Wv	 ���N�ve��C�clm�&Ao# �~|$finde�0�STD te�r FiLA�NG���R��
p��n3��z0Cen����r,������J�� ��� ���K��Ú�=���_Ӛ��r� "FNDR�� 3����f��tguid��䙃N�."��J�tq �� �������������J����_������c���	m�Z��\fndr.��n#>
B�2p��Z�CP M1a�����38A��� c��6� (���N� B������� 2�$�81��m_���"ex�z5�.Ӛ��c��bSа�e�fQ��	��RB�T;�OPTN  �+#Q�*$�r*$��*$ r*$%/s#C�d/.,P���/0*ʲDPN`��$���$*�Gr�$�k Exc�'IF��$MASK�%93� H5�%H558��$548 H�$4 -1�$��#1(�$�0 E�$��$-b�$��>�!UPDT �B�4 �b�4�2�49�0�4a��3�9j0"M�49�4�  ��4�4t�psh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4��3�adq\�5K97�9":E�ajO l "DQ^E^�3i�D!q ��4ҲO ?R�? ��q�5��T��32rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F���4��.�5y N� �2i�l(in�4��31� JH1�2Q4�251<ݠ�4rmal� �3)�REo�Z_�æOx�����4��^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg0���4�$HCd\�fͲ �eڱ�4�REM���4�yݱ"u@�RER59�32fO��47Z��5lity,�U��e"�Dil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe� =$�^�
E��u�IAymptm�U��BU��vste�y\�3��m e�b�DvI�[�Qu�:F��Ub�*_�
E,�sIu��_ Er���ox���4huse�E-�?�sn�������8FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��@�b���(��1� ��c��Y�R�� �>� P���W��������'�0ɵ�[��͂����  � ,�[@� �A^�bumpšf��B*�Box%��7A�ǰ60�BBw���MC�� (6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`����)��\bbk96�8 "�4�ω�b5b�9va69����'etbŠ��X����F�ed	�F��u�Lf� �sea"������'�\��,���b�Dѽ�o6�H�
�x�$�f���!y���Q[�! tperr��fd� TPl0o� _Recov,��3|D��R642 � 10��C@}s� N@��(U�rro���y�u2r��  �
�  ����$�$CLe� ��������������$z�_DIGIT\������� �.�@�R�d�v����� ����������* <N`r���� ���&8J \n������ ��/"/4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_@�_�_ oo$j��+c�:PRODUCT�M�0\PGSTK�D��V&ohozf9�9��D���$�FEAT_IND�EX��xd���  
�`I�LECOMP ;���#��`�c�SETUP2 �<�e�b� � N �a�c_AP2BCK 1=�i?  �)wh0"?{%&c����Q �xe%�I�m� ��8��\�n���� !���ȏW��{��"� ��F�Տj���w���/� ğS���������B� T��x������=�ү a������,���P�߯ t������9�ο�o� ϓ�(�:�ɿ^��� Ϗϸ�G���k� �� ��6���Z�l��ϐ�� ����U���y���� D���h��ߌ��-��� Q���������@�R� ��v����)�����_� ����*��N��r ��7��m��&�3\�i
pP� 2#p*.cVRc�*���� /��PC�/1/FR6:D/].��/+T�` �/�/F%�/�,�`r/?�*.F�8?	H#&?e<�/�?;STM �2�?�.K ��?�=iPe�ndant Pa'nel�?;H�?@O��7.O�?y?�O:GIF�O�O�5�OoO�O_:JPG _J_�56_��O_�_�	PAN?EL1.DT�_��0�_�_�?O�_2 �_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEIN�S.XML���0\���qCus�tom Tool�bar	��PA?SSWORDy?FRS:\L��� %Passw�ord Config���֏e�Ϗ� B0���T�f������ ����O��s������ >�͟b��[���'��� K��򯁯���:�L� ۯp�����#�5�ʿY� �}��$ϳ�H�׿l� ~�Ϣ�1�����g��� �� ߯���V���z�	� s߰�?���c���
�� .��R�d��߈��� ;�M���q������<� ��`������%���I� �������8���� n���!��W� {"�F�j| �/�Se�� /�/T/�x//�/ �/=/�/a/�/?�/,? �/P?�/�/�??�?9? �?�?o?O�?(O:O�? ^O�?�O�O#O�OGO�O kO}O_�O6_�O/_l_ �O�__�_�_U_�_y_ o o�_Do�_ho�_	o �o-o�oQo�o�o�o �o@R�ov�� ;�_���*�� N��G������7�̏ ޏm����&�8�Ǐ\� 돀��!���E�ڟi� ӟ���4�ßX�j��� �����įS��w��𛯭�B�#��$FI�LE_DGBCK� 1=��/���� (� �)
SUMM?ARY.DGL���OMD:������Diag Su�mmary��Ϊ
CONSLOG��������D�ӱCo�nsole lo�gE�ͫ��MEMCHECK:�!ϯ����X�Memor?y Data��ѧ߁{)��HADOW�ϣϵ�J����Shadow ChangesM��'�-��)	F�TP7Ϥ�3ߨ����Z�mment T�BD��ѧ0=4)�ETHERNE�T�������T�ӱ�Ethernet� \�figura�tionU�ؠ��DCSVRF�߽߫������%�� v�erify alyl��'�1PY���DIFF�����[����%��dif!f]������1R�9�K��� ���{X��CHGD������c��r���2ZAS� 1��GD����k��z��F�Y3bI[� 1�/"GD����s/����/*&�UPDATES.�� �/��FRS:�\�/�-ԱUpd�ates Lis�t�/��PSRBW�LD.CM(?����"<?�/Y�PS_R?OBOWEL��̯ �?�?��?&�O-O�? QO�?uOOnO�O:O�O ^O�O_�O)_�OM___ �O�__�_�_H_�_l_ o�_�_7o�_[o�_lo �o o�oDo�o�ozo �o3E�oi�o� ��R�v��� A��e�w����*��� я`���������O� ޏs������8�͟\� ����'���K�]�� �����4���ۯj��� ���5�įY��}��� ���B�׿�x�Ϝ� 1���*�g�����Ϝ� ��P���t�	�ߪ�?� ��c�u�ߙ�(߽�L� ���߂���(�M��� q� ���6���Z��� ���%���I���B�� ���2�����h����$FILE_� {PR� ��������MDONLY 1�=.�� 
 ���q������� ���~%�I� m�2��h ��!/�./W/�{/ 
/�/�/@/�/d/�/? �//?�/S?e?�/�?? �?<?�?�?r?O�?+O =O�?aO�?�O�O&O�O JO�O�O�O_�O9_�O�F_o_
VISBC�KL6[*.V�Dv_�_.PFR:�\�_�^.PVi�sion VD file�_�O4oFo \_joT_�oo�o�oSo �owo�oB�of �o�+���� ���+�P��t�� ����9�Ώ]�򏁏�� (���L�^������� 5���ܟk� ���$�6� şZ��~�����
�MR_GRP 1�>.L��C4�  B���	 �W�����*u����RHB� ��2 ���� ��� ��� B�����Z�l���C����D�������Ŀ��K���/J�G4I����TX�;F�5UPlf0����ֿ Fl�G��E(	!�;�':t=E�@���@�߶@��ef1�@���@�n�*�E�� F�@ �������J���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6\b��+�&�(�a�hL߅�p�A��A��� ��v���r������
� C�.�@�y�d����� ����������?�Z�,lϖ�BH��8���Ж�������
0�PS?@�P�X��ܿ�� �B���/ ��@'�33:��.�g.N�UUU�U��q	�>u.�?! rX��	�-�=[z�=�̽�=V6<�=��=�=$q������@8�i�7G��8�D��8@9!�7��:����D��@ D�� CϬ���C������' /0-��P/����/N� �/r��/���/�?? ;?&?_?J?\?�?�?�? �?�?�?O�?O7O"O [OFOOjO�O�O�O�O �гߵ��O$_�OH_3_ l_W_�_{_�_�_�_�_ �_o�_2ooVohoSo �owo�o�i��o�o�o ��);�o_J� j������� %��5�[�F��j��� ��Ǐ���֏�!�� E�0�i�{�B/��f/�/ �/�/���/��/A�\� e�P���t�������� ί��+��O�:�s� ^�p�����Ϳ���ܿ � ��OH��o�
ϓ� ~ϷϢ���������� 5� �Y�D�}�hߍ߳� ���������o�1�C� U�y��߉����� ��������-��Q�<� u�`������������� ��;&_J\ ���������� ڟ�F�j4��� ������!// 1/W/B/{/f/�/�/�/ �/�/�/�/??A?,? e?,φ?P�q?�?�?�? �?O�?+OOOO:OLO �OpO�O�O�O�O�O�O _'__K_�o_�_�_ �_l��_0_�_�_�_#o 
oGo.okoVoho�o�o �o�o�o�o�oC .gR�v��� ��	���<�`� *<��`����� ޏ��)��M�8�q�\� ������˟���ڟ� ��7�"�[�F�X���|� ��|?֯�?�����3� �W�B�{�f�����ÿ ���������A�,� e�P�uϛ�b_������ �_��߀�=�(�a�s� Zߗ�~߻ߦ������� � �9�$�]�H��l� ������������#� �G�Y� �B������� z�������
ԏ:�C .gRd���� ��	�?*c N�r����� /̯&/�M/�q/\/ �/�/�/�/�/�/�/? �/7?"?4?m?X?�?|? �?�?�?�?��O!O3O ��WOiO�?�OxO�O�O �O�O�O_�O/__S_ >_P_�_t_�_�_�_�_ �_�_o+ooOo:oso ^o�o�op��o��  ��$��o�o� ~������� 5� �Y�D�}�h����� ��׏����
�C� .�/v�<���8����� �П����?�*�c� N���r��������̯ ��)��?9�_�q��� JO�����ݿȿ�� %�7��[�F��jϣ� ���ϲ�������!�� E�0�i�T�yߟߊ��� ���߮o�o��o>� t�>��b������ �����+��O�:�L� ��p������������� 'K6oZ� Z�|�~����� 5 YDi�z� �����/
// U/@/y/@��/�/�/�/ ���/^/???Q?8? u?\?�?�?�?�?�?�? �?OO;O&O8OqO\O �O�O�O�O�O�O�O_��O7_��$FNO ���VQ��
F�0fQ kP FLA�G8�(LRRM_�CHKTYP  �WP��^P��WP�{QOM�P_MsIN�P����P��  XNPSS�B_CFG ?�VU ���_���S ooIUT�P_DEF_OW�  ��R&hI�RCOM�P8o�$�GENOVRD_�DO�V�6�flT[HR�V d�edkdo_ENBWo k`�RAVC_GRP� 1@�WCa X "_�o_1U< y�r����� 	��-��=�c�J��� n��������ȏ�� ��;�"�_�F�X���ib�ROU�`FVX�P��&�<b&�8�?��埘��������  D�?�јs���@@g�B��7�p�)�ԙ���`S+MT�cG�mM����� �LQHOSTC��R1H���P�\�at�SM��f��\���	12�7.0��1��  e��ٿ����� ǿ@�R�d�vϙ�0�*��	anonymous����������֣�[�� � � ����r����ߨߺ��� ��-���&�8�[�I� �π������ 1�C��W�y���`�r� �����ߺ������� %�c�u�J\n�� �������M�" 4FX��i��� ���7//0/B/ T/���m/��/ �/�/??,?�/P?b? t?�?�/�?��?�?�? OOe/w/�/�/�?�O �/�O�O�O�O�O=?_ $_6_H_kOY_�?�_�_ �_�_�_'O9OKO]O__ Do�Ohozo�o�o�o�O �o�o�o
?o}_R dv���_�_oo !�Uo*�<�N�`�r� �o������̏ޏ�?�Q&�8�J�\���>�E�NT 1I�� sP!􏪟  ����՟ğ������� A��M�(�v���^��� ��㯦��ʯ+�� � a�$���H���l�Ϳ�� ���ƿ'��K��o� 2�hϥϔ��ό��ϰ� ������F�k�.ߏ� R߳�v��ߚ��߾����1���U��y�<�QUICC0��b�t����1�����%����2&���u�!ROUTERv�R�d����!PCJOG�����!192�.168.0.1�0��w�NAME �!��!ROB�OTp�S_CF�G 1H�� ��Auto�-started^�tFTP�� ����� 2 D��hz���� U��
//./�v� ��/���/�/�/ �/�/�!?3?E?W?i? �/?�?�?�?�?�?�? ���AO�?eO�/�O �O�O�O�?�O�O__ +_NO�OJ_s_�_�_�_ �_
OO.OoB_'ovO Ko]ooo�oP_>o�o�o �o�oo�o5GY k}�_�_�_�� 8o��1�C�U�$y� �������ӏf���	� �-�?�����Ə ���ϟ����� ;�M�_�q���.�(��� ˯ݯ��P�b�t��� ��m���������ǿٿ �����!�3�E�h�� {ύϟϱ����$�6� H�J�/�~�S�e�w߉� ��jϿ��������*߀��=�O�a�s��YT_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������OYC�R.RDzVTA{��OGBOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G_BUFF 1X�]	��2	աϸ��� ���������!�N� E�W߄�{ߍߺ߱��� �������J����DCS Zr� =����^�+�ZE��������a�IO ;1[
{ ُ!�� �!�1�C�U�i�y� ��������������	 -AQcu��Ы����EfPTM  �d�2/A Sew����� ��//+/=/O/a/�s/�/�/��SEVt����TYP��/??y͒�R�S@"��×�FL 31\
������?��?�?�?�?�?�?/?T�P6��">�NGNAM�ե�U`�7UPS��GI}�����mA_LOAD��G %�%DF_MOTN����O�@MAXUALRM<��J��@sA�QD����WS ��@C �]m�-_���MP2�7�]^
{ ر�	�!+P�+ʠ�;_/�ƅRr�W�_�WU �W�_��R	o�_o?o "ocoNoso�o�o�o�o �o�o�o�o;&K q\�x���� ���#�I�4�m�P� ��|���Ǐ���֏�� !��E�(�i�T�f��� ��ß��ӟ���� � A�,�>�w�Z������� ѯ����د���O� 2�s�^�������Ϳ����ܿ�'��BD_L?DXDISAX@	���MEMO_AP�R@E ?�+
 � *�~ϐϢϴ�����������@ISCw 1_�+ �� IߨT��Q�c�Ϝ߇� �ߧ�����w����>� )�b�t�[����{� ���������:���I� [�/������������ o�����6!ZlS ��s��� �2�AS'�w ����g��./�/R/d/�_MST�R `�-w%SC/D 1am͠L/�/ H/�/�/?�/2??/? h?S?�?w?�?�?�?�? �?
O�?.OORO=OvO aO�O�O�O�O�O�O�O __<_'_L_r_]_�_ �_�_�_�_�_o�_�_ 8o#o\oGo�oko�o�o �o�o�o�o�o"F 1jUg���� �����B�-�f��Q���u�����ҏh/MKCFG b�-�㏕"LTARMu_��cL��� σQ�N�<�M�ETPUI�ǂ����)NDSP_CMNTh���|� ' d�.��ς��ҟܔ|�POSCF�����PSTOL� 1e'�4@�<#�
5�́5�E�S� 1�S�U�g�������߯ ��ӯ���	�K�-�?����c�u�����|�SI�NG_CHK  y��;�ODAQ,��f��Ç��DEV� 	L�	MC}:!�HSIZEh���-��TASK �%6�%$123456789 ������TRIG 1]g�+ l6�%܀��ǃ�����8�p�Y�P[� ��EM_I�NF 1h3�� `)AT&FV0E0"����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ������H�����A���AI�q�,��|����� ���ߵ��� ��J���n������W� ����������"���� X��/����e�� ����0�T; x�=�as�� /�,/c=/b/�/ A/�/�/�/�/��? ���^?p?#/�?�/ �?s?}/�?�?O�?6O HO�/lO?1?C?U?�O y?�O�O3O _�?D_�O�U_z_a_�_�ONIwTOR��G ?5��   	EX�EC1Ƀ�R2�X3��X4�X5�X���V7*�X8�X9Ƀ�RhB Ld�RLd�RLd�RLd
b LdbLd"bLd.bLd:b�LdFbLc2Sh2_h2�kh2wh2�h2�h2��h2�h2�h2�h3�Sh3_h3�R�R_�GRP_SV 1�in���(����C�?BPP�A4��>%��gY��>r��x�_�D=R^��PL_N�AME !6���p�!Defa�ult Pers�onality �(from FD�) �RR2eq �1j)TUX)TsX��q��X dϏ 8�J�\�n��������� ȏڏ����"�4�F�@X�j�|������2'� П�����*�<�N�`�r��<�������� ү�����,�>�P�tb� �Rdr 1o�y� �\�, ��3���� @D��  ��?�����?x䰺��A'�6�����;�	lʲ	� �xJ������ �< ��"�� �(pK��K ��K=�*�J���J���JV���Zό����rτ́p@j�@T;f��f��ұ]�l��I���������������b��3��´  ��`��>����bϸ�z���Ꜧ���3Jm��
� B�H��˱]���q�	� ~p�  P�p�Q�p��p|  �Ъ�g���c�	'�� � ��I�� �  ��ނ�:�È
�È�=���"�nÿ�	��ВI  �n @B�cΤ�\���B���q�y�o�N���  '������@2��@���X��/�C��C�C�@ C����=��
�A��* #  @<�UP�R�
h�B�"b�A��j�����������Dz۩��߹������j��( �� -���C���'�7�������Y����� �?�ff ��gy> �����o�:a��
>+�  	PƱj�(�����7	���|�?�嚧�xZ�p<
6�b<߈;܍��<�ê<� <�&Jσ��AI�ɳ+���?f7ff?I�?&�k��@�.��J<?�`�q�.� ˴fɺ�/��5/��� �j/U/�/y/�/�/�/��/�/?�/0?q��F�?l??�?/�?�+)�?�?�E�� �E�I�G+� F��?)O�?9O_OJO��OnO�Of�BL޳B �?_h�.��O�O��%_ �OL_�?m_�?�__�_��_�_�_�
�h��<�g>��_Co��_goRodo�o�GA��ds�q�C�o�o�o|����$]H�q���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?�$��?�K/�±�
=ç>�����3�W
=�#��W��e�צ�@�����{�����<��(��B�u���=B0�������	L��H�F��G���G���H�U`E����C�+���I�#�I��H�D�F��E���RC�j=��
�I��@H��!H�( E<YD0q�$� �H�3�l�W���{��� �����՟���2�� V�A�z���w�����ԯ ��������R�=� v�a������������ ߿��<�'�`�Kτ� oρϺϥ�������� &��J�\�G߀�kߤ� ���߳�������"�� F�1�j�U��y���� ���������0��T��?�Q����(��ٙ3/E����u�������M3��8�����M4Mgqs&IB+2�D�a���{�^^	�������uP2P7Q 4_A��M0bt��R������/   �/�b/ P/�/t/�/ *a)_3/�/�/�%1a?�/�?;?M?_?q?   �?�/�?�?�?�?O �2 F�$�vGb�/�A��@�a�`�qC��C@�o�Ot����KF� Dz�H@�� F�P �D���O�O�ys�<O!_3_E_W_i_s?_���@@pZ�4�22!2~
 p_�_�_�_ 	oo-o?oQocouo�o��o�o�o��Q ���+��1��$M�SKCFMAP � �5�� �6�Q�Q"~�cONREL  
�q3�bEXC/FENB?w
s1u�XqFNC_QtJO�GOVLIM?wdtIpMrd�bKEY?wu�u�bRUN�|��u�bSFSP�DTY�avJu3sS�IGN?QtT1M�OT�Nq�b_C�E_GRP 1p�5s\r���j� ����T��⏙���� ��<��`��U���M� ��̟��🧟�&�ݟ J��C���7������� گ�������4�V�`�TCOM_CFG 1q}�Vp������
P�_ARC_�\r
jyUAP_�CPL��ntNOCHECK ?{ 	r�� 1�C�U�g�yϋϝϯπ��������	��({N�O_WAIT_L��	uM�NTX�r�{�[m�_ERR�Y�2sy3�  &�������r�c� ��T_MO��t>��, 62$�k�3�PARAM��u{�	�[����u?�� =9@345?678901�� &���E�W�3�c�����`{�������������=�UM_RSPACE �Vv���$ODRDS�P���jxOFFSET_CARTܿαDIS��PE?N_FILE� �q���c֮�OPTIO�N_IO��PW�ORK v_��ms �P(�R��@�6$j.j	 ���Hj(6$�p=�_DSBL  �5�Js�\��RIE�NTTO>p9!CᴧPqfA� UT__SIM_D
r��b� V� LCT ww�bc��U)+$�_PEXE�d&R�ATp �vju�p��2�X�j)TUX)T�X�##X d -�/�/�/??1?C? U?g?y?�?�?�?�?�?��?�?	OO-O?O�H2 �/oO�O�O�O�O�O�O�O�O_]�<^O;_M_ __q_�_�_�_�_�_�_`�_o���X�OU[��o(��(����$o�, ���IpB` @D��  Ua?�[cAa?p]a]�DWcUa쪞�l;�	lmb�`�xJ�`�p���a�</ ��`�m�a���H(��H3k�7HSM5G�2�2G���Gp
1��
���'|���CR�>�>q��GsuaT�3���  �4spBpyr  �]o�*SB_�����j]��t�q� ��rna� �,���6  ���PQ�
|N�M�,k���	'� � ���I� �  ���%�=���Э���ba	���I�  �n @@��~���p��������N	 W�  '�!o�:q�pC	 C�A@@sBq�|��� m��
�!�h@ߐ"�n����*�B	 �qA���p� �-�qbz��P��t�_�������( ?�� -��� ��n�ڥ[A]Ѻ�b4��'!5�(p �?��ff� ��
����OZ�R*�85�z����>΁  Pia��( 5���@���ک�a�c�d^F#?��5�x���*�<
6b<���;܍�<����<� <�&�o&�)�A�lcΐ|I�*�?fff?��?&c���@�.�uJ<?�` ��Yђ^�nd��]e�� [g��Gǡd<����1� �U�@�y�dߝ߯ߚ� ���߼�	���-�������&��"�E�� �E��G+� Fþ�����������@&��J�5��bB��AT�8�ђ��0�6��� >���J�n�7��[�m�0��h��<1��>�M��I
�@��A�[��C-�)��?���� /�YĒ��Jp��vaFv`CH/�������}!@I�Y�'��3A�A�AR�1AO�^?��$�?�������
=ç>�����3�W
=�s#����+e��ܒ������{�����<��.(��B�u���=B0�������	�*H�F��G���G���H�U`E����C�+�-I�#�I��H�D�F��E���RC�j=U>
�I��@H��!H�( E<YD0/�?�? �?�?�?O�?3OOWO BOTO�OxO�O�O�O�O �O�O_/__S_>_w_ b_�_�_�_�_�_�_�_ oo=o(oaoLo�o�o �o�o�o�o�o�o' $]H�l�� �����#��G� 2�k�V���z���ŏ�� �ԏ���1��U�g� R���v�����ӟ��������-��(��ٙ�����a�����Q�c�,!3��8�}���,!4Mgqs����ɢIB+կ�篴a���{���A�/�e�S����w��P!�P���� ���7��ӯ�ϑ�R9�Kτ�oχϓ���  ���χ�� ��)��M������z���{߉ߛ���ߒ���������   )�G�q�_����2 F�$�&Gb���n�[ZjM!C�s�@j/�A��S�=�F� Dz���� F�P �D��W����)������������x?_���@@
9�=�=��=��
 v�� �����*�<N`�*P ����˨�1��$P�ARAM_MEN�U ?-���  �DEFPULSE�l	WAITT�MOUT�RC�V� SHE�LL_WRK.$�CUR_STYLv�,OPT�N/PTB./("C�R_DECSN� ��,y/�/�/�/�/�/ �/?	??-?V?Q?c?�u?�?�USE_P�ROG %�%��?�?�3CCR������7_HOST7 !�!�44O��:T̰�?PCO)A�RC�O�;_TIME��XB�  �GDEBUGV@��3�GINP_FLMSK�O�IT`��O�EWPGAP �L���#[CH�O�HTYPE����?�?�_ �_�_�_�_oo'o9o bo]ooo�o�o�o�o�o �o�o�o:5GY �}����������1�Z��EWO�RD ?	7]	�RS`�	PNeS�$��JOE!�>�TEs@WVTR�ACECTL 1�x-�� ��� ������ɆDT Qy�-���D �{ ���4�P :�L :�GP :�D :�@ :�8�,� >�P�b�����П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�V�(�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_d��_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п�_ ���*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ //�$)�$PGTRA�CELEN  �#!  ���" �8&_UP z���g!�o S!h 8!_�CFG {g%Q#"!x!�$J �#�|"DEFSPD �|�,!!J ��8 IN TRL +}�-" 8�%�!�PE_CONFI�� ~g%��g!�$�%�$LID�#�-74GRP� 1�7Q!��#!A ���&f�f"!A+33D��� D]� C�O� A@+6�!�" �d�$�9�9*1*0� 	 +9�(�&�"��? ´	C�?�;B @3AO�?OIO3OmO�"!>�T?�
�5�O�O�N�O =?��=#�
�O_ �O_J_5_n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_ Roxoco�o�o�o�o�o �o�o>)bM���;
V7.1�0beta1�$�  A�E>�rӻ�A " �p�?!G��q>�嚻r��0�q��޻qBQ��qA\��p�q�4�q�p�"�BȔ2�D�V�h�w�!�p�?�?)2{ȏ w�׏���4��1� j�U���y�����֟�� ����0��T�?�x� c�������ү����!o �,�ۯP�;�M���q� ����ο���ݿ�(π�L�7�p�+9��sF@ �ɣͷϥ�g% ������+�!6I�[� �������ߵߠ����� ����!��E�0�B�{� f����������� ��A�,�e�P���t� ����������� =(aL^��� ����'9$ ]�Ϛ��ϖ����� ��/<�5/`�r߄� �ߏ/>�/�/�/�/�/ ?�/1??U?@?R?�? v?�?�?�?�?�?�?O -OOQO<OuO`O�O�O �O�O���O_�O)__ M_8_q_\_n_�_�_�_ �_�_�_o�_7oIot ���o�o���o�o �o(/!L/^/p/�/{ *o������� ��A�,�e�P�b��� �������Ώ��+� =�(�a�L���p����� �Oߟ񟠟� �9�$� ]�H���l�~�����ۯ Ư���#�No`oro�o n��o�o�o�oԿ�� �8J\ng���� vϯϚ�������	��� -��Q�<�u�`�r߫� ���ߺ�������;� M�8�q�\�������� z������%��I�4� m�X���|��������� ��:�L�^���Z�� ���������$� 6�H�Swb� ������// =/(/a/L/�/p/�/�/ �/�/�/?�/'??K? ]?H?�?��?�?f?�? �?�?O�?5O OYODO }OhO�O�O�O�O�O�O &8J4_F_��� �_�_��_�_"4 -o�O*ocoNo�oro�o �o�o�o�o�o) M8q\���� �����7�"�[� m��?����R�Ǐ��� ֏�!��E�0�i�T� ��x��������_$_ V_ �2�l_~_�_������R�$PLID_�KNOW_M  ��T�|����SV ��U�͠�U ��
��.�ǟR�=�O������mӣM_GROP 1��!`0u���T@ٰo�ҵ�
���Pзj��` ���!�J�_�W�i�{� �ϟϱ����������V��MR�����T��s�w� s��ߠ޴� �߅��ߩ߻�����A� ��'������ ��������=��� #���������}�������S��ST��1 1Ն�U# ���0�_ A .��,> Pb������ ��3(iL^�p�����2r*���<-/�3/)/;/M/4 f/x/�/�/5�/�/�/�/6??(?:?�7S?e?w?�?8�?�?�?�?MAD  d#`�PARNUM  �w�%OSCH?J ME
�G`A�Iͣ�EUPD`OrE
a��OT_CMP_0��B@�P@'˥T�ER_CHK'U���˪?R$_6[RS8l�¯��_MOA@�_�U_�_RE_RES_G ��>�o o8o+o\oOo�oso�o �o�o�o�o�o�o�W �\�_%�Ue B af�S� ����S 0����SR0�� #��S�0>�]�b��S�0�}������RV 1�x����rB@c]��}t�(@c\��}��D@c[�$����RTHR_IN�Rl�DA��˥d,�M�ASS9� ZM�M�N8�k�MON_QUEUE ���X˦��x� RDNP�UbQN{�P[��ENqD���_ڙEXE韌ڕ�@BE�ʟ��O�PTIOǗ�[��P�ROGRAM %��%��ۏ�O��?TASK_IAD0�OCFG ���xtO��ŠDATA��]�Ϋ@��27� >�P�b�t���,����� ɿۿ�����#�5�G�^��INFOUӌ�������ϭϿ����� ����+�=�O�a�s� �ߗߩ߻��������4^�jč� yġ~?PDIT �ί|c���WERFL
���
RGADJ ��n�A����?�����@���IORI�TY{�QV���MPGDSPH�����Uz�y���OTOEy��1�R� (!�AF4�E�P]����!tcph����!ud��!�icm��ݏ6�XYm_ȡ�R��ۡ)� *+/ ۠�W:F�j ������%@7[B�*��OPORT#�BC۠�����_CAR�TREP
�R� S�KSTAz��ZSS�AV���n�	2500H863��P�r�$!�R����q�n�}/�/�'^� URGE�B��6rYWF� DO{�r�UVWV��$�A�WR�UP_DELAY� �R��$R_HOTk��%O]?�$�R_NORMAL�k�L?�?p6SEMI�?�?�?3AQSKI�P!�n�l#x 	1/+O+ OROdO vO9Hn��O�G�O�O�O �O�O_�O_D_V_h_ ._�_z_�_�_�_�_�_ 
o�_.o@oRoovodo �o�o�o�o�o�o�o *<Lr`����n��$RCVT�M�����pDC�R!�LЈqB���C*J�C�$�>�$ >5>�;��04M�¹�O��ǃ��������~���9On�Y�<
6b�<߈;܍��>u.�?!<�&{�b�ˏݏ ��8�����,�>�P� b�t���������Ο�� �ݟ��:�%�7�p� S������ʯܯ� � �$�6�H�Z�l�~��� ����ƿ���տ��� 2�D�'�h�zϽ��ϰ� ��������
��.�@� R�d�Oψߚ߅߾ߩ� ��������<�N�� r����������� ��&�8�#�\�G��� ��}����������� S�4FXj|�� �������0 T?x�u�� ��'//,/>/P/ b/t/�/�/�/�/�/�/ �?�/(??L?7?p? �?e?�?�?��?�? O O$O6OHOZOlO~O�O �O�?�?�O�O�O�O _ _D_V_9_z_�_�?�_ �_�_�_�_
oo.o@o�Rodovo�X�qGN_�ATC 1��� AT&F�V0E/� A�TDP/6/9/�2/9�hATA��n,AT%G1%B960/�_+++�o,�a�H,�qIO_T?YPE  �u�s�n_�oREFPO�S1 1�P{ 'x�o�Xh_� d_�����K�6� o�
���.���R����^{{2 1�P{����؏V�ԏz����q3 1��$�6�p���ٟ���S4 1� ����˟���n���%�S5 1�<�N�`������<���S6 1�ѯ���/�����|ѿO�S7 1�f��x���ĿB�-�f��S8 1�����Y��������y�SMAS�K 1�P  
89�G��XNOM����a~߈ӁqMOT�E  h�~t��_CFG ���������rPL_RANG��ћQ��POWER� ��e��S�M_DRYPRG %i�%��J��TART �
��X�UME_PRO�'�9��~t_EXE�C_ENB  <�e��GSPD����8��c��TDB���sRM��MT_!��T���`OBO�T_NAME �i���iOB_�ORD_NUM �?
�\qH863  �T���������bPC�_TIMEOUT��� x�`S232���1��k L�TEACH PENDAN �ǅ��}���`Ma�intenanc?e Cons�R}��m
"{�dKCLC/Cg��Z ��n�� No U�se}�	��*N�PO��х�z��(CH_L��3�����	�m?MAVAIL���{��ՙ�SPAC�E1 2��| d��(>��&����p��M,8�?�ep/eT/�/�/ �/�/�W//,/>/�/ b/�/v?�?Z?�/�?�9 �e�a�=??,?>?�? b?�?vO�OZO�?�O�O(�Os�2�/O *O<O�O`O�O�_�_u_ �_�_�_�_[3_#_ 5_G_Y_o}_�_�o�o@�o�o�o[4.o @oRodovo$�o�o�����"�	�7�[5 K]o��A��� �	�̏�?�&�T�[6h�z�������^�ԏ ���&��;�\�C�q�[7��������͟{� ��"�C��X�y�`���[8����Ưد� ���0�?�`�#�uϖ�x}ϫ�[G �iۧ �ϋ
G� ����$�6�H�Z� l�~ߐ��8 ǳ�����߈��d(��� M�_�q������ �����?���2�%�7� e�w������������� �������!�RE�W� ����������?Q `�� @0��ߖrz	�V_�� ���
/L/^/|/2/ d/�/�/�/�/�/�/? �/�/�/*?l?~?�?R? �?�?�?�?�?�?�?2O��?
��O[_M?ODE  �˝I/S ���vO,�*ϲ�O-_��	�M_v_#dCWORK�_AD�Mxq�^%aR  ��ϰ��P{_�P_INTV�AL�@����JR_�OPTION�V ��EBpVAT_�GRP 2���;�(y_Ho �e_vo�o�oYo�o �o�o�o�o*<� bOoNDpw��� ���	���?�Q� c�u�����/���Ϗ� �����)�;���_�q� ��������O�ɟ�� �՟7�I�[�m�/��� ����ǯٯ믁��!� 3���C�i�{���O��� ÿտ���ϡ�/�A� S�e�'ωϛϭ�oρ� ������+�=���a� s߅�Gߕ߻����ߡ� ��'�9�K�]��߁� ����y�����������5�G�Y��E�$SCAN_TIM�A�Yuew�R ��(�#((�<0�.aaPaP
Tq>��Q���o�����OO2/��:	�d/JaR��WY ��^���^R^	r�  P���; �  8�P�x	�D�� GYk}���������Qp�/@/R//)P;G�o\T��Qpg-��t�_Di�KT��[  � l v%������/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OWW�#�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_olO~Od+No `oro�o�o�o�o�o�o �o&8J\n�������u�  0�"0g�/�-�?� Q�c�u���������Ϗ ����)�;�M�_� q�����$o��˟ݟ� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�����Do���� ����ҿ�����,� >�P�b�tφϘϪϼ����������w
�   58�J�\�n߀ߒߜ� ����������	��-� ?�Q�c�u����� ��-�����  �2�D�V�h�z��������������������& ��%	�1234567�8�" 	��/� `r��������( :L^p���� ��� //$/6/H/ Z/l/~/��/�/�/�/ �/�/? ?2?D?V?h? �/�?�?�?�?�?�?�? 
OO.O@Oo?dOvO�O �O�O�O�O�O�O__ *_YON_`_r_�_�_�_ �_�_�_�_ooC_8o Jo\ono�o�o�o�o�o �o�oo"4FX j|���������	��s3�E��W�{�Cz  B}p��   ���2���z�$SCR�_GRP 1�(��U8(�\x�^ @}  	�!�	 ׃���"�$� Հ�-��+��R�w����D~������#����O���M�-10iA 89�09905 Ŗ5 M61C >4��TJׁ
� ��� 0�����#�1�	"�z�������¯Ҭ ���c�� �O�8�J��������!�����ֿ��B��y���������A��$�  @��<� �"R�?��d���Hy�u��O���F@ F�`�§�ʿ�϶����� ��%��I�4�m��<��l߃ߕߧ߹�B� ��\����1��U�@� R��v�������� ������;���*<=��
F���?�d�<�>73�����@�:���7 B���ЗЙ����EL_DEFAULT  �����B��MIPOWERFL  �$�1 WFDO �$��ERVENT? 1�����"��pL!DUM�_EIP��8��j�!AF_INEx �=�!FT����!��4 ���[!RP?C_MAIN\>q�J�nVISw�=���!TP&�PU��	d�?/�!
PMON_POROXY@/�e./��/"Y/�fz/�/!�RDM_SRV��/�	g�/#?!R� C?�h?o?!
�pM�/�i^?�?!RLSYNC�?�8�8�?O!R3OS�.L�4�?SO "wO�#DOVO�O�O�O �O�O_�O1_�OU__ ._@_�_d_v_�_�_�_��_o�_?oocoiI�CE_KL ?%�y (%SVCPRG1ho8��e����o�m3�o�o�`4� �`5(-�`6PU�`7x}�`�$��l9��{�d:? ��a�o��a�oE��a �om��a���aB�� �aj叟a���a� 5��a�]��a����a 3����a[�՟�a���� �a��%��aӏM��a�� u��a#����aK�ů�a s���a��mob�`�o �`8�}�w�������ɿ ���ؿ���5�G�2� k�VϏ�zϳϞ����� �����1��U�@�y� dߝ߯ߚ��߾����� ��?�*�Q�u�`�� ����������� ;�&�_�J���n�����������sj_DE�V y	��MC:��_.OUT",~REC 1�Z�� d    ]	�     ��@�������A����
� �PSD#6S r��O� �� %�� `�� �Z�{*� �� *��  +X- � I�- �- !- � ��X�YZ�PSJ;�4 �? Z (�  � ԣ�R ��� E- � �/e/�l4�/�R�� X� (,/�>/P/�/�/�""4�R =�!� � ؀ � ?"S1��'!V�/���("- �� \?�?$=�=�?�?�?"O OFO4OjO|O^O�O�O �O�O�O�O�O_ __ T_B_x_f_�_�_�_�_ �_�_�_oooPo>o to�oho�o�o�o�o�o �o(
L:\� p���w,� ���4�"�X�F�|� ��p�����֏ď�� ��0��@�f�T���x� ����ҟ�Ɵ���,� �<�b�P���h�z��� ���ί��(�:�� ^�L�n�p�������ܿ �п� �6�$�Z�H� jϐ�rϴϢ������� ���2�D�&�h�Vߌ� z߰ߞ����������� 
�@�.�d�R��ZjoV 1�w P������ 
�� ����
TY�PEVFZN_�CFG ��5�d�4�GR�P 1�A�c �,B� A� D;� B���  �B4RB2�1HELL:�(
��?���<%RS'!��H 3lW�{��� ���2VhV������%w ����#!�1�L����7�2�0�d����HK 1��� �k/f/ x/�/�/�/�/�/�/�/ ??C?>?P?b?�?�?��?�?��OMM ���?��FTOV�_ENB ���+�H�OW_REG_U�IO��IMWAI�TB�JKOUTr;F��LITIM;Ew���OVAL[O>MC_UNITC�F�+�MON_ALI�AS ?e�9 ( he��_&_8_ J_\_B_�_�_�_�_ j_�_�_oo+o�_Oo aoso�o�oBo�o�o�o �o�o'9K] n����t�� �#�5��Y�k�}��� ��L�ŏ׏������ 1�C�U�g�������� ��ӟ~���	��-�?� �c�u�������V�ϯ ������;�M�_� q��������˿ݿ�� ��%�7�I���m�� �ϣϵ�`�������� ��3�E�W�i�{�&ߟ� �������ߒ���/� A�S���w����X� ����������=�O� a�s���0��������� ����'9K] ����b��� #�GYk}� :������/ 1/C/U/ /f/�/�/�/ �/l/�/�/	??-?�/ Q?c?u?�?�?D?�?�? �?�?O�?)O;OMO_O 
O�O�O�O�O�OvO�O�__%_7_�C�$S�MON_DEFP�RO ����`Q �*SYSTEM�*  d=OUR�ECALL ?}�`Y ( �}
�xyzrate �61 *.* v�irt:\tmp�back\�P=>�192.168.�4�P46:224�4 �Q�_�_�_�K}��W�^5288 ��_�_couo�ob9c�opy frs:�orderfil.dat�\*o<a�o��o�ol0�bmdb:�_�o<a�obt�rc6�o�hemp:1660 W��:�.�v*.d��~ �`�r���e�Y+�=� O�����o)o҂�� ҏc�u����o�o5�w ٟ���"���xџ�b�t����4x��: �Q�_;�M�V�����}5��a����7�ׯ h�z������:�կ� ��
����A�ӿd�v� �ϛ�.�;�ѯ����� ��ϼ�O�`�r߄ߗ� ��2�Ϳ������'� ��K�\�n��ϥ�8� ���������#ߴ�G� �j�|����_3�E�W�������� �Hf472 ����bt��8�߲�*< ����/ �3	�as��3���/T� �	/��(��6�f/ x/�/��//A/S/�/�/?�>|54>o�/a? s?�?�ߪ349�?�? �?�"�?58�?bOtO �O��?��85=`WO �O�O�O��O�J�Oa_ s_�_�/��<_N_�_�_ o?(?�S�_�_couo �o�?�?5O�G�o�o�o O"O�o�H�obt� ��/�/QdV������8 �g�y� ���o�o9T���	� ��@ҏc�u�������$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1����?���%֟ ��&�	��\�?�f� ��u��������ϯ�� "��F�)�;�|�_��� ����ֿ��˿��� B�%�f�I�[Ϝ�Ϧ� �ϵ�������,��6� b�E߆�i�{߼ߟ��� ��������L�/�V� ��e��������� ���6��+�l�O�v� �������������� 2V9K�o� ������& R5vYk��� ��/��<//F/ r/U/�/y/�/�/�/�/ ?�/&?	??\???f? �?u?�?�?�?�?�?�? "OOFO)O;O|O_O�O �O�O�O�O�O_�O_ B_%_f_I_[_�__�_ �_�_�_�_�_,oo6o boEo�oio{o�o�o�o �o�o�oL/V �e������ ��6��+�l�O�v��������PARAM� ����� ��	��P�����OFT_K�B_CFG  �⃱���PIN_S_IM  ����C�U�g�����RVQSTP_DSB,��򂣟����SR ��/�� & gCAR������TOP_ON_E�Rސ���P_TN /�@��A	�RIN�G_PRM� ���VDT_GRP� 1�ˉ�  	������������Я �����*�Q�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߣߠ� ������������0� B�i�f�x������ �������/�,�>�P� b�t������������� ��(:L^p �������  $6HZ�~� ������/ / G/D/V/h/z/�/�/�/ �/�/�/?
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O�__&_8___\_��V�PRG_COUN�T��@���RENBU��UM�S��__UPD 1�/�8  
s_�o o*oSoNo`oro�o�o �o�o�o�o�o+& 8Jsn���� �����"�K�F� X�j���������ۏ֏ ���#��0�B�k�f� x���������ҟ���� ��C�>�P�b����� ����ӯί������UYSDEBUG��P�P�)�d�YH�S�P_PASS�U�B?Z�LOG ���U�S)��#�0�  ��Q)�
MC:\��6���_MPC���U�ϒ�Qñ8� �Q�S_AV �����lǲ%�ηSV;��TEM_TIMEw 1��[ (�P�)�T��{�ؿT1S�VGUNS�P�U'��U���ASK_?OPTION�P�U��Q�Q��BCCF�G ��[u� n�X�G�`a�gZo� �߃ߕ��߹������ �:�%�^�p�[��� ������� �����6� !�Z�E�~�i���������%�������&8 ��nY�}�?� �ԫ ��( L:p^���� ���/ /6/$/F/ l/Z/�/~/�/�/�/�/ �/�/�/2?8 F?X? v?�?�??�?�?�?�? �?O*O<O
O`ONO�O rO�O�O�O�O�O_�O &__J_8_n_\_~_�_ �_�_�_�_�_o�_ o "o4ojoXo�oD?�o�o �o�o�oxo.T Bx��j��� �����,�b�P� ��t�����Ώ��ޏ� �(��L�:�p�^��� ����ʟ��o�� 6�H�Z�؟~�l����� ��د���ʯ ��D� 2�h�V�x�z���¿�� �Կ
���.��>�d� Rψ�vϬϚ��Ͼ��� ����*��N��f�x� �ߨߺ�8�������� �8�J�\�*��n�� �����������"�� F�4�j�X���|����� ��������0@ BT�x�d��� ��>,Nt b������/ �(//8/:/L/�/p/ �/�/�/�/�/�/�/$? ?H?6?l?Z?�?~?�? �?�?�?�?O�&O8O VOhOzO�?�O�O�O�O �O�O
__�O@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<o^o�o ro�o�o�o�o�o�o  J8n$O�� ���X���4��"�X�B�v��$TB�CSG_GRP �2�B���  �v� 
 ?�  ������ ׏�������1��U��g�z���ƈ�d�, ���?v�	 �HC��d�>�����e�CL  Bጙ�Пܘ������\)��Y  3A�ܟ$�B�g�B�#Bl�i�X�ɼ���>X��  D	J���r�����C����үܬ���D�@v�=�W� j�}�H�Z���ſ���������v�	�V3.00��	�m61c�	�*X�P�u�g�p�>�d��v�(:�� ���p͟�  O�����p�����z�JCFoG �B���Y ���������=��=�c�q� K�qߗ߂߻ߦ����� ���'��$�]�H�� l������������ #��G�2�k�V���z� ������������ �p*<N���l� ������#5 GY}h��� �v�b��>�// / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?d? R?t?v?�?�?�?�?�? O�?*OO:O`ONO�O rO�O�O��O�O�O_ &__J_8_n_\_�_�_ �_�_�_�_�_�_�_o Fo4ojo|o�o�oZo�o �o�o�o�o�oB0 fT�x���� ���,��P�>�`� b�t�����Ώ����� ��&�L��Od�v��� 2�����ȟʟܟ� � 6�$�Z�l�~���N��� ��دƯ�� �2�� B�h�V���z�����Կ ¿����.��R�@� v�dϚψϪ��Ͼ��� ����<�*�L�N�`� �߄ߺߨ����ߚ�� �����\�J��n�� ���������"��� 2�X�F�|�j������� ��������.T Bxf����� ��>,bP �t�����/ �(//8/:/L/�/�� �/�/�/h/�/�/�/$? ?H?6?l?Z?�?�?�? �?�?�?�?O�?ODO VOhO"O4O�O�O�O�O �O�O
_�O_@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<oro`o �o�o�o�o�o�o�o &�/>P�/�� �������4� F�X��(���|����� ֏����Ə0��@� B�T���x�����ҟ�� ����,��P�>�t� b������������� ��:�(�^�L�n��� ����2d�����̿ �$�Z�H�~�lϢϐ� �������Ϻ� ��0� 2�D�zߌߞ߰�j��� �������
�,�.�@� v�d��������� ����<�*�`�N��� r������������� &J\�t�� B������ F4j|��^����/�  2 6# 6&J/6"��$TBJOP_�GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� ƞ6$ @2 �"	� �C�� �&b�  Cق'�!�!>ǌ��
559>��0+1�33=��CL� fff?>+0?�ffB� J1��%Y?d7�.��/>;��2\)?0��5���;��h{CY� �  @� ~�!B�  A�P?��?�3EC�  D��!�,�0*BO���?�3JB��
:�/��Bl�0��0�$��1�?O6!Aə�3AДC�1D�G6Ǌ=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__<�O�O>B�\JU�O�HH�1ts�A@g33@?1� C�� ��@�_�_&_8_>��D�UV_0�LP�Q30O<{�zR� @�0 �V�P!o3o�_<oRifo Po^o�o�o�oRo�o�o �o�oM(�ol��p~��p4�6&��q5	V3.0}0�#m61c�$�*(��$1!6�A�� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�IR�CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;S@;Q�U�|8�`rz@/&�8�6&<��1��w�^$ESTPAR�S  *({ _#H�R��ABLE 1%�p+Z�6#|�Q�Q � 1�|�|�|��5'=!|�	|�
|��|�˕6!|�|�:|���RDI��z!ʟܟ� ��$���O������¯ԯ�����S��x# V���˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���U-����ĜP�9� K�]�o��-�?�Q�c��u���6�NUM  ��z!� �>  Ȑ����_CF�G �����!@�b IMEBF_T�T����x#��a�VE�R��b�w�a�R {1�p+
 (3�6"1 ��  6!�� �������� �9�$�:� H�Z�l�~���������@������^$��_���@x�
b MI_�CHANm� x� >kDBGLV;0o��x�a!n ETHE�RAD ?�
� �y�$"�\&�n ROUT��!�p*!*�SN�MASK�x#�255.h�fx�^$OOLOFS_�DI��[ՠ	OR�QCTRL � p+;/���/+/=/ O/a/s/�/�/�/�/�/���/�/�/!?��PE?_DETAI���PON_SVOF�F�33P_MON� �H�v�2-9S�TRTCHK ����42VTCOMPATa8�24�:0FPROG =%�%CA)&O~�3ISPLAY���L:_INST_M�P GL7YDUS8���?�2LCK�LPKQUICKMEt ��O�2SCRE�@}�
tps�@�2�A�@�I��@_Y����9�	SR_GR�P 1�� ���\�l_zZg_@�_�_�_�_�_�^�^� oj�Q'ODo/ohoSe ��oo�o�o�o�o�o �o!WE{i�������	1234567�h�!���X�E1�V[�
 �}ipn�l/a�gen.htmno��������ȏ�~�Panel� setup̌}��?��0�B�T�f� ��񏞟��ԟ� ��o����@�R�d�v� �����#�Я���� �*���ϯůr����� ����̿C��g��&� 8�J�\�n�����϶� ��������uϣϙ�F� X�j�|ߎߠ����;� ������0�B��*N�UALRMb@G ?�� [��� ���������� ��%� C�I�z�m�������v�SEV  �����t�ECFG CՁ=]/BaA$�   B�/D
 ��/C�Wi{� ������4 PRց; �To�\o�I�6?K0(%����0���� �//;/&/L/q/\/`�/�/�/l�D ��Q�/I_�@HIS�T 1ׁ9  �(  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1�?v?�?�?�?�� >?P=71c?�?	OOx-O�?�:edit[2CAR�?|O�O�O�O8AO�?]0962kO _�_$_6_�O�O�A36 �O�_�_�_�_IR�_�_ �_oo+o=o�_aoso �o�o�o�oJo�o�o'9I|��a81�o u������o� ��)�;�M��q��� ������ˏZ�l��� %�7�I�[������� ��ǟٟh����!�3� E�W����������ï կ�v���/�A�S� e�Pb������ѿ� �����+�=�O�a�s� ϗϩϻ�������� ��'�9�K�]�o߁�� �߷��������ߎ�#� 5�G�Y�k�}���� �����������1�C� U�g�y���v������� ����	�?Qc u��(���� )�M_q� ��6���// %/�I/[/m//�/�/ �/D/�/�/�/?!?3? �/W?i?{?�?�?�?�� ���?�?OO/OAOD? eOwO�O�O�O�ONO`O �O__+_=_O_�Os_ �_�_�_�_�_\_�_o o'o9oKo�_�_�o�o �o�o�o�ojo�o# 5GY�o}�������?��$UI�_PANEDAT�A 1������  	�}�0�B�T�f�x��� )����mt� ۏ����#�5���Y� @�}���v�����ן�� �����1��U�g�N�\����� �1�� Ïȯگ����"�u� F���X�|�������Ŀ ֿ=������0�T� ;�x�_ϜϮϕ��Ϲ� �����,ߟ�M�� j�o߁ߓߥ߷���� ��`��#�5�G�Y�k� �ߏ���������� ����C�*�g�y�`� ��������F�X�	 -?Qc����߫ ����~; "_F��|�� ���/�7/I/0/ m/�����/�/�/�/�/ �/P/!?3?�W?i?{? �?�?�??�?�?�?O �?/OOSOeOLO�OpO �O�O�O�O�O_z/�/ J?O_a_s_�_�_�_�O �_@?�_oo'o9oKo �_oo�oho�o�o�o�o �o�o�o#
GY@ }d��&_8_�� ��1�C��g��_�� ������ӏ���^�� �?�&�c�u�\����� ��ϟ���ڟ�)�� M�����������˯ ݯ0�����7�I�[� m����������ٿ� ҿ���3�E�,�i�P� �ϟφ��Ϫ���Z�l�}���1�C�U�g�y���)߰�#�������  ��$�6��Z�A�~� e�w��������� ��2��V�h�O������v�p��$UI_P�ANELINK �1�v� � �  ���}1234567890����	 -?G ���o�� ���a��#5G�	����p&���  R��� ��Z��$/6/H/ Z/l/~//�/�/�/�/ �/�/�/
?2?D?V?h? z??$?�?�?�?�?�? 
O�?.O@OROdOvO�O  O�O�O�O�O�O_�O �O<_N_`_r_�_�_�0,���_�X�_�_�_  o2ooVohoKo�ooo �o�o�o�o�o�o� �,>r}����� �������/� A�S�e�w�������� я���tv�z��� �=�O�a�s������� 0S��ӟ���	��-� ��Q�c�u�������:� ϯ����)���M� _�q���������H�ݿ ���%�7�ƿ[�m� ϑϣϵ�D������� �!�3�Eߴ_i�{�
 �߂����߸������ /��S�e�H���~� ��R~'�'�a��:� L�^�p����������� ���� ��6HZ l~���#�5�� � 2D��hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?�/�?�?�?�? �?�?m?OO&O8OJO \O�?�O�O�O�O�O�O �O[�_��4_F_)_j_ |___�_�_�_�_�_�_ o�_0ooTofo��o ��o��o�o�o ,>1bt��� �K����(�:� ���{O������ʏ ܏�uO�$�6�H�Z� l���������Ɵ؟� ���� �2�D�V�h�z� 	�����¯ԯ����� �.�@�R�d�v���� ����п���ϕ�*� <�N�`�rτ��O�Ϻ� Io���������8�J� -�n߀�cߤ߇����� �����o1�oX��o |����������� ��0�B�T�f���� ����������S�e�w� ,>Pbt��' �����: L^p��#�� �� //$/�H/Z/ l/~/�/�/1/�/�/�/ �/? ?�/D?V?h?z? �?�?�???�?�?�?
O O.O��ROdO�߈OkO �O�O�O�O�O�O_�O <_N_1_r_�_g_�_7O�M�m�$UI�_QUICKME�N  ���_AobRESTORE 1��  ��|��Rto�o�im �o�o�o�o�o: L^p�%��� ���o����Z� l�~�����E�Ə؏� ��� �ÏD�V�h�z� ��7�������/���
� �.�@��d�v����� ��O�Я�����ß ͯ7�I���m������� ̿޿����&�8�J� �nπϒϤ϶�a��� ����Y�"�4�F�X�j� ߎߠ߲������ߋ����0�B�T�gSC�RE`?#m�u1sco`uU2��3��4��5��6��7��8��bUGSERq�v��Tp঑�ks����4��5*��6��7��8��`�NDO_CFG ��#k  n` �`PDATE ����Non�ebSEUFRA_ME  �TA��n�RTOL_AB�RTy�l��ENB�����GRP 1��ci/aCz  A�����Q�� $�6HRd��`U������MSK  ������Nv�%��U�%���bVI�SCAND_MA�X�I��FAIL_IMG� ��PݗP#��IM�REGNUM�
�,[SIZ�n`��A�,VONT�MOU��@����2��a���a����F�R:\ � �MC:\�\wLOG�B@F� !�'/!+/O/�U�z MCV��8#UD1r&E�X{+�S�PPO�64_��0'f�n6PO��LI�b�*�#V���,�f@�'�/� =	��(SZV�.�����'WAI�/ST�AT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_�JMPERR 1��#k
  �23�45678901 dF�ψO{O�O�O�O�O �O_�O*__N_A_S_x�_
� MLOWc>8
 �_TI�=��'MPHASOE  ��F��P�SHIFT�15 9�]@<�\� Do�U#oIo�oYoko�o �o�o�o�o�o�o6 lCU�y�� ��� ��	�V�-��e2����	VSwFT1�2	V�M�� �5�1G� ����%A�  BU8̀̀�@ pك�Ӂ˂�у��z�ME�@�?�{��!c>&+%�aM1��k�0��{ �$`0TDI�NEND��\�O � �z����S��w���P���ϜRELE�Q��Y���\�?_ACTIV��<:�R�A ��e���e�:�RD� ���YBOX �9��د�6��02����190.0m.�83���254��QF�	� �X�j��1�robot����   px�૿�5pc�� ̿�����7�����-�^f�ZABC�����,]@U��2ʿ�eϢ� �ϛϭϿ����� �� �V�=�z�a�s߰�E�	Z��1�Ѧ