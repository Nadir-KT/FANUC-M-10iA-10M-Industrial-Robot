��   ?3�A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�DUM�MY10  � &SOP_T  � $��EMGO��R�ESET�MOT|�HOLl���12�STAR^ PDI8G9G�AGBGC�TP;DS�REL�&�U� �� �E�ST���SFSP�C���C��C�NB��SP)*$8*$3%)4%)5%)6%)7%)S��PNSTRz�"D|�  �$$CLr   ����!������ VIR�TUAL�/�!;L�DUIMT  ~�����~�$MAXDRI� b��5�%.1 �%� � �d%Open ?hand 1�����% a?�? �" � �!�# �%CloseQ?d?�?��?�9�7RelaAx�?�?)OOO�9�6L82QO2O�OVO�3 @�?�O�O
_�O�4O �O�Ol__�6�Fh_@�_d_�_�[�3���_ o�_:o�_�_poomo �oUogo�o�o �o�o 6H3l-�Q �u����2�� �h����;�M���ԏ ��������.�ݏR�d� �%���I���m���� ���*�ٟ�`���� 3�E���̯��𯟯�� &�կJ����E���A� ��e�w�쿛�Ͽ�ѿ �X��|�+�=ϲ�a� ���ϗϩ����B��� �x�'�u߮�]�o��� ������>�P�;�t� #�5��Y���}���� ���:�����p���� C�U������� ���� 6��Zl-�Q �u����2� �h�;M�� ����./�R// /M/�/I/�/m//�/ �/?�/�/?`??�? 3?E?�?i?�?�?�?�? &O�?JO�?O�O/O}O �OeOwO�O�O_�O�O F_X_C_|_+_=_�_a_ �_�_�_�_o�_Bo�_ oxo'o�oKo]o�o�o �o�o�o>�obt #5�Y�}�� ��:���p���� C�U�ʏ܏Ǐ ����� 6��Z�	��U���Q� Ɵu������� �ϟ� �h����;�M�¯q� �������.�ݯR�� ���7�����m���� ���ǿٿN�`�Kτ� 3�EϺ�i��ύϟ��� &���J���߀�/ߤ� S�eߟ��ߛ����� F���j�|�+�=��a� �������	�B��� �x�'���K�]����� ������>��b #]�Y�}� �(��#p� CU�y� /�� 6/�Z/	//�/?/�/ �/u/�/�/�/ ?�/�/ V?h?S?�?;?M?�?q? �?�?�?�?.O�?ROO O�O7O�O[OmO�O�O �O_�O�ON_�Or_�_ 3_E_�_i_�_�_�_o �_oJo�_o�o/o�o Soeo�o�o�o�o�o F�oj+e�a �����0��� +�x�'���K�]�ҏ�� �����ɏ>��b�� #���G���Ο}���� ��(�ן�^�p�[��� C�U�ʯy����� 6��Z�	����?��� c�u������� �Ͽ� V��zό�;�M���q� �ϕϧ�����R����
Send E�ventU�5�SENDEVNT���3�i��%	�}�Data�ߘ�D�ATA�߿���%�}�SysVar<��SYSVY��}1�%Get�ߞZ�GET�����%Request Menu�����REQMENU!�����?߀�;ߤ� _������������ F��j+�O� ����0�� fxc�K]�� ����>/�b// #/�/G/�/k/}/�/? �/(?�/�/^??�?�? C?U?�?y?�?�?�?$O �?!OZO	OO�O?O�O cOuO�O�O�O _�O�O V__z_)_;_u_�_q_ �_�_�_o�_@o�_o ;o�o7o�o[omo�o�o �o�oN�or! 3�W����� �8���n���k��� S�e�ڏ���������� F���j��+���O�ğ s��������0�ߟ� f������K�]�ү�� ������,�ۯ)�b�� #���G���k�}��� �(�׿�^�ς�1� C�}���y��ϝϯ�$� ��H���	�Cߐ�?ߴ��c�u��$MACR�O_MAX:��  ��������SOPENB�L ��� ��՗�r�r�A���?PDIMSK���3�Y�SUc�u��TPDSBEX Q \�p�q�U�� ��n����