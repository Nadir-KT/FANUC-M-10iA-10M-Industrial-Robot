��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETGss�ET�H_FLTR.�  $� �  �FTP�_CTRL. �@ $LOG_�8	�CMO>$�DNLD_FIL�TE� � SUBD�IRCAP� o �HO��NT.� 4� H_NA�ME !A?DDRTYPA �H_LENGTH�' �z +L�S D $?ROBOTIG �PEER^� MA�SKMRU~O]MGDEV#� �RDM*�DIoSABL&� OTCPIG/ 3 �$ARPSIZ�&_IPF'W�_MC��F_I�N� FA~LAS�Ss�HO_� I�NFO��TEL�K PV��b	 WORD  �$ACCES�S_LVL?TI�MEOUTuOR�T � �ICEUmS=  ��$#  ����!��� � � VIRTUAL�/�!'0 �%_
���F��d����$�%��;�+ ����#�$�� �-2%;��SHARED 1��)  P!�!�?���!|?�?�? �?�?O�?%O�?1OO ZOOBO�OfO�O�O�O �O_�O�OE__i_,_ �_P_�_t_�_�_�_o �_/o�_SooLo�oxo �opo�o�o�o�o�o *Os6�Z� ~�����9�� ]� ���D�V���z�ۏ ����#���Y�H��}�@���)7z _LI�ST 1=x!1.ܒ0��d�ە�1�d�255.�$������%ړ2 ��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I����o�������O�6���8��0���� �$�� �-� ���-�(�%���&!Ò�)�0H�!� ���r?j3_tpd���!� � �!!KC�� e�0ٙ��&W�!�Cm ��w߉�S�!CON� ��1�==�smon��W�