��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG �ET�H_FLTR.�  $� �  �FTP�_CTRL. �@ $LOG_�8	�CMO>$�DNLD_FIL�TE� � SUBD�IRCAP� o �HO��NT.� 4� H_NA�ME !A?DDRTYPA �H_LENGTH�' �z +L�S D $?ROBOTIG �PEER^� MA�SKMRU~O�MGDEV#PC_3�RDM*��DISABL&>���TCPIG/ �3 $ARPS�IZ&_IPF�'W_MC��F�_IN� FA~L�ASSs�HO_ބ INFO��T;ELK PV��b	 WORD�  $ACCESS_LVL?TIMEOUTu�ORT � �IC�EUS= �   ��$#  �����!�� � � VIRTUAL�/�!'|0 �%
���F�����$�%����+ ������$�� �-2�%;�SHARED� 1�)  CP!�!�?���!|? �?�?�?�?O�?%O�? 1OOZOOBO�OfO�O �O�O�O_�O�OE__ i_,_�_P_�_t_�_�_ �_o�_/o�_SooLo �oxo�opo�o�o�o�o �o*Os6� Z�~����� 9��]� ���D�V��� z�ۏ����#����Y�H�}�@���)7z _LIST 1=_x!1.ܒ0���d�ە1�d�25c5.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I���� o�������O�6����8������ �$ ���-� ���-�!��%�%��&!Ò�)��0H!� ����rj3_tpd����! � �!!KC� e�0ٙ��&W�!Cm ��w߉�~S�!CON� ���1�=�smon��W�