��   %��A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���D�MR_GRP_T�  � $�MA��R_DON�E  $OT�_MINUS o  	GPLN^8COUNP T gREF>wPOO�tlTpBCKLSH_SIGo�SEACHMST�>pSPC�
�M�OVB RADAP�T_INERP ��FRIC�
CO�L_P M�
GR�AV��� HIS���DSP?�H�IFT_ERRO��  �NApM�CHY SwARM�_PARA# ]d7ANGC M=2pCLDE�_CALIB� DB�$GEAR�2�� RING��<��PLCL*; ��STA� m�TRQ_M��LgINK"2&SX<*UY<*Z/)II*IW*�Ie$ �RV*� < $� EN�BpV_DEBU:��!PNU;%� �UNEVEox�  �$�ASS  ����!������ VIR�TUAL�/�!' �1 5�/ ��� �  B?��>?w?b?�?�?�?�?�?�?�5��I�=��!8O&L��{4��V����l�����v� f|n %O�O!OKL�O�O�O�O�O�OzK1_7R _]_o_Z_�_��d�_�_�_<�_��=L���_o3?�o��@�3oXo jo|o�o�o�o5�o�o �o�o#�$�R)SAw62k��� ����#�5�G��" � M�s���������͏�ߏ���'�9��#��$% 1521D}U%a{��� �_��}_ԟ������ ��R�=�v�a����� ��ͯ��������<� '�`�K�]��������� ޿ſϯ�ӿ8�Ͽ\� Gπ�kϤϏϡ����� ����"�	��U��|� ߠߋ��߯������� �	�B�-�f�M�Wߙ� [���W��������,� �)�b�M���q����� ��������(L 7p[m���� ����!�H�l W�{����� /�2//#e/'/�/ #/�/�/�/�/�/�/�/�.??R?=?v?;g�$kRV[�b�8k?��?c?  BFo;gx �?O(O:OLO^OpO�O�O  h 
�  :  B`�����������S������������@$����\�����C���@�@r���C��O__,_>_P_b_ t_�_�_�_�_�_�?�_ �_o(oOLo^opo�o �o�o�o�o�o�o  $6HZl~�� �����o=o2� �V�1oz������� ԏ���
��.�@�R� d�v���������П� ����*�<�C�`�G� Y���q���̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|σ��χ� �ϟ�������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ���(�:�L�^�p��� ������������  $6HZl~�� �������2 �Bhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??<?N?5?r? M�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_jQ