��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1����|UREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"(�AS�BN_CFG1 � 8 $CN?V_JNT_* |�$DATA_C�MNT�!$FL�AGS�*CHE�CK�!�AT_C�ELLSETUP�  P $HOME_IO,�G�%�#MACR=O�"REPR�(-�DRUN� D|�3SM5H UTO�BACKU0 �� $ENAB���!EVIC�T]I � D� �DX!2ST� ?0B��#$INTERV�AL!2DISP_�UNIT!20_D�On6ERR�9FR�_F!2IN,G�RES�!0Q_<;3!4C_WA�471��8GW+0�$Y �$DB� 6COMW!2MO� H.o	 \rVE�1�$F�RA{$�O�UDcB]CTMP�1_FtE2}G1_P�3�B�2�XD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za4 q;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6�_�7_�8_�9�CO�$ <� �o�op�hK3 1#`O_Mc@�AC t � E�#6NGPvABA � �c1�Q8��`,��@Bnr1�� d�P�0Xe���axnpUP@&Pb26���p�"J�pS_R�rPBC��J�rĘߜJV�@U� B��`s}�g1�"YtP_*0wOFS&R @� �RO_K8T��aIT<�3T�NOM_�0�1�p�34 >��D !�� Ќ@��hPV��mCEX�p� �0g0ۤ<�p�r
$TF�2Co$MD3i�TO�3��0U� F� R��Hw2tC1(�Ez�g0#E{"F�"F�F40CP@�a2 �@$�PPU�3N�)ύRևAXd�!DU��AI�3�BUF�F=�@1c |pp���pPIT�� PP�M�M��y��F�SIMQSI�"ܢVAڤT�9I=�w T�`(z�M��P�B�qFAC5Tb�@EW�P1��BTv?�MC�k �$*1JB`p�*1DEC��F���y=�� �H0�CHNS_EMP�1�$G��8��@_�4�3�p|@P��3�TCc�(r/�0-sx���ܐ� MBi��!����J�R� i�SEGFRR��Iv �aR�Tp9N�C��PVF�?�>bx &��f {uJc!�Ja��� !28�pץ�AJ���SIZ�3S�c�B�TM���g��>JaRSINFȑb� ��q�۽�н�����L�3�B���CRC�e�3CCp���� c��mcҞb�1J�cѿ��.����D$ICb�C q�5r�ե��@v�'���SEV���zF��_�եF,pN��ܫ�p?�4�0A�! �r ���h�Ϩ��p�2��@�a�� �د�R�Dx Ϗ��oH"27�!ARV�O`C�'$LG�pV�B�1�P��@�t�aA�0'�|�b+0Ro�� MEp`0"1 CRA 3 CAZV�g6p�O �#FCCb�`�`F�`K�8������ADI��a �A�bA'�.p��p�`�c�`S4PƑ�a�A�MP��-`Y�3P�M���CUR��QU�A1  $@TITO1/S@S�!����"0�DBPXWO��zB0!5�$SK����2G=�DBq�!"�"�PR�� 
p� =����!# S 6q1$2�$z���eL�)$�/PAE���� %�/��PC�!&�?4ENE�q.i'*?PA�!RE�p�2(H ��O��0#$L|3$$@�#�B[�;���FOs_D��ROSr��#������3RIG7GER�6PApS��>��ETURN�2�c�MR_8�TUw�\�0EWM��M�cGN�P���BLAH��<E���P��&$�P� �'P@�Q3�CkD{��DQ���4�1�1��FGO_AWA�Y�BMO�ѱQ#!��DCS_�)7  �PIS� I  gb {s�C��A��[ �B$�S��AbP�@r�EW-�TNTVճ�BV�Q[C�(c`�UW�r�P�J��P�$0��S�AFE���V_SV>�bEXCLU�砝nONL2��SY��*a&�OT�a'�HI_V�4��B����_ *P0� 9�_�z��p �"�@SG�� +nrr�@�6Acc*b��G�#@E�V�.iHb?fANNUNX$0.$fdID�U�2�SC@�`�i�a��jP�f��z��@I$2,O��$FibW$}�OT�9@�1 $DUMMYk��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6�a�!M�SW�E. 8Q�KgEYI5���TM�100s�qA�vIN��#��b��/ D��H7OST_P!�rk���ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  �8	=ȳ���DT�k0�!1 � $|S��ESAMPL��@j�۰f璱f���I�0|��[ $SUB��k�#0�C��T�r#a�SAVʅ��c���CX��P�fP$n0E��w YN_B#2 M0Q�DI{dlpO(���9#$�R_I��� �ENC2s_S� 3  5�C߰�f�- �SpU����!4�"g�޲�19T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9�g�DSP�v��PC���r"��(���ƓV7ALUߗHE�ԕ�M+�IPճ��OP5P ��TH��֤D��P�S� �۰F�B�df�J� ��мC1+6 H�bLL_DUs�~a3@{�0�3:���OTX"����sʡR_N_OAUTO�!7�pC$)�$�*��c4�*(�Cy�8�C, �"��q&�L�� 8/H *8�LH < 6����c"�`, `Ĭ� kª�q��q��sq��T~q��7��8��9���0����1��1̺1�ٺ1�1�1 �1*�1�2(�2����U2̺2ٺ2�2�U2 �2�2�3(ʥ3��3��̺3ٺ3��3�3 �3�3��4(�a��?��!9� <�9�&�z��I`��1���M��QFE@�'@� : ,6��Q?g �@P?9��5�9�E�@A�q��A� ;p$T�P�$VARI�:�Z���UP2�P< ���TDe����K`Q���"���BAC�"= T�p��e$�)_,�bn�kp+ IF�IG�kp�H  ��P°Y�@`�!>Gt ;E��sC�ST�D� D���c�<� 	C��{�� _���l���R  ���FORCEUP?b^��FLUS�`H��N>�F ���RD_CM�@E������ ��@vMP��REMr F �Q��1�����7Q
�K4	NJ�5EFF�ۓ:�@IN2Q��O�VO�OVA�	TgROV���DTՀ�DTMX� � �@�
ے_PH"p��CL��_TpE�@d�pK	_(�Y_T��Tv(��@A;QD� ������!0tܑ&0RQ���_�a��2��M�7�CL�dρ�RIV'�{��EAmRۑIOHPC�@d����B�B��CM9@����R �GCLF�e!DYk(M�a6p#5TuDG��8� �%aFSSD �s�? P�a�!�1����P_�!�(�!1��E��3�!3�+5�&�GSRA��7�@��;ᚔPW��ONn��EBUG_SD2HP��{�_E A �L����TERM�`5Bi5R�O�RI#e0Ci5K@�GSM_�P��e0Di5��0TA�9E�9U}P\�F� -�A�{�AdPw3S@B$gSEG�:� EL{UwUSE�@NFIJ�B$�;1젎4�4C�$UFlP=�$,�|QR@��_G90qTk�D�~SNST��PAT����APTHJ3Q�E�p%B�`�'EC���ARx$P�I�aSHFTy��A�A�H_SHOR(Р꣦6 �0$�7P9E��E�OVR=��aRPI�@�U�b �Q�AYLOW���I�E"�r�A��?���ERV��XQ�Y��mG>@@�BN��U���R2!=P.uASYMH�.uFAWJ0G�ѡEq��A�Y�R�Ud>@��EC���EP;�uP;��6WOR>@M`��0SMT6�G3�G1R��13�aPAL@���P��q�uH � :���TOCA�`yP	P�`$OP����p�ѡ�`0O,��RE�`R4C�A�O�p낎Be�`R��Eu�h�A��e$P�WR�IMu�RR�_�cN��q=B I�&2H���p_ADD�R��H_LENG��B�q�q�q$�R��S��JڢSS��SK�N��u���u̳�uٳS�E�A�jrS��MN�!K�����b����OLX��p�<���`ACRO3pJ� �@��X�+��Q��6�OUP3�b_�IX��a�a1��}򚃳� ��(��H��D��ٰ���氋�IO2S��D�����	�7��L $l��`Y!_O�FFr�PRM_����aTTP_�+�H:�M (|pOcBJ]"�p��$���LE~Cd���N � ��֑AB_�TqᶔS�`H�LVh�KR"uH�ITCOU��BG�LO�q���h�`����`��`SS� ����HW�#A:�O�ڠ<`INCPU>2VISIOW�͑���n��to��to�ٲ ��IOLN��P �8��R��p$S�Lob PUT_&n�$p��P& ¢���Y F_AS�"Q��$L������Q"  U�0	P4A��^����ZPHY��-���y��UOI �#R `�K����$�u�"pPpk���$�X������UJ5�S-�v��NE6WJOGKGN̲DIS����Kp�L��#T (�uAVF��+`�CTR�C
�FgLAG2��LG�d�U ���؜�13LG_SIZ����bŰ4�a��a�FDl�I `�w� m�_�{0a�^� �cg���4�����Ǝ����{0��� SCH_H���a7�N�d�VW���E�"����4��UM�Aљ`LJ�@�DAUf�EAU�p��d�|�r�GH�ba���B�OO��WL ?�6 IT��y0�wREC��SCR �ܓ�D
�\���MARGm�!��զ ��dH%�����S����W���U� �JGM[�M�NCHJ���FNK�EY\�K��PRGƂ�UF��7P��FW�D��HL��STP���V��=@��А�RES��HO`����C9T@��b ��7�[�UL����6�(RD� ����Gt��@PO��������MD�FOCU��RwGEX��TUI��	I��4�@�L� ����P����`���P��NE��CANAx��Bj�VAILI��CL !�UDCS_CHII4��s�O�D(!�S���S�x�D���BUFF�!�X�?PTH$�m���v`�ěԬ�A
trY�?P��j�3���`OS1Z2Z3�Z��� Z � ���[aEȤ��ȤIKDX�dPSRrO�X��zA�STL�R}��Y&�� Y$E�C���K�&&p+P|�� [ LQ� �+00�	P���`#qdt�
�U�dw<���_ \ �`4Г�\���t�#\0C4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#�1D���'B�LD�%�$�%ORGڰ5�2�P VŇVY8�s�T�r�$}d^ ���$6��$�%�S�`T� �B0�4>�6RCLMC�4]?0o?�9세�MI�p}dg_ d=њRQ�=�DSTB�p�c ;F�HHAX�R� JHdLEXCE�SrWPCM!p�a`�/B�Ta�B��`5a�p=F_A7Ji���KbOtH� K�db q\Q���v$MBC��LI|�)SREQU�IR�R�a.\o�AXD�EBUZ�ALt M��c�b�{P����2�ANDRѧ`�`d0;�2�ȺSDC��N�INl�K�x`��X� �N&��aZ���UP�ST� ezrL�OC�RIrp�E�X<fA�p�9A����`AQ��f XfY�OND�rMF,� �Łf�s"��}%�e/�� �a�FX3@IGG>�� g ��t"���ܓs#N�s$R�a%��iL��hL�v�@��DATA#?pE��%�tR��Y�Nh t $MD`qI}�)nv� ytq�yt�HP`�Pxu��(�zsANSW)�yt@��yu�D+�)Yr���0o�i[ �@CUw�V�p� 09AARR2��j� Du�{Q��7Bd$OCALIA@��G�:�2��RIN��"��<E�NTE��Ck��r^�آ9AA]���_N�qlk���9�D����Bm��DIVFD�H�@���qnI$�V,��S�$���$Z�X�o�*�����oH �$�BELT�u!ACCEL�.�~�=��IRC�� ���D�T<�8�$PS�@�"L�@�r��#^�S�xEы T�PATH3����I���3x�p�A_@W��ڐ���2nC���4�_MG�$D�D��T���$FW��Rp9��I�4��D}E7�PPABN��ROTSPEE�[g�� J��[�C@�4��@$USE_d+�VPi��SYY����1 �aYN!@A��ǦOFF�qǡM�OU��NG���O9L����INC�tMa�6��HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]�ౌB��VE��#�y�2�3_UP񕋳LOWL���p� B���Du�9B#P`�x ����BCv�r�MOSI���BMOU��@�7P�ERCH  ȳOV��â
ǝ���� D�ScF�@MP����B� Vݡ�@y�j�LU0k��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A���x�����N`�F�RT1I�A$��MOUІЀHB�BS0�p7D5����ë�Z�DUM2�ԓS_BCKLSH_Cx�k���� ϣ���=���ޡ �	ACLAL"q��1М�@��CHK� �S�RTY��^�%�E1Qq_�޴_UM��@�C#��SCL�0�r�LMT_J1_L��9@H�qU�EO�p�b�_�e�k�e�SPC��u���N�PC�N�Hz \P�2�C�0~"XT��CN_:�N9��I�SF!�?�V���U� /���x�T���CB!�SH�:��E�E1TрT����y���T��P�A ��_P��_ � =������!�����J6 L�@��OG|�G�TORQU��ONֹ��E�R��H�LE�g_W2���_郠����I�IJ�I��Ff`xJ�1X�~1�VC3�0BD:B�1�@SB�JRKF9�0D�BL_SM��2M��P_DL2GR�V����fH�_��d���COS���LNH� �������!*,��aZ���fMY��_(�TH��)T�HET0��NK2a3���"��CB�&CB�CAA�B�"�0�!��!�&SB� 2N�%GTS�Ar�CI Ma�����,4#97#$DU���H\1�  �:Bk62�:AQ(rSf'$NE�D�`I��HB+5��$̀�!A�%��5�7���LPH�E�2���2SC% C%�2-&FC0JM&̀EV�8V�8߀LVJUV!KV/KV=KVKKVYKVgIH�8FRPM��#X!KH/KH=KUHKKHYKHgIO�<�O�8O�YNOJO�!KO/KO=KOKKO
YKOM&F�2�!+i%�0d�7SPBALA�NCE_o![cLE60H_�%SPc� &��b&�b&PFUL�C�h�b�g�b%p�1=k%�UTO_���T1T2�i/�2N ��"�{�t#�Ѱ`�0(�*�.�T��OÀ<�>v INSEG"�ͱ�REV4vͰl�DI�F�ŕ�1lzw��1m�0OBpq�я?��MI{���nLCHgWARY�_�AB��~!�$MECH�!�o ��q�AX��P�����7Ђ�`n 
p�d(�U�ROB���CRr�H���o(��MSK_f`�p� P �`_��R /�k�z�����1S�~��|�z�{���z��qIN�Uq�MTCOM�_C� �q  ����pO�$NO�REn����pЂ7r 8p GRe�u�SD�0AB�$?XYZ_DA�1a���DEBUUq�������s z`$��COD�� L���p��$BUFIwNDX|�  <��MORm�t $فUA��֐����r�<��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p�=�C�}pt�@b�D��FRIrӚ�T��RO@ \�E�}��y�OPWO�Yq�v0Y�SY�SBU/@v�$SO!Pġd���ϪUΫ}p�PRUN����PA�D���rɡL�_O�Uo顢q�$^)�IMAG��w���0P_qIM��L�I�Nv�K�RGOVCRDt��X�(�P*�J�|��0L_�`]�L�0�RB1�0��M��ED}��p J��N�PMֲ��\c��w�SL�`q�w x $OVSL4vwSDI��DEX�@���#���-�V} *�N4�\#�B�2�G�4B�_�M�y�q|�E� x Hw���p��ATUSW����C�0o�s���BT�M�ǌ�I�k�4p��x�԰q�y Dw�!E&���@E�r��p7��жЗ�EXE���ἱ�����f q�z3 @w���UP'��3$�pQ�XN����������� �PG�΅{ h $S#UB����0_���!��MPWAIv�PL7ã�LOR�٠F\p�˕$RCVFA�IL_C��٠BW�D΁�v�DEFS}P!p | Lw����Я�\���UN!I+�����H�R�+�V}_L\pP����	P��p�}H�> �*��j�(�s`~�N�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��G���PLI��p� � $ˀP_S�WI�pq�J_PL~��AL_ ���J��A��B��� C���D�$E���.�C_�U�� � � ���*��J3K0����TIA�4��5��6��MOM��������ˀB��AD��������6��PU� NR�������?H��m��� A$PI�6 q��	�����K4��)6�U��w`��S/PEEDgPG�� ������Ի�4T��� � @��SA�Mr`��\�]��MOV_�_$�npt5�H�5���1���2��@������'�S�Hp�IN�'�@�+�����4($4+T+G�AMMWf�1'�$GGET`�p���Da�z��

pLIBR>ѺII2�$HI=�_�g�t��2�&E;��(A�.� �&LW�-6<��)56�&]��v�p��V���$PDCK���q��_?�����q�&���7��4����9+� �$_IM_SR�pD�s0�rF��r�rLE���aOm0H]��0�-ܬpq��PJqUR_SCRN�FA����S_SAVE_DX��dE@�NOa�CA A�b�d@�$q�Z�Iǡ s	�I� �J�K� ��� �H�L��>�"hq� �����ɢ�� @bW^US�A�G�L�0m����a��)q`��3��WW�I@v�_�q�.M�UAo�� � $sPY+�$W�P�vNG�{��P:��R`A��RH��RO�PL��@���q� ��s'�X;�	OI�&�Zxe ���m�G� p��ˀ�3s��O�O�O�O�O�aa�_т� |��q�d@�� .v��.v��d@��[wFvr��E���% Z��r;B�w�|�tPn���PMA�QUa ��Q8��1٠wQTH�HOLG�oQHYS��ES�F�qUE�pZB��Oτ�  ـPܐ(�AP����v�!�t�O`�q��u�"���FA��IGROG�����Q2����o�"��p��INFOҁ�׃V����R��H�OI��� (�0SLEQ����@��Y�3����Á��P�0Ow0���!E�0NU��AUT<�A�COPY�=�(/�'��@Mg�N��=��}1������ ��RG4��Á���X_�P�C$;ख�`��W���P��@�������E�XT_CYC b�HᝡRpÁ�r��_NAe!А����ROv`	�� �s ���POR_�1�E2�SRV �)l_�I�DI��T_� k�}�'���dЇ�����U5��6��7��8i��H�SdB���2�$R��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,�0FL`�o@SYN��K�M��Ck��PWR+�9ᘐ���DELA}�dY��pAD�av�Q�SKIP4� ĴA�$�OB`NT����P_$�M�ƷF@ \bIpݷ�ݷ�ݷd� ���빸��Š�Ҡ��ߠ�9��J2�R� ��� 4V�EX� TQQ����TQ������� ��`���R;DC�V� �`��X)�R�p�����r���m$RGEAR_� IOBT�2FLG���fipER�DTC����Ԍ���2TH2yNS}� 1����G T\0 �$��u�M\Ѫ`I�d PA�REF��1Á� l�h��E�NAB��cTPE �04�]����Y�]��� �Qn#��*��"�����
��2�Қ�߼�����(����3�қ'�9�K�]�o���4�Ҝ�������������5�ҝ!�3�E�W�i�{�
�6�Ҟ��������(�����7�ҟ-�?Qcu�8�Ҡ �������P�үSMSKÁ�l�Ԁa��EkA��REoMOTE6������@�݂TQ�IOD}5�ISTP�QR�9W@��� �pJ� ���p����E�"�$DSB_SIG!N�1UQ�x�C\�TP~���RS232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+�TQ��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�P��S�0�����p_�XPC)�$FRE?EFROMS	pna��GET�0��UP%D�A�2E#P� :�ߧ� !$USAN�na&�����ERI�0�RpRY$q5*"_j@�Pm1�!N�6WRK9KD����6��QFRIEND�Q�RUFg�҃�0oTOOL�6MY�t�$LENGTHw_VT\�FIR�p�C�@ˀE> +IUF�IN-RM��RGyI�1ÐAITI�b$GXñ3IvFG2v7�G1���p3�B�GP1R�p�1F�O_n 0��!RE��p�53҅�U�TC��3A�A�F��G(��":��� e1n!��J�8�%���%�]��%�� 74�XS O0�L��T�3�H&��8���%b453G�E�W�0�WsR�TD ����T��M����Q�T�]�$V 2�����1�а91�8�02*�;2k3�;3�:i fa�9-i�aQ��NS���ZR$V��2BVwEVD�2A Q�B;�����&�S�`��F�"�kX�@�2a�PS�E���$r1C��_$Aܠ6wPR��7vMUb�cS�t '�16�9�� 0G�aV`��p�d`���50�@���-�
25S�� E��aRW����B��&�N�AX�!�A�:@LAh��rTHI�C�1I���X�d1T�FEj��q�uIF_CH�3�qI܇7�Q�pG1RxV���]�岺:�u�_JF~�P�RԀƱ�RVAT��� ��`���0�RҦ�DOfE��CO9UԱ��AXI����OFFSE׆TRIGNS���c����h����H�Y��IGGMA0PA�pJ��E�ORG_UNE9V�J� �S����?�d �$CА�=J�GROU�����TOށ�!��DSP���JOGӐ�#��_	Pӱ�"O�q����@n�&KEP�IR��dܔ�@M}R��AP�Q�^�Eh0��K�SY�S�q"K�PG2�B�RK�B��߄�p`Y�=�d����`AD_�<����BSOC����N��DUMMY1�4�p@SV�PDE�_OP�#SFSP_D_OVR-���1C��ˢΓOR٧3�N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1q"�LCHDL��REGCOVʤc0��Wq@1M������RO�#��rȐ_+��� @0��e@VER�$O�FSe@CV/ �2WD�}��Z2����TR�!���E_�FDO�MB_CiM���B��BL�bܒ#��adtVQR�$0�p���G$�7�AM�5��� eŤ��_M�;��"'����8$C�A��'�E�8�8$HcBK(1���IO<�q����QPPA�ʀ����
��Ŋ����DVC_DBhC;�� #"<Ѝ�r!S�1[ڤ��S�3[֪�ATIO"q 1q� ʡU�3���CABŐ�2�CvP ��9P^�B���_� �?SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW�_C��U��S@��SA��A�pl$UNITm�l_�AT���e��ƐCYCLq�NE�CA���FLTR_2_FIO�7(�ӌ)&B�LPқ/�.�_�SCT�CF_`�F0b�l���|�FS(!E�e�CHA�1��4�D��"3�RSD��$"}�����_Tb�PR�O����� EMi_䙰a�8!�a �!�a��DIR0�R�AILACI�)RM�r�LO��C���Q`q��#q�դ�PR=�%S�A�pC/�c =	��FUNCq�0rRINP�Q�0��2f�!RAC �B ��p[���[WARn�F��BL�Aq�A����DAk�\���LD0���Q�d�qeq�TI"rp��K�hPRIA�!r"AF��Pz!=�;@��?,`�RK���Mǀ9I�!�DF_@B�l%1n�LM�FAq@OHRDY�4_�P@�RS�A�0� �MU�LSE@���aG ��ưt��m��$�1$�1$�1o����� x*�EG00�����!AR���Ӧ�09p�2,%� 7�AXE���ROB��WpA��_l-��SY[�W!‎&MS�'WRU�/-1��@�STR������Eb� 	�%��J��AB� ���&9�����kOTo0 	$��ARY�s#2��Ԓ��	ёFI@��$�LINK|�qC1��a_�#���%kqj2XYZ��t;rq�3��C1j2^8'0B��'�4����+ �3FI���7�q����'��_Jˑ���O3�Q'OP_�$;5���A#TBA�QBC��&��DUβ�&6��TURN߁"r�E11:�p��9GFL�`_���* Ȩ@�5�*7��Ʊ +1�� KŐM��&�8���"r��ORQ��a�(@#p=� j�g�#qXU�����mT'OVEtQ:�M��i�@��U��U��VW�Z �A�Wb��T{�, ��@ ;�uQ���P\�i��UuQ��We�e�SERʑe	��E� O���UdAas��4S�/7����AX��B� 'q��E1�e��i��i rp�jJ@�j�@�j�@�j P�j@ �j�!�f��i ��i��i��i��i �y�y�'y�7y�TqHyDEBU8�$32���qͲf2G + AB����رnS9VS�7� 
#�d� �L�#�L��1W��1W� JAW��AW��AW�QW��@!E@?D2�3LAB�29U4�Aӏ��Co 0 o�ERf�>5� � $�@_ mA��!�PO���à�0#�
�_MR}At�� d � 9T��ٔERR����;TY&���I��V8�0�cz�TOQ�d�PL[ �d�"�� ?�w��! � pp`T8)0���_V1Vr�a(Ӕ����2ٛ2�E�ĺ��@�H�E���$QW�����V!��$�P��o�cI��a�Σ	 HELL_�CFG!� }5��B_BASq��SR3��� �a#Sb���1�%���2��3��4��5*��6��7��8����RO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CYO. U�OUG�P~ �����m�������TPհ_KAR�l�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h��]��l0SEM�4�(�Ml4�6�TYN�SO���DIZ�~�A������m_TM�MAN�RQ��k0E�����$KEYSWIT�CH���m���HE���BEAT��EF- LE~�����U���F!Ĳ���B�O_H�OM=OGREFUPPR&��y!� [��C��O��-ECO�C��Ԯ0_IOCMWD
�a���m���� � Dh1���U�X���M�βgPgCFgORC��� ���m�OM.  � Q@�5(�U�#P, Q1��, 3��45���NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�� �� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E'��V�P��UPDs� � �`NЦ�5�Y�SLOt�� � �L��d���A�aT�A�0d��|�ALU�:ed�~�CUѰjgF�!aID_L�ÑeH�I�jI��$FILcE_���d��$2�vfSA>�� hO�~�`E_BLCK���b$��hD_CPU yM�yA��c�o�db�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA�i�J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP��_(�g����pr��� `�`GROU�w`��B��NFL�IC��f�REQUwIRE3�EBU�0�qB���w�2����p����q5�p�� \^��APPR��C}��Y�
ްEN٨CL9O7��S_M��H����u�
�qu�� ���MC�����9�'_MG��C�Co��`pM�в�N�BRKL�GNOL|�N�[�R���_LINђ�|�=�J����Pܔ�������� ���������6ɵ��̲8k�+��q���G� ��
��q)�<�7�PATH3�L�@B�L��H�wࡠ�J�CN�CA�Ғ�ڢ6B�IN�rUCV�4aZ��C!�UM��Y,���aE�p����������PAYLOAJ2L`R_A	N�q�Lpp����$�M�R_F2LS3HR��N�LOԡ��Rׯ�`ׯ�ACRL�_G�ŒЛ� ��H�j`߂$HM���FWLEXܣ�qJ�u� :���� ���������1�F1�V�j�@�R�d�v�������E����ȏ ڏ����"�4�q��� 6�M���~��U�g�y�$ယT��o�X��H� �����藕?����� ǟِݕ�ԕ�����%�7��JJ�� �� V�h�z���`A�T�採@�EL�� �S��J|�Ŝ�J�Ey�CTR��~�T�N��FQ��HAN/D_VB-���v`n�� $��F2M�X���ebSW�q#��'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aDM)F�AW�Z`i�Aw�AA��X X�'pi�Dw��D��Pf�G�p�)S�Tk��!x��!N��DY�pנM�9$`%Ц� H��H�c�׎���0� ��Pѵڵ������������� ����1��R�6��QA'SYMvř���v���J���cі�_SH >��ǺĤ�ED����������J�İ%��C��IDِ�_VI��!X�2PV_UNIX�FThP�J��_R�5 _Rc�cTz�pT�V��@�@��İ�߷��U ��������Hqpˢ���aEN�3�DI����O4d �`J��� x g"IJAA ȱz�aabp�coc�`as�cr�a� ��/OMME��� �b4�RqT(`PT�@� S��a7�;�Ƞ�@�h��a�iT�@<� $DUMMY9Q��$PS_��RF�C�E`$v p�p���Pa� XƠ����STE���S�BRY�M21_V�F�8$SV_ER�F�O��LsdsCLR�JtA��Odb`O��p � D �$GLOBj�_LO���u�q�cAp�r�@�aSYS�qADR�``�`TCH  �� ,��ɩb�W7_NA���7���SR���l ���
*?�&Q� 0"?�;'?�I)?�Y)�� X���h���x������) ��Ռ�Ӷ�;��Ív��?��O�O�O�D(�`XOSCRE栘p�����ST��s}Hy`���Ea/_H�A�q� TơgpTYP�b���G�a�G���Od0ISb_䓀dEaUEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI� m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1A�ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���}АVSHIF��Nc�P�`ג�E��ȐR����OSURz��Wk`RADIL����_�a��:�9a���`a�r��LULQ$�OUTPUT_BM����IM�AB ��@�rTILSCO��C7��� ����&��3�� A���q���m�I�E2G�o�y@Md�}���yDJU��N�/WAIT֖�}���{�%! NE�u�Y�BO�� ��� $`�t�SB�@TPE��NEC�p�J^FY�nB_T��R�І�a$�[$YĭcB��dM����F� �p�$�pb�O�P?�MAS�_DUO�!QT�pD���ˑ#%��p!"DELcAY�:`7"JOY� @(�nCE$��3@ 0�xm��d�pY_[�!"��`�"��[���P?{ �ZABC%�?�  $�"R���
E`�$$CL�AS�������!E`n�� � VIRqT]��/ 0ABS�����1 5�� < �!F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZi{0-�GAXL�p2��!�637  �{tIN��q�ztPRE�����v��p�uLARMRE?COV 9�r�wtNG�� .;	? =#�
�.��0PPLIC��?�5�p��Handling�Tool o� �
V7.50P/�23 �!�PBv��
��_SWt�w UP�!� x�#F0��t���An�v� 864��� �it�y� N��" 7wDA5�� j� ?QB@ϐo��Noneisͅ�˰ ��T�]~�!LAAxyr�P_l�V�uT��s9�UTO�"�Њt�y~��HGAPON
0�g�1��Uh�D 1-581�����̟ޟry����Q 1���p�,�� ����;�@��q_��"��" ��c�.�H���D�?HTTHKYX��" �-�?�Q���ɯۯ5� ���#�A�G�Y�k�}� ������ſ׿1���� �=�C�U�g�yϋϝ� ������-���	��9� ?�Q�c�u߇ߙ߽߫� ��)�����5�;�M� _�q�������%� ����1�7�I�[�m� ���������!���� -3EWi{� �����) /ASew��� �/��/%/+/=/ O/a/s/�/�/�/�/? �/�/?!?'?9?K?]? o?�?�?�?�?O�?�?`�?O#O]���TO��E�W�DO_CLE�AN�����CNM ; � �_�_/_A_S_�DSP�DRYR�O��HIc��M@�O�_�_�_�_ oo+o=oOoaoso�o`�o���pB��v �u���aX�t������9�PLUGG���G���U�PRCvPB�@"��_�orOr_^��SEGF}�K[ mwxq�O�O����8�?rqLAP�_�~ q�[�m��������Ǐ�ُ����!�3�x�T�OTAL�f yx�U�SENU�p�� ��H���B��RG_S�TRING 1~u�
�Mn��S5�
ȑ_ITwEM1Җ  n5� � ��$�6�H�Z�l� ~�������Ưد����� �2�D�I/�O SIGNAL�̕Tryou�t Modeӕ�Inp��Simu�latedבO�ut��OVE�RR�P = 10�0֒In cy�cl��בPro?g Abor��ב���Status�Փ	Heartb�eatїMH �Faul��Aler'�W�E�W�i�{���ϟϱ������� �CΛ�A����8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j�|���WOR{pΛ�� (ߎ����� ��$�6� H�Z�l�~���������������� 2PƠ�X ��A{� ������ /ASew���8��SDEV[� o�#/5/G/Y/k/}/ �/�/�/�/�/�/�/?�?1?C?U?g?y?PALTݠ1��z?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O8�O_�?GRI�`Λ DQ�?_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o2_l�R��a\_�o"4 FXj|���� �����0�B�T��oPREG�>��  f���Ə؏���� � 2�D�V�h�z��������ԟ���Z��$A�RG_��D ?	����;���  	]$Z�	[O�]O���Z�p�.�SBN_�CONFIG �;�������C�II_SAVE � Z�����.�T�CELLSETU�P ;�%H?OME_IOZ�Z�?%MOV_���
�REP�lU�(�U�TOBACKܠ���FRA;:\z� \�z�Ǡ'`�z���ǡ�i�INI�0z����n�MESSA�G���ǡC���OD�E_D������%�Ox�4�n�PAUSX�!�;� ((O>��ϞˈϾϬ��� �������*�`�N����rߨ߶�g�l TSK  wͥ�_�q��UPDT+��d�!�A�WSM_CF��;���'�-�GRP 2:�?�� N�BŰA��%�XoSCRD1�1
7�' �ĥĢ���� ������*������� r�����������7��� [�&8J\n���*�t�GROUN��UϩUP_NA��:�	t��_�ED�17�
 ��%-BCKEDT-�2�'K�`���-t�z�eq�q�z���A2t1�����q��k�(/��ED3 /��/�.a/�/;/M/ED4�/t/)?�/�.?p?�/�/ED5 `??�?<?.�?O�?�?ED6O�?qO�?�.MO�O'O9OED7 �O`O_�O.�O\_�O�OED8L_,�_�^�-�_ oo_�_ECD9�_�_]o�_	-09o�oo%oCR_  9]�oF�o�k� ~� NO_DEL���GE_UNUS�E��LAL_OUT ����WD_ABOR���~��pITR_R�TN��|NON�Sk���˥CA�M_PARAM �1;�!�
 8�
SONY XC�-56 2345�67890 �ਡ@���?�>�( А\�
�Ԫ�{����^�HR�5q�̹��ŏR57�ڏ�Aff���KOWA SC3W10M
�x�̆�d @<�
�� �e�^��П\�����*�<��`�r�g�CE_RIA_I��!�=�F���}�z� ��_LI�U�]�����<z��FB�GP 1��Ǯ�M�_�<q�0�C*  �����C1��9��@��G����CR�C]��d*��l��s��R��翪��[Դm��v���������� C�����(�����=�H=E�`ONFIǰ��B�G_PRI 1�{V���ߖϨ�������������CH�KPAUS�� 1K� ,!uD�V� @�z�dߞ߈ߚ��߾� �����.��R�<�b�4���O������^��_MOR��� ���BZ?�<���� 	 ��� ��*��N�`����䡑��?��q?;�;�����K��9�P��|�ça�-:���	�

��M��@�pU�ð��<��,~���DB���튒)�
mc:cpmi�dbg�f�:�/  ��¥��p�/�  �U�U�	s� )�� �s>�  .�/U�?���p#�p$Ug��/���p�Uf��M/w�O/�
DEFg l��s)��< buf.txt s/�t/��ާ�)��	`�����=L�m��*MC��1��a��?43��1����t�īCz  B�HH�CPUeB���CF�;.�<C���C�5rY
K�D�ny�DQ��D���>��D�;�D���=F���>F�$G}�RB�Gz&�0��Y	��!�&w�K1���s���V�������BDLw�M@x8��1Ҩ�����g@D�p@�0E�YK�EX�E�Q�EJP F��E�F� G���>^F E��� FB� H�,- Ge��H�3Y,!5��  >�33 ���N~  n8�~@��#5Y�E>�ðA��Yo<#�
"Q ����+_�'RSMOF�S�p�.8��)T1>��DE ��F� 
Q��;�(P � B_<_��R��X��	op6C4P�Y
�s@ ]AQ�2s@CR�0B3�MaC{@@*c�w��UT�pFPROG %�z�o�o�igI�q���v��ldK�EY_TBL  ��&S�#� �	
��� !"#�$%&'()*+�,-./01i�:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������vq���͓���������������������������������耇���������������������p`LCK�l4�p`�`�STAT ��S_A�UTO_DO����5�INDT_ENB!���R�Q?�1��T2}�^�STOP�b���TRLr`LE�TE��Ċ_SCREEN �Z�kcsc��U���MMENU 1� �Y  < �l�oR�Y1�[���v� m���̟�����ٟ� 8��!�G���W�i��� �����ïկ��4�� �j�A�S���w����� 迿�ѿ����T�+� =�cϜ�sυ��ϩϻ� ������P�'�9߆� ]�o߼ߓߥ������ ��:��#�p�G�Y�� ����������$��� �3�l�C�U���y��� �������� ��	V�Y)�_MANUAyL��t�DBCO[��RIGڇ
�DBN�UM� ��B1 e
��PXWORK 1!�[�_U/�4FX�_AWA�Y�i�GCP r b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�mg�&/�~&lMZ�IdPx@|P@#ONTIMه�� d�`&�
��e�MOTNEN�D�o�RECOR/D 1(�[g2�/{�O��!�/ky "?4?F?X?�(`?�?�/ �??�?�?�?�?�?)O �?MO�?qO�O�O�OBO �O:O�O^O_%_7_I_ �Om_�O�_ _�_�_�_ �_Z_o~_3o�_Woio {o�o�_�o o�oDo�o /�oS�oL�o ����@��� +�yV,�c�u���� ����Ϗ>�P����� ;�&���q���򏧟�� P�ȟ�^������I� [����� ���$�6��������jTOL�ERENCwB����L�͖ CS_CFG )��/'dMC:\�U�L%04d.C�SV�� c��/#A� ��CH��z� �//.ɿ��(S�RC_OUT *���1/V�SGN �+��"��#��17-FEB-20 18:570�27-JANp�2�1:48+ P;��ɞ�/.���f�pa�m���PJPѲ��V�ERSION �Y�V2.0�.�ƲEFLOG�IC 1,� 	:ޠ=�ޠL���PROG_ENqB��"p�ULSk'� ����_WRS�TJNK ��"fE�MO_OPT_S�L ?	�#
 	R575/# =�����0�B����TO  �ݵϗ��V_F EX�d��%��PATH ;AY�A\����\�5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAqU��z�^"MSWX��.�<�4,#�Y�/�
!J�6%Z�I~m��$SBL__FAUL(�0�^9'TDIA[�1<��<� ���1�234567890
��P��HZ l~������ �/ /2/D/V/h/�Z� P� ѩ� yƽ/��6�/�/�/? ?/?A?S?e?w?�?�?��?�?�?�?�?�,/�U3MP���� �A�TR���1OC@PM�El�OOY_TEM=P?�È�3F���G�|DUNI��.�Y�N_BRK 2�_�/�EMGDI_�STA��]��ENC�2_SCR 3�K7(_:_L_^_l& _�_�_�_�_)��C�A14_�/oo/oAo�Ԣ�B�T5�K� ϋo~ol�{_�o�o�o '9K]o� �������� #�5��/V�h�z��л` ~�����ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T���x��������� ү�����,�>�P� b�t���������ο� ���(�f�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������:� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ���*<N` r������� &8J\n� ���������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?��?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O��O__NoETMO�DE 16�5��Q �d�X
�X_j_|Q�PRROR�_PROG %fGZ%�@��_  �U�TABLE  �G[�?oo)oRjR�RSEV_NUM�  �`WP��QQY`�Q_AUT�O_ENB  ��eOS�T_NOna �7G[�QXb W *��`��`��`	��`d`+�`�o�o�o�dHISUc�aOP�k_ALM 18G[� �A��l�P+�ok}����r�o_Nb�`  G[��a�R
�:PTCP_VER !GZ�!�_�$EXTL�OG_REQv9�i\�SIZe�W��TOL  �aD}zr�=#דQ?XT_BWD�p���xf́t�_DI�� 9�5�d�T�a<sRֆSTEP��|:P�OP_DOv��f�PFACTO�RY_TUNwd�M�EATURE �:�5̀rQ�Handlin�gTool �� �\sfmEn�glish Di�ctionary���roduA�A Vis�� M�aster�����
EN̐nalo�g I/O����g�.fd̐uto �Software� Update � F OR�ma�tic Back�up��H596�,�ground� Editޒ  �1 H5Ca�mera�F��OwPLGX�ell�ީ�II) X�om�mՐshw���co�m��co���\typ���pane���  opl��ty�le selec�t��al C��n�J�ՑonitorΧ�RDE��tr~��Reliab����6U�Diagn�os(�푥�552�8�u��heck� Safety �UIF��Enha�nced Rob� Serv%�q �) "S�r�Use�r Fr[�����a���xt. DIOm �fiG� sŢendx�Err��LF� pȐĳr�됮� ����  !���FCTN Menu`�v-�ݡ����TP Inېfa�c�  ER J�GC�pבk �Exct�g��H5�58��igh-S�pex�Ski1�  2
P��?����mmunic'�ocns��&�l�ur�ې��ST Ǡ�¯conn��2��TwXPL��ncr��stru����"F�ATKARE�L Cmd. L�E�uaG�545\~��Run-Ti���Env��d
!����ؠ++�s)�S�/W��[�Li�censeZ��� �4T�0�ogBoook(Syڐm)���H54O�MACR�Os,\�/Off�se��Loa�MqH������r, k��MechStop� Prot���� �lic/�MiвS�hif����ɒMi�xx��)���xSP�S�Mode Sw�itch�� R5�W�Mo�:�.�� G74 ���g���K�2h�ulti-�T=�M���LN (�Pos�Regiڑ������d�ݐ�t Fun�ǩ�.8�����Num~����� lne��ᝰ Adjup�����  - W��t�atuw᧒T�oRDMz�ot��_scove U��9���3Ѓ�ue�st 492�*�oز����62;�SN�PX b ���8 �J7`���Libr���J�48���ӗ� ȾԄ�
�6O�� P�arts in /VCCMt�32����	�{Ѥ�J990���/I� 2 P~��TMILIB���H���P�Acc�D�L�
TE$T�X�ۨ�ap1S�Tye����pkey��蟑wգ�d��Unexceptx�motnZ������f��є�� O����� 90J�єS?P CSXC<�f���Ҟ� Py�We�}���PRI�>v�r�t�men�� ^��iPɰa��x���vGrid�play��v��0��)�H1�M-10�iA(B201 z�2\� 0\k/�_Ascii�l��8��ɐ/�Col��ԑoGuar� 
��� /P-�ޠ"K��s�t{Pat ��!�S�Cyc�҂�o�rie��IF8�ata- quҐ�� xƶ��mH574���RL��am���P~b�HMI De3�1(b����PCϺ�?Passwo+!��7"PE? Sp$�[����tp��� ven���Tw�N�p�YELLOW BOE	�k$Arc��vis���3*�n0Wel=dW�cial�7��V#t�Op����1�y� 2F�a�p�ortN�(�p�T1��T� �� ��xy�]�&TX��tw�i�gj�1� b� ct�\�JPN ARCPSU PR���oݲOL� Sup�2fil� &PAɰ�אcro�� "PaM(����O$SS� �eвtex�� r����=�t�ssaIgT��P��P@�0Ȱ�锱�rtW��8H'>r�dpn��nG1
t�!� z ���ascbin4Opsyn��+Aj��M HEL�NC�L VIS PKGS PLOA`��MB �,�4VW��RIPE GE�T_VAR FI�E 3\t��FL�[�OOL: AD�D R729.F_D \j8'�CsQ�QE��DVvQ�sQ�NO WTWTE|��}PD  �^�ѼbiRFOR ��E�CTn�`��ALS�E ALAfPCP�MO-130  �M" #h�D: �HANG FRO�MmP�AQfr��R�709 DRAM� AVAILCH�ECKSO!��sQV�PCS SU�@L?IMCHK Q +P~~dFF POS���F�Q R593�8-12 CH�ARY�0�PROG�RA W�SAV�EN`AME�P.SeV��7��$En*�p�p?FU�{�TRC|�� SHADV0UP?DAT KCJўR�STATI�`�P _MUCH y�1���IMQ MOTN�-003��}�RO�BOGUIDE DAUGH�a����*�tou����I� :Šhd�ATH�Pep�MOVET�ǔV�MXPACK M�AY ASSER�T�D��YCLfqT�A�rBE CORg vr*Q3rAN�p�RC OPTIO�NSJ1vr̐PS_H-171Z@x�tcǠSU1�1Hp^9R!�Q�`_T�P���'�j�d{tby �app wa 5I�~d�PHI���p�a�TEL�MXSPOD TB5bLu 1���UB6@�qENJ`C�E2�61��p��s>	�may n�0�� R6{�R� �Rt�raff)�� 4�0*�p��fr��s�ysvar sc�r J7��cj`DJU��bH V��Q�/�PSET ER9R`J` 68��P�NDANT SC�REEN UNR�EA��'�J`D�pP�A���pR`IO Y1���PFI�pB�p_GROUN�PD���G��R�P�QnRSVI�P !p�a�PDIGIT VERS�r�}BLo�UEWϕ �P06  �!��M�AGp�abZV�D�I�`� SSUE��ܰ�EPLAN� JOT` DEL��pݡ#Z�@D͐C�ALLOb�Q phx��R�QIPND���IMG�R719޺�MNT/�PES� �pVL�c��Ho�l�0Cq���tPG:t�`C�M�canΠ޹�pg.v�S: �3D mK�vie�w d�` �p��e�a7У�b� of ��Py���ANNOT� ACCESS �M��Ɓ*�t4s �a��lok��Fl�ex/:�Rw!m-o?�PA?�-������`n�pa SNB�PJ AUTO-��06f����TB��PI�ABLE1q 63}6��PLN: RG�$�pl;pNWFM�DB�VI���tWI�T 9x�0@o��Q�ui#0�ҺPN R;RS?pUSB�� �t & remo�v�@ )�_��&AxnEPFT_=� 7<`��pP:�OS-1w44 ��h s�g��@OST� � �CRASH DU{ 9��$P�p�W� .$��LOGIN��8&�J��6b�046 issu�e 6 Jg��:� Slow �s�t��c (Hos�`�c���`IL`IM�PRWtSPOT:�Wh:0�T�STYzW ./�VMGR��h�T0CAT��ho�s��E�q��� �O�S:+pRTU�' k�-S� ����E�:��pv@�2�� t�\hߐ��m ��a3ll��0�  $�H�� WA͐��3 C�NT0 T�� W�roU�alarm���0s�d � �0SE�1���r R{�OM�EBp���K� 55f��REàSEst��g     ��KANJI�no����INISIT�ALIZ-p�dn1w�eρ<��dr�� �lx`�SCII �L�fails �w�� ��`�YST�Ea���o��Pv� I�IH���1W�Gro�>Pm ol\wpS�h@�P��Ϡn c�flxL@АWRI �OF Lq��p?��F�up��de-�rela�d "kAPo SY�ch�A�betwe:0IN�D t0$gbDOȲ��r� `�Gi�gE�#opera�bilf  PAbH�i�H`��c�lead�\etf�Ps�r�OS 030�&: �fig��GLA �)P ��i��7Np �tpswx�B��If�g������5a}E�a EXCE#dxU�_�tPCLOS��o"rob�NTdp�FaU�c�!���P�NIO V750ªQ1��Qa��DB� ��P M�+P�QE�D�DET��-� �\rk��ONLI;NEhSBUGIQ �ߔĠi`Z�IB�S �apABC JA'RKYFq� ���0�MIL�`� R�pNrД �p0GAR���D*pR��P�"! 	jK�0cT�P�Hl#�n�a�ZE V�� �TASK�$VP2 (�4`
�!�$�P�`W�IBPK05�!F�ȐB/��BUSY� RUNN�� "��򁐈��R-p�L�O�N�DIVY�CsUL��fsfoaBW�p���300	V��ˠIT`�ao505.�@OF᠏UNEX�P1b�af�@�E��SVEM�G� NMLq� D�0pCC_SAFE�X 0c�08"qD �P�ET�`N@�#J8	7����RsP�A'��M�K�`K�H �GUNCHG۔M�ECH�pMc� T�  y, g@�$ �ORY LEAKpA�;�ޢSPEm�tJa��V�tGRIܱx�@�CTLN��TRk�FpepR�j5m0�EN-`IN�����p �`�Ǒk!���T3/dqo�STOR�0A�#�L�p �0�@�Q�АY�&�;p�b1TO8pP�s���F`B�@Yp`�`DU�B�aO�supk�t4 � 2P�F� Bnf�Q�P?SVGN-1��VN�SRSR)J�U�P�a2�Q�#D�q l� O��QBRKCTR5Ұ�|"-�r��<pc�j!INVP�D ZO� ��T`h#�Q<�cHset,|D��"DUAL� w�2�*BRVO117 A]�TNѫt�+bTa2473��q.?��s�AUz�i�B�com�plete��60�4.� -�`h�anc�U� F:��e8��  ��np�JtPd!q��`��� �5h596p�!5 d�� "p�P�P�Q�0�P�2�p�A� xP��R(T}\xPe� aʰI���E��1��p� j�  � �xSP�^P� �A�AxP�q 5 s�ig��a��"AC�;a��
�bCexPb;_p��.pc]l<b�Hbcb_circ~h<n�`tl1�~`xP�`o�dxP�b]o2�� cb�c�ixP�jup�frm�dxP�o�`e�xe�a�oFdxPtp�ed}o��u`�cpt�libxzxP�lcr �xrxP\�blsazEdxP_fm�}gcxP��x���o|sp�o�mc�(��ob_jzop��u6�wf��t��wm2s�1q��sld�)���jmc�o\�n��nuhЕ��|st�e��>�cpl�qp�iwck���uvf0uߒ��l�visn�Cgac�ulwQ
E F w ! Fc.fd�Q�v�� qw���Da�ta Acqui�si��nF�|1�RR�631`��TR�QD�MCM �2�P7u5H�1�P583xPm1��71��59`�5�P57<PxP�Q�����(���Q��o ypxP!daq\�1oA��@�� ge/��etdms�"DM�ER"؟,�pgdD���.�m���-��q�aq.<᡾xPmo���h���f{�u�`13���MACROs,7 Sksaff�@z����03�SR�Q(��Q6��1�Q9ӡ�R�Z�Sh��PxPJ643��@7ؠ6�P�@�PRS�@���e �Q�UС� PIK�Q52 �PTLC�W��xP3; (��p/O��!��Pn �xP5��0�3\sfmnmc? "MNMCq�<�ԔQ��\$AcX�FM ���ci,Ҥ�X���װcdpq+�
�sk�S�K�xP�SH560�,P��,�y�ref?p "REFp�d��A�jxP	�of�O�Fc�<gy�to�T�O_����ٺ����+je�u��caxCis2�xPE�\�e�q"ISDTc��]��prax ��MN���u�b�isde�܃h�\�w�xP! i�sbasic��B�� P]��QAxes�R6������.��(Ba�Q�ess ��xP���2�D�@�z�atis���(�@{�����~��m��FMc�u�{�
ѩ�MNIS��ݝ����x�������ٺ��x� j�75��Devic��� Interf�ac�RȔQJ75a4��� xP�Ne` ��xP�ϐ2�б�����dn� "DN�E���
tpdnui5UI��ݝ	�bd�bP�q_r�sofOb
dv_aro��u��|���stchkc���z	 �(}on1l��G!ffL+H��J(��"l"/�n��b��z�hamp���T�C�!i�a"�5�9��S�q��0 (��+P�o�u�!2��xp}c_2pcchm�ЏCHMP_�|8бp�evws��2쳌p�csF��#C Se=nxPacro�U���-�R6�Pd�xPk�����p��gT�L��1d M�2`��8�1c4�ԡ�3 qem��G�EM,\i(��Dgesnd�5���H{�}H�a�@sy���c�Is1u�xD��Fmd��I���7�4���u���AccuCal�P�4� ���ɢ7ޠB0��6j+6f�6��99\aFF q�S(�U��2�
�X�p�!Bd��cb�_�SaUL��  ��� ?�ܖto��o�tplus\tsCrnغ�qb�Wp���t���1��Tool� (N. A.)0�[K�7�Z�(P�m� ���bfcls� k94�"K4p��q�tpap� "P�S9H�stpsw�o��p�L7��t\ �q����D�yt5�4�q���w�q��� �M�uk��rkey����s���}t�sfeatu6�EA��� cf)t�\Xq�����d�h5���LRC0�md��!�587���aR�( ����2V��8c?u3l\�pa3}H�&r-�Xu���t,�� �q "�q�Ot��~,����{�/��1c�}����y �p�r��5���S�XA�g�-�y���Wj87�4�- iRViys���Queu� � Ƒ�-�6�1���	(����u���tӑ�����
�tpvtsn "VTSN�3�C�+�� v\pRDVx����*�prdq\�yQ�&�vstk=P0������nm&_����clrqν���get�TX��Bd��aoQϿ�0qst!r�D[� ��t�p'Z�����npv��@�enlIP0��D!x�'��|���sc ߸��tvo/��2�q���vb����q���!����h]��(� Co�ntrol�PR�AX�P5��556l�A@59�P56.@�56@5A�J6�9$@982 J552 IDVR7� hqA���16�H���La�� ��Xe��frlparm.�f�FRL�am0��C9�@(F�����w6{���A��QJg643�� 50�0�LSE
_pVA�R $SGSYS�C��RS_UNITS �P�2�4tA��TX.$VNUM?_OLD 5�1�xP{�50+�"�`? Funct���5@tA� }��`#@�`3�a0�cڂ��9���@�H5נ� �P���( �A����۶}����0ֻ}��bPRb�߶�~ppr4�TPSP`I�3�}�r�10�#@;A� t�
`���1����96�����%C��� Aف��J�bIncr�	����\���1�o5qni4�MNINp	xP�`���!���Hour  �� 2�2�1 �AAV1M���0 ���TUP ��J�545 ��61�62�VCAM�  (�CL�IO ��R6x�N2�MSC �"P �ST�YL�C�28~ 1�3\�NRE "�FHRM SCH~^�DCSU%�ORSR {b�0�4 �EIO�C�1 j 542� � os| � egist������7�1�MA�SK�934"7 <��OCO ��"%3�8��2����� 0 HB��� 4v�"39N� Re��� �LCHK
%O�PLG%��3"%M7HCR.%MC  ; �4? ��6 dPI��54�s� DSW�%MD� pQ�K!6C37�0�0p"�1��֠"4 �6<27 �CTN K � 5 J���"7��<25�%z/�T�%FRDM� �Sg!��9309 FB( NBA�P� �( HLB  Me�n�SM$@jB( PgVC ��20v�α2HTC�C�TMIL��\@PA�C 16U�hAJ`S9AI \@ELN��<2�9s�UECKy �b�@FRM �b��OR���IPL���Rk0CSXC \���VVFnaTg@�HTTP �!2�6 ��G�@ob�IGUI"%IP�GS�r� H863� qb�!�07r�!34� �r�84 \s`o`! Qx`CC3 Fbr�21�!96 rb�!51 ���!53R% 1!s3!��~��.p"9js VATFUJ775"��pLRu6^RP�WSMjU'CTO�@xT58 F�!80���1XY <ta3!770 ��7885�UOL  GT�So
�{` LCM9 �r| TSS�EfP�6 W�\@CPE `��0VR� l�Q�NL"��@001 oimrb�c3 =�`�b�0���0�`6 w�b-P- R-�b8nn@5EW�b9 �Ҁ�a� ���b�`ׁ�b2� 2000��`3$��`4*5�`5!�c��#$�`7.%�`8 oh605? U0�@�B6E"aRp7� !Pr8 t�a@�>tr2 iB/�1vp�3�vp5 Ȃtr9�Σ�a4@-p�r3 F��r5&�re`Lu��r7 ��r8�U��p9 \h738|�a�R2D7"�)1f��2&�7� �O3 7iC��4>wq5Ip�Or60 CҲL�1bEN�4 I�p�yL�uP��@N�-PJ�8�N�8NeN�9 PH�r`�E�b7]��|���8�Вࠂ9 �2��a`0�qЂ5~�%U097 0��@1�0���1 (<�q�3 5R��� �0���mpU��0�0�7*�H@(q�\P�"RB6�q124��b;��@���@06l� x�3 pB/x��u ��x�6 H60�6�a1� ��7 �6 ���p�b1�55 ����7jUU�162 �3 �g��4*�65 2�e "_��P�4U1H`���B1���`0'�174 �q��P�E?186 R ��P��7 ��P�8&�3 }(�90 B/�s�191����@202��6 3���A��RU2� d��2 �b2h`��4�᪂2��4���19v Q�2T��u2d�Tpt2� ���H�a2hP�$�5����!U2�p�p
�2�p��@5�0-@��i8 @�9��TX@�t� �e5�`rb26Af�2^R�a�2Kp��1Dy�b5Hp�`
�5��0@�gqGA���a52hѐ�Ḳ6�60ہ)5� ׁ2��8�E��M9�EU5@ٰ\�qQ5hQ`S�2ޖ5�p\w�۲�pJ �-P��M5�p1\t�H�4���PCH�7j��phi�w�@��P�x��559 ldu� P�D��@�Q�@������� �`�.��P>��8�58�1�"�q58�!AM�۲T�A iC�a5�89��@�x����5 �a��12׀0.�1���,�2����,�!P'\h8��Lp ��,��7��6�0840\���ANRS 0C�}A��p��{��ran��FRA��Д� �е���A%���ѹ� �Ҍ�����(����� ����З�������� �ь����$�G��1�Čը���������� xS�`q� c �����`64���M��iC/50T-H������*��)p46��� C��N�����m75s֐� 1Sp��b46��v�x���ГM-71?�a7�З����42������C��-�а�7�0�r�E��/h ����O$��rD���c7c7C�q�䈌Ѕ���L��/��2\imm7c7�@g������`��� (��e�����"�������a r��c�T	,�Ѿ�"��,�� ���x�Ex�m77t ����k���5������)�iC��-HS -� B
_�>���+�Т�7U�]���TMh7�s��7�������-9?�/260L_������Q�������]�9pA/@���q�S�х���h�621��c��92�������.�)92c0�g$�@������)$��5$���pylH"O"
�21���t?�350�����p��$�
�� �350!���0��9��U/0\m9��M9�A3��4%� s"��3M$��X%u���"him98J3����� i d�"m4~�10�3p�� ����h79!4̂�&R���H�0�� ��\���g�5AU��� ���0���*2��00��#06�АՃ�,�է!07{r ��� �����kЙ@����EP�#�������?��#!�;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/�p�?�ҽCD25L�����0�"l�2�BL
#��B��\20 �2_�r�re���X���1��N����A@��z��`C�pU��`F��04��DyA�\�`fQ��sU����\�5  ���; p�^P��<$�85���+P=�ab;1l��1LT��lA8�!uDnE(�2�0T��J�1 e�bHC85���b�Ռ�5[�16Bs���������d2��x��m6t!`Q����bˀ��8�b#�(�6iB;S�p �!��3� ��b�s ��-`�_�W8�_�L���6I	$�X5�1��U85��R�p6S ����/�/+q�!�q��`�6o��5m[o)�m6sW��Q�?��set06p ��3%H�5��10p$�����g/�JrH���  ��A�85!6����F�� ���p/2��h�܅�✐)�5��̑v��(�&�m6��Y�H�ѝD̑m�6�Ҝ��a6�DM����-S�+��H2�����Ҽ�� �r ̑��✐��l���p1���F���2��\t6h T6H ����Ҝ�'Vl�� �ᜐ�V7ᜐ/����
;3A7��p~S��������4�`圐�V����!3��2�PM�[��%ܖO�chn��vel5����Vq���_arp#��̑��.���2l_hempq$�.�'�6415� ��5���?����F�����5g�L�ј[���!1��𙋹1����M7NU�М��e(ʾ����uq$D;��B-�4��3&H�f�c�� ��h������u� ��㜐��ZS�!ܑL4���M-����S�$ ̑�ք �� 0��<�p����07shJ�H�v�À�sF��S*� ������̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(U L�&�(�,���0�\�?����̑�a�� xSP���a�e�w��2��(�	�2�C��A/���\�+p������21 (ܱ�CL S����B̺��7FГ��?�<�lơ1L@����c� ���u9�0����e/q��O���q9�K��r9 (�� ,�Rs�ז�5�G�m20c��i��w�2��:�0`�$��2 �2l�0�k�X�S� ,�Bι2��O���1!�41w���2T@� _std��G�y� ��x��H� jdgm�� ��w0\� �1L���	� P�~�W*�b��t �5������3�,���E{�������L��5\L��3 �L�|#~���~!���4�#��O����h�LA6A�������2�����44�����>[6\j4s��·����#��ol�E"w�8 Pk�����?0xj�H1��1Rr�>��]�2aF�2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l���0�&�"��|�`Am1��2��ػ��3�HqB ��K�R��ˑb� W���Fs���)�ѐ�@!���a�1����5��;16�16C��xC����0\imBQ@��d����b��\B5�-���DiL���O� _�<ѠPEtL�E�R�H�ZǠPgω�am1l��u���̑�b�<����<�$�T�̑�F ����Ȋ�Dpb��X�"��hr��p� .���^P��9�0\�� j971\kc/krcfJ�F�s������c��e "CTME�r���ɛ��a�`main.[��g��`run}�_vc �#0�w�1Oܕ_u��<��bctme��Ӧx�`ܑ�j735��- KAREL /Use {�U���AJ��1���p� Ȗ�9�B@��L�9���7j[�atk208 "K��Kя�
�\��9��a��̹8����cKRC�a�o ��kc�qJ�&s�� ���Grſ�fsD��:`y��s�ˑ1X\j|�&�rdtB�, ��`.v�q�� �sǑIf\�Wfj52�TKQuto Set���J� H5K53M6(�932���91�K58(�9�BA�1(��74O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v����! conre�;a#�Contro�l Re�ble��CNRE(�T�<р4�2���D�)���S�5�52��q(g�� (�򭂯4X�cOux�\�sfuts�UTAS`�i�栜���t�棂��? 6�T�!�GSA OO+D6� ��������,!���6c+� igt�t6�i��I0�TW8` ���la��vo58�o��bFå򬡯i�Xh���!Xk�0Y!8\m;6e�!6EC���v��6���������B<16�A���A�6s� ���U�g�T|ώ����r1�qR��˔Z4 �T�����,#�eZp)g����<ONO0���uJ��tCR;��F�a�� xSP�f��pr?dsuchk �1"��2&&?���t��*D%$�r(�✑�娟:r��'�s�qO��<�scrc�C�\At�trldJ"o�\��V����Paylo>�nfirm�l�!�87��7��A�3ad�! �?ވIЯ?plQ��3��3"0�q��x pl�`��p�d7��l�calC��uDu���;��mo�v�����initX�:s8O��a�r4 ���r67A4|�e �Generati�ڲ���7g2q$��g{ R� (Sh��$�c ,|�bE��$Ԃ�\�:�"��4b��4�4�. sg��A5�F$d6"e;Qp "SHAP��TQ ngcr pG�C�a(�&"� ��"gGDA¶��r6��"aW�/�$dat�aX:s�"tpadx��[q�%tput;a __O7;a�o8�1�yl+s�r�?�:�#�?�5Ix�?�:c O�:y O��:�IO�s`O%g �qǒ�?�@0\��"o��j92;!�Ppl.�Collis�QSkip#��@5��@J� �D��@\ވ�C@XJ�7��7�|s2���ptcls�LS��DU�k?�\_ ects�`�< \�Q ��@���`dcKqQ�FC;��J,�n��`# (��4eN����T�{���'j(�c �����/IӸaȁ��̠�H�����зa��e\mcclm?t "CLM�/�¾� mate\��lmpALM�?>p�7qmc?����2vm��q��%�3s��_svx90�_x_msu�2�L^v_� K�o�{i�n�8(3r<�c_l�ogr��rtr)cW� �v_3��~yc��d�<�te���der$cCeN� Fiρ�R���Q�?�l�ent�er߄|��(Sd���1�TX�+fK�r�a99sQ9+�5��r\tq\� "F�NDR����STDn$LA�NG�Pgui��D�⠓�S������sp�!ğ֙uf�ҝ�s ����$�����e+�=� ��������������<w�H�r\fn_�ϣ���$`x�tcpma>��- TCP���~��R638 R�X�Ҡ��38��M7p,���Ӡ�$Ӡ�8p0а��VS,�>�tk��99�a��B3���PզԠ`��D�2�����UI�� t���hqB���8�����0���p���re�ȿ��exe@4φ�B�ࠓe38�ԡG�rmp8WXφ�var@�π��3N�����vx�!�ҡ��q�RBT� $cOPTN? ask E0�Ӿ1�R MAS0�H�593/�96 HY50�i�480�5�!H0��m�Q�K��7�
0�g�Pl�h0ԧ�<2�ORDP��@"���t\mas��0��a��"�ԧ�����k@�գR����ӹ`m�՘b��7�.f��u�d���r��spla�yD�E���1w�UP�DT Ub��887� (��Di{���v �Ӛ�Ԛ⧔��#�B���㟳��o  �@���a�䣣��60q���B����qscaan��B���ad@�������q`�䗣��#��К�`2�� vlv��Ù�$�>�b����! S��Ea�sy/К�Util���룙�511 JȘ����R7 ��No�r֠��inc),(<6Q�� �`c��"84�[���986FVR�x So����q�nd6����P��4�a\ �(��
  �������d���K�bdZ���meyn7���- Me`CtyFњ�Fb�0�8TUa�577?Ai3R��\�5�u?��!� n���f�x�����l\mh����űE|hmn�	��<\O����e�1�� l!��y(��Ù�\|p����0�B���Ћmh�@�� :.aG!���/� t�55�6�!X�l�.�us��Y/k)ensSubL���eK�h��  �B\1;5g?y?�?0�?D��?*rm�p�?Ktbox O2K|`?�G��C?A%ds���?1ӛ#� �TR�� /��P�4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R�?Ă�Q3t.�P׀a�l��P+OP517��IN0a��Qq(}g��PESTf3ua�PB�l�ig�h��6�aq��P �� xS��`  <n�0mbumpP�Q7969g�69�Qq���P0�baAp�@Q�� BOX��,>vc�he�s�>vetux㒣=wffse�3���]�;u`aW��F:zol�sm<ub�a0-��]D�K�ibQ�c�ெ�Q<twaǂ tp��Q҄Taror �Recov�b�O�P�642����a`�q��a⁠QErǃ��Qry�з`�P'�T �`�aar������	{'��pak971��7�1��m���>�pj�ot��PXc��C�1�a�db -�ail��n�ag���b�QR62�9�a�Q��b�P  �
  �P���$$CL[q �����������$�PS_D�IGIT���"�!�4�F�X� j�|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� �������*璬1:PRO�DUCT�Q0\P/GSTK�bV,n�99�\����$FEAT_�INDEX��~�?� 搠�ILECOMP +;��)��"���SETUP2 �<����  N !�_A�P2BCK 1=~�  �)}D6/E+%,/i/�� W/�/~+/�/O/�/s/ �/?�/>?�/b?t?? �?'?�?�?]?�?�?O (O�?LO�?pO�?}O�O 5O�OYO�O _�O$_�O H_Z_�O~__�_�_C_ �_g_�_�_	o2o�_Vo �_zo�oo�o?o�o�o uo
�o.@�od�o ���M�q� ��<��`�r���� %���̏[������� !�J�ُn�������3� ȟW������"���F� X��|����/���֯ e������0���T�� x������=�ҿ�s� ϗ�,ϻ�9�b�� �P/ 2) *�.VRiϳ�!�*�����������P�C�7�!�FR6�:"�c��χ��T ��߽�Lը��ܮx�<��*.F��>�" �	N�,�k��ߏ��STM ������Qа���!�iP�endant POanel���H��F���4������GIF�������u����JPG&P���<����	PANEL1.DT��������2�Y�G��
3w�����//�
4�a/�O//�/�/�
TPEI?NS.XML�/����\�/�/�!Cu�stom Too�lbar?�PASSWORD/~�FRS:\R?�? %Pass�word Config�?��?k?�? OH�6O�?ZOlO�?�O O�O�OUO�OyO_�O �OD_�Oh_�Oa_�_-_ �_Q_�_�_�_o�_@o Ro�_voo�o)o;o�o _o�o�o�o*�oN�o r��7��m ��&���\���� �y���E�ڏi���� ��4�ÏX�j������ ��A�S��w����� B�џf�������+��� O���������>�ͯ ߯t����'���ο]� 򿁿�(Ϸ�L�ۿp� ��Ϧ�5���Y�k� � ��$߳��Z���~�� �ߴ�C���g����� 2���V����ߌ��� ?����u�
���.�@� ��d������)���M� ��q�����<��5 r�%��[� &�J�n� �3�W��� "/�F/X/�|//�/ �/A/�/e/�/�/�/0? �/T?�/M?�??�?=? �?�?s?O�?,O>O�? bO�?�OO'O�OKO�O oO�O_�O:_�O^_p_ �O�_#_�_�_Y_�_}_�o�_�_Ho)f�$F�ILE_DGBCK 1=��5`��� �( �)
SUMMARY.DGRo��\MD:�o�o�
`Diag S?ummary�o�Z�
CONSLOG��o�o�a
J�aC�onsole l�ogK�[�`ME?MCHECK@'��o�^qMemory Data���W�)�qHADOW���P���sShadow� Changes�S�-c-��)	FTP=��9����w�`qmment �TBD׏�W0<��)ETHERNET̏�^�q�Z��a�Etherne�t bpfiguration[��P��?DCSVRFˏ���Ïܟ�q%�� �verify a�llߟ-c1PY���DIFFԟ��̟�a��p%��diCffc���q��1X�8?�Q�� �����X��CHGD ��¯ԯi��px���� ���2`�G�Y��c ��� �GD��ʿܿq��p���Ϥ��FY3h�O�a���c ��(�GD������y��p�ϡ�0��UPDATES�.�Ц��[FRS�:\�����aUp�dates Li�st���kPSRB?WLD.CM.��\���B��_pPS_ROBOWEL�� �_����o��,o!�3� ��W���{�
�t���@� ��d�����/��S e�����N� r� =�a� r�&�J��� /�9/K/�o/��/ "/�/�/X/�/|/�/#? �/G?�/k?}??�?0? �?�?f?�?�?O�?O UO�?yOO�O�O>O�O bO�O	_�O-_�OQ_c_ �O�__�_:_�_�_p_ o�_o;o�__o�_�o �o$o�oHo�o�o~o �o7�o0m�o�  ��V�z�!�� E��i�{�
���.�Ï R����������.�S� �w������<�џ`� �����+���O�ޟH� �����8���߯n�����$FILE_���PR����������� �MDONLY �1=4�� 
 ���w�į��诨� ѿ�������+Ϻ�O� ޿sυ�ϩ�8����� n�ߒ�'߶�4�]��� ��ߥ߷�F���j��� ��5���Y�k��ߏ� ��B�����x���� 1�C���g������,� ��P���������?���Lu�VISB�CKR�<�a�*.�VD|�4 FR�:\��4 V�ision VD file� : LbpZ�#�� Y�}/$/�H/� l/�/�/1/�/�/�/ �/�/ ?�/1?V?�/z? 	?�?�???�?c?�?�? �?.O�?ROdOO�OO �O;O�O�OqO_�O*_ <_�O`_�O�__%_�_��MR_GRP �1>4�L�UC�4  B�P	 �]�ol`�*�u���RH�B ��2 ���� ��� ���He�Y�Q`orkbIh��oJd�o�Sc�o�o�L,�MVS��K?�F�5U�aS��i�o�o� E=aEP���E!�-����9?6">_�Z`}@6�A��a$lq?_���A�\�xq0~�� F@ �r�d�a�}J��NJk��H9�Hu���F!��IP��s}?�`�.9��<9�8�96C'6<?,6\b�1�@,.�g�R���v�A�PA�����|�ݏx�� �%��I�4�F��j� ����ǟ���֟��!�`�E�`r�UBH�P �~�������W�
6�PJ��PQØ�˯�o�oB�x�P5���@�33@����4�m�T�UUU�U�~w�>u.�?!x�^��ֿ����3��=[z��=�̽=V6�<�=�=��=$q��~��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�Ϡ Cϫo��C�
�P��P'�6��_V�  m�o��To��xo�ߜo ������A�,�e�P� b���������� ���=�(�a�L���p� ���������������� *��N9r]�� ������8 #\nY�}�� �����/ԭ//A/ �e/P/�/p/�/�/�/ �/�/?�/+??;?a? L?�?p?�?�?�?�?�? �?�?'OOKO6OoO�O HߢOl��ߐߢ��O��  _��G_bOk_V_�_z_ �_�_�_�_�_o�_1o oUo@oyodovo�o�o �o�o�o�oN u����� ����;�&�_�J� ��n�������ݏȏ� �%�7�I�[�"/�� ������ٟ������� 3��W�B�{�f����� ��կ�������A� ,�e�P�b��������O �O�O��O�OL�_ p�:_�����Ϧ����� ���'��7�]�H߁� lߥߐ��ߴ������� #��G�2�k�2��V w�����������1� �U�@�R���v����� ��������-Q �u���r��6 ��)M4q \n������ /�#/I/4/m/X/�/ |/�/�/�/�/�/?ֿ �B?�f?0�BϜ?f� �?���/�?�?�?/OO SO>OwObO�O�O�O�O �O�O�O__=_(_a_ L_^_�_�_�_���_�� o�_o9o$o]oHo�o lo�o�o�o�o�o�o�o #G2kV{� h������� C�.�g�y�`������� ���Џ���?�*� c�N���r�������� ̟��)��M�_�&? H?���?���?�?�?�� ��?@�I�4�m�X�j� ����ǿ���ֿ��� �E�0�i�Tύ�xϱ� ����������_,��_ S���w�b߇߭ߘ��� ��������=�(�:� s�^��������� ��'�9� �]�o��� ��~����������� ��5 YDV�z ������1 U@yd��v� ����/Я*/��
/ �u/��/�/�/�/�/ �/�/??;?&?_?J? �?n?�?�?�?�?�?O �?%OOIO4O"�|OBO �O>O�O�O�O�O�O!_ _E_0_i_T_�_x_�_ �_�_�_�_o�_/o�� ?oeowo�oP��oo�o �o�o�o+=$a L�p����� ��'��K�6�o�Z� �����ɏ��폴�  ��D�/ /z�D/�� h/ş���ԟ���1� �U�@�R���v����� ӯ������-��Q� <�u�`���`O�O�O�� �޿��;�&�_�J� oϕπϹϤ������ ��%��"�[�F��Fo �ߵ����ߠo��d�!� ��W�>�{�b��� ������������A� ,�>�w�b����������������=���$FNO ����\_�
F0l q � FLAG>�(�RRM_CHKT_YP  ] ���d �] ��O=M� _MIN� 	����� �  �XT SSB_CF�G ?\ �����OTP_DEF_OW  	���,IRCOM�� >�$GENO�VRD_DO���<�lTHR� �d�dq_ENB�] qRAVC_GRP 1@�I X(/ %/ 7//[/B//�/x/�/ �/�/�/�/?�/3?? C?i?P?�?t?�?�?�? �?�?OOOAO(OeOpLO^O�OoROU��F\� ��,�B,�8�?����O�O�O	__  D�UPE_�Hy_�\@@m_B�=�vR/���I�O�SMT�G
���
�oo+l�$HOSTC�s1H�I� ���zMSM�l[�bo�	127�.0�`1�o  e�o�o�o#z�o�FXj|�l60s	�anonymou�s������Q%ao�&�&��o �x��o������ҏ� 3��,�>�a�O�� ��������Ο�U%�7� I��]����f�x��� �����ү����+� i�{�P�b�t������ ������S�(�:� L�^ϭ�oϔϦϸ��� ���=��$�6�H�Z� ����Ϳs�������� ��� �2���V�h�z� ��߰���������
� �k�}ߏߡߣ���� ����������C�* <Nq�_���� ��-�?�Q�c�eJ ��n����� ��/"/E�X/j/ |/�/�/�%'/ ?[0?B?T?f?x?� �?�?�?�?�??E/W/�,O>OPObO�KDaEN�T 1I�K P�!�?�O  �P �O�O�O�O�O#_�OG_ 
_S_._|_�_d_�_�_ �_�_o�_1o�_ogo *o�oNo�oro�o�o�o 	�o-�oQu8 n������� �#��L�q�4���X� ��|�ݏ���ď֏7����[���B�QUICC0��h�z�۟���1ܟ��ʟ+���2�,���{�!ROUTER|�X�j�˯!PCJOG̯���!192.�168.0.10���}GNAME �!�J!ROBO�T�vNS_CFG� 1H�I ��Auto-started�$/FTP�/���/ �?޿#?��&�8�J� �?nπϒϤ�ǿ��[�������"�4�G�#� ��������������� �������&�8�J�\� n����������� ��/�/�/F���j��� �������������� 0S�T��x�� ���!�3��G, {�Pbt��C� ���/�:/L/ ^/p/�/���	/ �/=?$?6?H?Z?)/ ~?�?�?�?�/�?k?�? O O2ODO�/�/�/�/ �?�O�/�O�O�O
__ �?@_R_d_v_�_�O-_ �_�_�_�_oUOgOyO �O�_ro�O�o�o�o�o �o�_&8Jmo �o�����o)o ;oMoO!��oX�j�|� ����oď֏���� /���B�T�f�x���^��ST_ERR �J;�����PDUS_IZ  ��^P�����>ٕWRD� ?z��� � guest���+�=�O�a�s��*�SCDMNGR�P 2Kz�Ð��۠\���K�� 	P01�.14 8�q �  y��B�    ;�����{ ���߇������������������~ �ǟI�4�m��X�|��  �i  �  
����� ����+��������
����l�.x����"�l�ڲ۰�s�d�������_�GROU��L��� ��	��۠07�K�QUPD  d���PČ�TYg������TTP_AUTH 1M��� <!iPeOndan���<��_�!KARE�L:*�����K�C%�5�G��VI�SION SETZ���|��Ҽߪ� ��������
�W�.��@��d�v���CTRL N��������
�FFF9�E3���FRS�:DEFAULT��FANUC� Web Server�
���� ��q��������������WR_CONFI�G O�� ����IDL_CP�U_PC"��B���= �BH#M�IN.�BGNR_IO��� ���% �NPT_SIM_�DOs}TPM�ODNTOLs >�_PRTY�=�!OLNK 1P���'9K�]o�MASTE�r �����O_CFG��UO����CYCLE���_ASG 1Q���
 q2/D/V/ h/z/�/�/�/�/�/�/��/
??y"NUM����Q�IPC�H��£RTRY�_CN"�u���SGCRN������1 ���R�����?��$J23_�DSP_EN������0OBPROqC�3��JOGV��1S_�@��8G�?�';ZO'??0C�POSREO�KANJI_�ϠuH�A#��3T ���E<�O�ECL_LM B2�e?�@EYLOGG+IN��������LANGUAGE� _�=� ,}Q��LG�2U���+�� �x�����P�C � �'0������MC:\�RSCH\00\�˝LN_DISP V������f�TOC�4Dz\�=#�Q�?PBOOK W+��o���o�o���Xi�o�o �o�o�o~}	x(y��	ne�i�ek�ElG_BUFF K1X���}2� ���Ӣ����� �'�T�K�]������� ����ɏۏ���#��P��ËqDCS }Zxm =���%| d1h`���ʟܟ�g��IO 1[+ �?'����'�7�I� [�o��������ǯٯ ����!�3�G�W�i��{�������ÿ׿�E^l TM  ��d�� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߈t��SEV�0m�TYP�� ��$�}�ARS"�(_�s�2�FL 1\��0�������������L�5�TP<P���}DmNGNAM�4��U�f�UPS`G�I�5�A�5s�_L�OAD@G %�j%@_MOV��u����MAXUALRMB7�P8��y���3�0]&q��Ca]s�3�~�� 8@�=@^+ طv	V��V0+�P�A�5d�r���U������ E(iTy��� ����/ /A/,/ Q/w/b/�/~/�/�/�/ �/�/??)?O?:?s? V?�?�?�?�?�?�?�? O'OOKO.OoOZOlO �O�O�O�O�O�O�O#_ _G_2_D_}_`_�_�_ �_�_�_�_�_o
oo Uo8oyodo�o�o�o�o��o�o�o�o-��D_LDXDISA^��� �MEMO_A�PX�E ?��
 �0y�����������IS�C 1_�� � O����W�i��� ��Ə�����}��ߏ D�/�h�z�a������ ��������@��� O�a�5���������� ��u��ׯ<�'�`�r� Y������y�޿�ۿ ���8Ϲ�G�Y�-ϒ� }϶ϝ�����m������4��X�j�#�_MS�TR `��}�S_CD 1as}�R� ��N��������8�#� 5�n�Y��}����� �������4��X�C� |�g������������� ��	B-Rxc ������� >)bM�q� ����/�(// L/7/p/[/m/�/�/�/ �/�/�/?�/"?H?3? l?W?�?{?�?�?�?n��MKCFG b���?��LTAR�M_�2cRuB �3WpTNBp�METPUOp�2�����NDSP_CMNTnE@F�EN�� d���N�2�A�O�D�EPOSC�F�G�NPSTOoL 1e-�4@�<#�
;Q�1;UK_ YW7_Y_[_m_�_�_�_ �_�_�_o�_oQo3o�Eo�oio{o�o�a�AS�ING_CHK � �MAqODAQ�2CfO�7J�eDE�V 	Rz	M�C:'|HSIZE�n@����eTASK� %<z%$12�3456789 ���u�gTRIG �1g�� l<u% ���3���>svv�YPaq��kEM_�INF 1h9G� `)�AT&FV0E0�(���)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ���ڄH������G�ֈAO�w�2�������џ �������� ͏ߏP��t������� ]�ί�����(�۟ �^��#�5�����k� ܿ� ϻ�ů6��Z� A�~ϐ�C���g�y��� �����2�i�C�h�� ��G߰��ߩ��ߙϫ� �������d�v�)ߚ� �߾�y�������� <�N��r�%�7�I�[� �����9�&��J�[�g��>ON�ITOR�@G ?�;{   	EOXEC1�3�2�3�4�5��p�U7�8�9�3� n�R�R�RR RR(R4RP@RLR2Y2eU2q2}2�2�U2�2�2�2��3Y3e3��aR�_GRP_SV �1it��q(�5�{
��5��۵MO~q_DCd~�1�PL_NAME �!<u� �!�Default �Personal�ity (fro�m FD) �4R�R2k! 1j)T?EX)TH��!�AX d�?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O�Ox2-?�O�O�O_�_0_B_T_f_x_�b< �O�_�_�_�_�_�_o@ o2oDoVoho&xRj"g 1o�)&0\�bO, �9��b�a� @D�  �a?���c�a?�`�a�aA�'�6�ew;��	l�b	 �xJp���`�`	p �<� �(p� ��.r� K�K ���K=*�J����J���JV���kq`q�P��x�|� @j�@wT;f�r�f�qx�acrs�I�� ��p���p�r�ph}��3��´  ��>��ph�`z��꜖"g�Jm�q� H��N��ac��$�dw�� � �  P� Q� �� |  �а�m�Əi}	'�� � �I�� �  �����:�È���=���(��#�a�	���I  �n @H�i~�ab��Ӌ�b�$w���"N<0��  'Ж�q��p@2��@�����r�q5�C�pC>0C�@ C��z��`
�A1�]w@B�V~X�
nwB0h�A��p�ӊa�p@����aDz����֏���Я	�pv��( �� -��I��-�=��A&�a�we_q�`�p� �?�ff ���m��� �����Ƽ�!@ݿ�>N1�  P�apv(�` ţ� �=�qst��/?���`x`�� �<
6b<߈�;܍�<�ê�<� <�&P�ό�AO��c1��ƾ��?fff?O�?y&��qt@�.���J<?�`�� wi4����dly�e߾g ;ߪ�t��p�[ߔ�� �ߣ����� ����6�wh�F0%�r�!�߷�1ى����E��� E�O�G+� F�!���/���?�e�P���t���lyBL�cB��Enw4��� ����+��R��s���������h�Ô�>��I�mXj�F��A�y�weC�p�������#/�*/c/N/wi�����fv/C�`� CHs/�`
=$�p�<!�!������'�3A�A��AR1AO�^?�$�?����±
=ç>�����3�W
�=�#�]�;e���?�����{����<�>�(�B�u�����=B0�������	R��zH��F�G���G���H�U`E���C�+��}�I#�I���HD�F���E��RC�j=��>
I��@�H�!H�( E<YD0w/ O*OONO9OrO]O�O �O�O�O�O�O�O_�O 8_#_\_G_�_�_}_�_ �_�_�_�_�_"ooo XoCo|ogo�o�o�o�o �o�o�o	B-f Q�u����� ��,��P�b�M��� q�����Ώ���ݏ� (��L�7�p�[���� ��ʟ���ٟ���6�@!�Z�E�W���#1( �g��9�K���ĥ �����Ư!�3�8���!4�Mgs��,�IB�+8�J��a���{�d�d�����ȿP���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ�����X�����  %�� � �h�Vߌ�z߰�&�g�@/9�$�������7�����A�S�e�w�  ��������������2 F�$N�&Gb������X���!C���@���8�����F� �DzN�� F�P D�������)#B�'9K]o~#?���@@v
�4$8�8��:8�.
 v� ��!3EWi�{����:� ���ۨ�1���$MSKCFMA�P  ��� ���(.��ONREL  ��!9��E�XCFENBE'
8#7%^!FNCe/W$�JOGOVLIM�E'dO S"d�KE�YE'�%�RU�N�,�%�SFSPDTY0g&P%�9#SIGNE/W$TO1MOT�/T!��_CE_GRP [1p��#\x� �?p��?�?�?�?�? O�?OBO�?fOO[O �OSO�O�O�O�O�O_ ,_�OP__I_�_=_�_ �_�_�_�_oo�_:o��TCOM_C_FG 1q	-��vo�o�o
Va_AR�C_b"�p)UA�P_CPL�ot$N�OCHECK ?=	+ �x� %7I[m� �������!��.+NO_WAITc_L 7%S2NT^a�r	+�s�_E�RR_12s	)9��� ,ȍޏ��x����&��dT_MO���t��, /��*oq�9�PARAM:��u	+��a��ß'g{�� =?�3�45678901 ��,��K�]�9�i��������ɯۯ��&g������C��cUM_RSPACE/��|����$ODR�DSP�c#6p(OF�FSET_CAR9T�o��DISƿ���PEN_FILE�尨!�ai��`OPT?ION_IO�/���PWORK ve7s# ��V������p�4�p�	 ����p��<���R�G_DSBL  ���P#��ϸ�R�IENTTOD �?�C�� !=#���UT_SIM_ED$�"���V��?LCT w}�h��iĜa[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ���� ��2�H(���H3k7HS�M5G�22G�?��Gp
͜��'f�/-,2�CR�>�D!�M#{Z/���3�����4y H "�c/u/�/�0B_����=jc��t�!�/ �/�"t32���~�/6  ��UP%�Q%��%�|T���S62�q?'e	'�� � �2I�� �  ��+==��ͳ?�;	��h	�0�I  �n @�2�.���Ov;��ٟ?&gN	 [OaA''�uD@!� Cb@C�@F#H!�/�O�O sb
�ATb@�@�@��@$�e`0Bb@QA�0Y�v: �13Uwz $oV_�/z_e_�_�_	���( �� -�2�1�1ta�UDa�c���:A-���~.  �?�ff���[o"o�_U�`oXâ�Q8���o�j>�1  Po�V(���eF0��f�Y���L�?˙���xb�P<
�6b<߈;����<�ê<�? <�&�,�/aA�;r�@Ov0P?offf?�0?&ipޘT@�.{r�J<?�`�u#	�B dqt�Yc�a�Mw �Bo��7�"�[�F� �j�������ُ� ���3����,���~(�E�� E��3?G+� F��a�� ҟ�����,��P�(;���B�pAZ�>� �B��6�<OίD���P� �t�=���a�s������6j�h��7o��>�S��O�����Fϑ�A�a�_���C3Ϙ�/�%?��?Ƀ��������#	���P �N||CH����Ŀ������@�I�_�'�3A��A�AR1A�O�^?�$�?���� �±
=�ç>����3�W
=�#� U���e���B��@���{����<����(�B��u��=B0�������	��b�H�F�G����G��H��U`E���C��+��I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻�������� � �9�$�]�H�Z��� ~�������������# 5 YD}h�� �����
C .gR����� ��	/�-//*/c/ N/�/r/�/�/�/�/�/ ?�/)??M?8?q?\? �?�?�?�?�?�?�?O �?7O"O[OmOXO�O|O �O�O�O�O�O�O�O3_:Q(������b���gUU��xW_i_2�3�8��_<�_2�4Mgs�_�_��RIB+�_�_�a?���{�mi�Go5okoYo�o}l��P'rP�nܡݯ�o=_`�o�_�[R?�Q�u���  �p���o��/�� S��z
uүܠ�������ڱ�����������  /�M�w��e��������l2 wF�$��Gb���t��a�`�p�S�C��y�@p�5�G�Y�۠F�� Dz��� F�P D��]����پ��ʯܯ�� ��~�?��ͫ@@�?�K��K���K���
 �|�������Ŀֿ �����0�B�T�f�ܽ�V� ���{���1��$PARA�M_MENU ?�3�� � DEF�PULSEr�	�WAITTMOU�T��RCV�� �SHELL_�WRK.$CUR�_STYL���	�OPT��PT�B4�.�C�R_DECSN���e��� �ߣ����������� !�3�\�W�i�{����USE_PROG %��%�����CCR���e�����_HOST !F��!��:���T�`�V��/�X����_TIME��^���  ��GDEB�UG\�˴�GINP_FLMSK�����Tfp����PGA�  ����)CH�����TYPE���������� � -?hcu �������/ /@/;/M/_/�/�/�/ �/�/�/�/�/??%?�7?`?��WORD �?	=	RS�fu	PNSU�Ԝ2JOK�DRT�Ey�]TRACE�CTL 1x3���� �`l m&�`�`�>�6_DT Qy3�%@��0D � [ `2@,6DU-6D.6D/6D06D16A�c2@�`8B V�8BR�8BM 8BJ�8BTF�8B6D6D	6DU
6D6D6D6DE6D6D^�8B6DU6D6D6D6D�8B6D6D~P8BA6DV�8Bj�8B6DA6DҀ8B�8B!6DE"6D#6D�8B%6DU&6D'6D(6D)6D*6D5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m�� ������Ǐن.A�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� r�����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ����������� �*��$PGT�RACELEN � )�  ���(��>�_�UP z��e�m�u�Y�n��>�_CFG {�m�W�(�n����PКӂ�DEFS_PD |���a�P��>�IN��T_RL }��(��8����PE_CO�NFI��~m�'�mњ��ղ�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�p�ح֚��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P;t _��������  Dz (�
 H�X~i�� ����/�/D/�//h/S/�/��
V�7.10beta�1��  A��E�"ӻ�Ay (�� ?!G��!/>���"����!����!BQ��!A\� �!���!2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?OO :O%O7OpO[O�OO�O �O�O�O�O_�O6_!_ Z_E_~_i_�_�_�_�_ �_�_'o2o�_VoAo So�owo�o�o�o�o�o �o.R=v1�<�/�#F@ �y�} ��{m��y=��1� '�O�a��?�?�?���� ��ߏʏ��'��K� 6�H���l�����ɟ�� �؟�#��G�2�k� V���z��������o ��ίC�.�g�R�d� ���������п	��� -�?�*�cώ���� �������B�;� f�x�������DϹ��� ���������7�"�[� F�X��|������� ����!�3��W�B�{� f��������� ��� ��/S>wbt ������ =OzόϾψ��� �ϼ� /.�'/R�d� v߈߁/0�/�/�/�/ �/�/�/#??G?2?k? V?h?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O���O�O�O_ _?_*_c_N_�_r_�_ �_�_�_�_o�_)oT fx�to���/ �o/>/P/b/t/ mo�|���� ���3��W�B�{� f�x�����Տ����� ��A�S�>�w�b��� �O��џ������+� �O�:�s�^������� ͯ���ܯ�@oRodo �o`��o�o�o��ƿ�o ���*<N�Y�� }�hϡό��ϰ����� ���
�C�.�g�Rߋ� v߈��߬�����	��� -��Q�c�N�ﲟ�� ��l��������;� &�_�J���n������� ����,�>�P�:L ����������� �(�:�3��0iT �x�����/ �///S/>/w/b/�/ �/�/�/�/�/�/?? =?(?a?s?��?�?X? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O*\&_8_r���_�_��$PL�ID_KNOW_�M  ��� Q�TSV ����P��?o"o4o�O�XoCoUo�o R�SM_GRP 1��Z�'0{`�@�`uf�e�`
�5� �g pk'Pe ]o�����������SMR�c�b�mT�EyQ}? yR ����������폯��� ӏ�G�!��-����� ������韫���ϟ� C���)���������`��寧���QST�a�1 1��)��v�P0� A 4� �E2�D�V�h������� ߿¿Կ���9��.� o�R�d�vψ��ϬϾϔ���2�0� Q�<3��3�/�A�S��4l�~ߐߢ��A5���������6
��.�@��7Y�k�}����8���������MAD  �)��PARNU/M  !�}o+���SCHE� S�
���f���S��UPD�f�x��_C�MP_�`H�� �'��UER_CHK-���ZE*�<RSr��_�Q_M�OG���_�X�__RES_G��!� ��D�>1bU �y�����/ �	/����+/ �k�H/g/l/��Ї/ �/�/�	��/�/�/� X�?$?)?���D?c?�h?����?�?�?�V� 1��U�ax�@c�]�@t@(@c�\�@�@D@c�[�*@��THR_INRr�J�b�U�d2FMASS?O �ZSGMN>OqCMO�N_QUEUE ���U�V P~P *X�N$ UhN�FV��@END�A��IEcXE�O�E��BE�@|�O�COPTIO�G���@PROGRAoM %�J%�@��?���BTASK_�IG�6^OCFG ���Oz��_�PDA�TA�c��[@Ц2=�DoVohozo�j 2o�o�o�o�o�o�);M jINFO
[��m��D�� ������1�C� U�g�y���������ӏ����	�dwpt�l �)�QE DIT ���_i��^WER�FLX	C�RGA�DJ �tZAЄ����?נʕFA��I�ORITY�GW�>��MPDSPNQ�����U�GD��OT�OE@1�X� _(!AF:@E� �c�Ч!tcp|n���!ud��>��!icm���?n<�XY_�Q�X�{��Q)� *�1�5��P��]�@� L���p��������ʿ ��+�=�$�a�Hυ�z��*��PORT)Q�H��P�E��_CARTREPP|X��SKSTA�H^�
SSAV�@�tZ�	2500H8�63���_x�
�'��*X�@�swPtS��ߕߧ���URGE��@B��x	WF��DO�F"[W\��������WRUP_DE?LAY �X��ԟR_HOTqX	B%��c���R_NOR�MALq^R��v�S�EMI�����9�Q�SKIP'��tUr�x 	7�1�1� �X�j�|�?�tU���� ����������$ J\n4���� ����4FX |j����� ��/0/B//R/x/�f/�/�/�/tU�$R�CVTM$��D��� DCR'����Ў!C`N�C��d�C��o?���>��L<|��{:��g�&���/���%��t����|���}'�:�o?�� �<
6b<߈�;܍�>u.��?!<�& �?h?�?�?�@>��?O  O2ODOVOhOzO�O�O �O�O�O�?�O�O__ @_+_=_v_Y_�_�_�? �_�_�_oo*o<oNo `oro�o�o�o�_�o�o �o�o�o8J-n ��_������ �"�4�F�X�j�U�� ����ď���ӏ�� �B�T��x������� ��ҟ�����,�>� )�b�M����������� �ïկ�Y�:�L�^� p���������ʿܿ�  ����6�!�Z�E�~� ��{ϴϗ�����-��  �2�D�V�h�zߌߞ� ����������
���.� �R�=�v��k��� �������*�<�N� `�r������������ ����&J\? �������� "4FXj|���!GN_ATC �1�	; �AT&FV0E0��ATDP/6/9/2/9��ATA�,�AT%G1%B�960�++U+�,�H/,�!�IO_TYPE � �%�#t�R�EFPOS1 1}�V+ x�u/�n�/j�/
=�/ �/�/Q?<?u??�?4?�?X?�?�?�+2 1�V+�/�?�?\O�?x�O�?�!3 1�O�*O<OvO�O�O_�OS4 1��O�O�O_��_t_�_+_S5 1�B_T_f_�_o	oBo>�_S6 1��_�_��_5o�o�o�oUoS7 1�lo~o�o�oH�3l�oS8 1� %_����SMASK 1��V/  
?�M��XNOS/�r�����~�!MOTE  n���$��_CFG ᢫��q���"PL_�RANG�����POWER ������SM_DRYPRG %o��%�P��TART� ��^�UME_PRO-�?����$�_EXEC_EN�B  ���GS�PD��Րݘ��T3DB��
�RM�
��MT_'�T�����OBOT_NA_ME o�����OB_ORD_�NUM ?��b!H863�  �կ����PC_TIMoEOUT�� x�oS232Ă1��� LTEA�CH PENDA1N��w��-���Mainte�nance Co#ns���s�"���?KCL/Cm��
�
���t�ҿ ?No Use-��8Ϝ�0�NPO�򁮋���.�C7H_L������q�	��s�MAVA#IL�����糅���SPACE1 2��, j�߂�D��s�߂� �{S�?8�?�k�v� k�Z߬��ߤ��ߚ�  �2�D���hߊ�|�� `����������  �2�D��h��|����`���������y���2����0�B���f� ����{���3);M_ ������/� /44FXj| */���/�/�/?(??=?5Q/c/u/�/ �/G?�/�/�?O�?$OEO,OZO6n?�?�? �?�?dO�?�?_,_�O A_b_I_w_7�O�O �O�O�O�_�O_(oIo@o^oofo�o8�_ �_�_�_�_�oo6oE�f){���Gw �o� �:��
M� ��� *�<�N�`�r������� w���o�収���d.��%�S�e�w��� ��������Ǐَ��� Θ8�+�=�k�}����� ��ůׯ͟����%� '�X�K�]��������� ӿ������#�E��W� `� @ �������x�����\�e����������� R�d߂�8�j߬߾߈� �ߤ����������0� r���X�������@������8����
�����_MODE � �{��S �"�{|�2�0��ψ��3�	S|)CWORK_AD���=9(+R  ��{�`� �� _?INTVAL���d����R_OPTI[ON� ��H �VAT_GRP �2��up#(N�k| ��_����� /0/B/��h�u/T�  }/�/�/�/�/�/�/? !?�/E?W?i?{?�?�? 5?�?�?�?�?�?O/O AOOeOwO�O�O�O�O UO�O�O__�O=_O_ a_s_5_�_�_�_�_�_ �_�_o'o9o�_Iooo �o�oUo�o�o�o�o�o �o5GYk-� ��u����� 1�C��g�y���M��� ��ӏ叧�	��-�?� Q�c������������ ���ǟ�;�M�_�����$SCAN_GTIM��_%}��R �(�#(�(�<04+d d 
!AD�ʣ��u�/X�����U��25�����dA�8�H�g��]	����������dd�x�  P~���� ��  8� ҿ�!���D��$�M�_�q� �ϕϧϹ��������8ƿv��F��X��/� ;�o�b��pm��t�_DiQ̡  � l�|�̡ ĥ�������!�3�E� W�i�{�������� ������/�A�S�e� ]�Ӈ����������� ��);M_q ������� r���j�Tfx� ������// ,/>/P/b/t/�/�/�/p�/�/�%�/  0�� 6��!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O *�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo �O�OJ�o�o�o�o�o �o�o 2DVh z�������
�7?  ;�>�P� b�t���������Ǐُ ����!�3�E�W�i��{�������ß � ş3�ܟ��&�8�J��\�n�������������ɯ����,�� �+�	12�345678��W 	� =5���@f�x���������� ���
��.�@�R�d� vψϚ�៾������� ��*�<�N�`�r߄� �Ϩߺ��������� &�8�J�\�n�ߒ�� �����������"�4� F�u�j�|��������� ������0_�T fx������ �I>Pbt �������! /(/:/L/^/p/�/�/ �/�/�/�/�2�/�?�#/9?K?]?�i�Cz  Bp˚ /  ��h2��*��$SCR_GR�P 1�(�U8�(�\x�d�@ � ��'�	 ?�3�1 �2�4(1*�&�I3�Fp1OOXO}m��CD�@�0ʛ)���H�UK�LM-10�iA 890?�9�0;��F;�M61�C D�:�CP��1

\&V�1	�6F� �CW�9)A7Y	(R�_��_�_�_�_�\���0i^�oOUO>o Po#G�/���o'o�o��o�o�oB�0ƐrtAA�0* C @�Bu&Xw?���ju�bH0{UzAF?@ F�`�r� �o�����+�� O�:�s��mBqrr����������B�͏b�� ��7�"�[�F�X���|� ����ٟğ���N��� AO�0�B�CU
L���xE�jqBq>HE����$G@�@pϯ BȆ��G�I
E�0E�L_DEFAUL�T  �T���E��MI�POWERFL � 
E*��7�WF�DO� *��1E�RVENT 1����`(�� L�!DUM_EI�P��>��j!AF_INE�¿C�O!FT�����r�!o:� ���a�!RPC_M'AINb�DȺPϭ�Nt�VIS}�Cɻ�����!TP��PU��ϫ�d��E�!
P�MON_PROX	YF߮�e4ߑ��_��f����!RD�M_SRV�߫�g��)�!R�IﰴYh�u�!
v�M���id���!RL�SYNC��>�8|���!ROS��4��4��Y�(�}��� J�\����������� ��7��["4F� j|����!��Eio�ICE_�KL ?%� �(%SVCPRG1n>���3��3���4//�5./3/�6V/[/��7~/�/��D�/�9�/�+�@��/�� #?��K?��s?�  /�?�H/�?�p/�? ��/O��/;O��/ cO�?�O�9?�O� a?�O��?_��?+_ ��?S_�O{_�)O �_�QO�_�yO�_� �Os����>o�o }1�o�o�o�o�o�o�o ;M8q\� �������� 7�"�[�F��j����� ��ُď���!��E� 0�W�{�f�����ß�� �ҟ���A�,�e� P���t��������ί��y_DEV ���MC:��@`!�OU�T��2��RE�C 1�`e�j�{ �� 	 � ����˿���ڿ��
 �`e���6�N� <�r�`ϖτϦ��Ϯ� ������&��J�8�n� ��bߤߒ��߶����� ��"��2�X�F�|�j� ������������� �.�T�B�x�Z�l��� ����������, P>`bt��� ���(L: \�d�����  /�$/6//Z/H/~/ l/�/�/�/�/.��/? �/2? ?V?D?f?�?n? �?�?�?�?�?
O�?.O @O"OdORO�OvO�O�O �O�O�O�O__<_*_ `_N_�_�_x_�_�_�_ �_�_oo8oo,ono \o�o�o�o�o�o�o�o �o "4jX� �������� �B�$�f�T�v����� �������؏��>��,�b�P�r���p�V [1�}� P
�l!������ �<��TYPE\���HELL_CFG� �.��� ���r�����RSR������ӯ����� ��?�*�<�u�`��������������/  �%�3�PE��Q�\�ӐM�Lo�p��d��2Ӑ�d]�K�:�HK 1�H� u����� ��A�<�N�`߉߄� �ߨ������������&�8��=�OMM ��H���9�FTOV_ENB&�1��OW_REG_U�I���IMWAI�T��a���OUTr������TIM��w���VAL��>��_UNIT��K��1�MON_ALI�AS ?ew� ( he�#������ ����Ӕ��);M ��q����d� �%�I[m �<����� �!/3/E/W//{/�/ �/�/�/n/�/�/?? /?�/S?e?w?�?�?F? �?�?�?�?�?O+O=O OOaOO�O�O�O�O�O xO�O__'_9_�O]_ o_�_�_>_�_�_�_�_ �_�_#o5oGoYokoo �o�o�o�o�o�o�o 1C�ogy�� H����	��-� ?�Q�c�u� ������� ϏᏌ���)�;�� L�q�������R�˟ݟ �����7�I�[�m� �*�����ǯٯ믖� �!�3�E��i�{��� ����\�տ����� ȿA�S�e�wω�4ϭ� �����ώ����+�=� O���s߅ߗߩ߻�f� ������'���K�]� o���>�������� ���#�5�G�Y��}����������o��$S�MON_DEFP�RO ������ �*SYSTEM�*  d=��R�ECALL ?}��� ( �}/�xcopy fr�:\*.* vi�rt:\tmpb�ack7=>in�spiron:12732 Ybt\�� }0.a6�HZ_��4�/s:orderfil.dat��Mbt�� }+/mdb:�MZ ��/�-�Qb/ t/�/�/�</�a/�/�??�!
xyzrate 61 �/@�/�/n?�?�?�%.7>M(4804 H?Z?�?�?O�(3.@�= aOsO�O�O� *�IO@�4YO�O�O_�)../ A?�8�On_�_�_%.�/ G_�1^_�_oo&O8O �O�Omoo�o�O�O�O Zo�o�o"_4_�_X_ i{��_�_C�_� ��o0oBoToe�w� ���o�oI��o���� �,�Pa�s����� �;��`����(? ��̟ޟo������?M*28�?Y�����!� 3�����a�s������� E���Y�����!�3� F�£ݿnπϒϥ�6� H�Š^�����&�8� ��ܿm�ߑߤ���ȿ Z������"�4���X� i�{��ϲ�C����� ����0�����e�w�0�������106�?X� ���� �2��������n�����92076GY��!�3� �߽as����E �Y��/!�3�F� ��n/�/�/��6/H/ � ^/�/??&8� �m??�?���Z?��?�?O!7�$SN�PX_ASG 1߸���9A�� P 0 �'%R[1�]@1.1O 9?�$3%dO�OsO�O�O �O�O�O�O __D_'_ 9_z_]_�_�_�_�_�_ �_
o�_o@o#odoGo Yo�o}o�o�o�o�o�o �o*4`C�g y������� 	�J�-�T���c����� ��ڏ�����4�� )�j�M�t�����ğ�� ����ݟ�0��T�7� I���m��������ǯ ٯ���$�P�3�t�W� i��������ÿ�� ��:��D�p�Sϔ�w� ���ϭ��� ���$�� �Z�=�dߐ�sߴߗ� �������� ��D�'� 9�z�]������� ��
����@�#�d�G� Y���}����������� ��*4`C�g y������ 	J-T�c�� ����/�4// )/j/M/t/�/�/�/�/��/�/�/?0?4,DPARAM �9E�CA �	���:P�4�0$HO�FT_KB_CF�G  q3?E�4P�IN_SIM  9K�6�?�?�?�0�,@RVQSTP_DSB�>�21On8�J0SR ��;�� & MULT�IROBOTTA�SK=Oq3�6T�OP_ON_ER�R  �F�8�AP_TN �5�@�A�BRIN�G_PRM�O �J0VDT_GRP� 1�Y9�@  	�7n8_(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2Dkhz�� �����
�1�.� @�R�d�v��������� Џ�����*�<�N� `�r���������̟ޟ ���&�8�J�\��� ��������ȯگ��� �"�I�F�X�j�|��� ����Ŀֿ���� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�tߛߘߪ߼��� ������(�:�a�^� p�����������  �'�$�6�H�Z�l�~���������������3V�PRG_COUN�T�6��A�5ENB�OM=�4J_UPD 1��;8  
q2� ����� )$ 6Hql~��� ��/�/ /I/D/ V/h/�/�/�/�/�/�/ �/�/!??.?@?i?d? v?�?�?�?�?�?�?�? OOAO<ONO`O�O�O �O�O�O�O�O�O__ &_8_a_\_n_�_�_�_�YSDEBUG�" � �Pdk	�PS�P_PASS"�B?�[LOG ���m�P��X�_  �g�Q
MC:\d�_b_MPCm��o�o��Qa�o �vfS_AV �m:dlUb�U\gSV�\�TEM_TIMEw 1�� (�`��Q�a�2o	T1S�VGUNS} #'�k�spASK_?OPTION" ��gospBCCF�G ��| 8�b�{�}`��� �a&��#�\�G���k� ����ȏ������"� �F�1�j�U���y��� ğ���ӟ���0��T�f��UR���S��� ƯA������ ��D� �nd��t9�l������� ��ڿȿ�����"� X�F�|�jϠώ��ϲ� ��������B�0�f� T�v�xߊ��ߦؑ��� ����(��L�:�\� ��p���������� � �6�$�F�H�Z��� ~������������� 2 VDzh�� �������4 Fdv���� ��//*/�N/</ r/`/�/�/�/�/�/�/ �/??8?&?\?J?l? �?�?�?�?�?�?�?�? OO"OXOFO|O2�O �O�O�O�OfO_�O_ B_0_f_x_�_X_�_�_ �_�_�_�_oooPo >otobo�o�o�o�o�o �o�o:(^L np�����O� �$�6�H��l�Z�|� ����Ə؏ꏸ���� 2� �V�D�f�h�z��� ��ԟ����
�,� R�@�v�d��������� ίЯ���<��T� f�������&�̿��ܿ ��&�8�J��n�\� �π϶Ϥ�������� ��4�"�X�F�|�jߌ� �ߠ����������� .�0�B�x�f��R��� ���������,��<� b�P�������x����� ����&(:p ^�������  6$ZH~l ��������/ &/D/V/h/��/z/�/��/�/�/�&0�$T�BCSG_GRP� 2��%��  �1 
? ?�  /?A? +?e?O?�?s?�?�?�?��?�;23�<d�, �$A?1	� HC���6>�@E�5CL  �B�'2^OjH4Jݸ�B\)LFY g A�jO�MB��?F�IBl�O�O�@�JG|_�@�  D	�15_ __$YC-P{_F_$`_j\��_�]@0�> �X�Uo�_�_6oSoo�0o~o�o�k�h�0	V3.00'2�	m61c�c	�*�`�d2�o�e>əJC0(�a�i �,p�m-  �0�����omvu1JC�FG ��%� 1 #0vz��rrBrv�x�� ��z� �%��I�4� m�X���|�������� ֏���3��W�B�g� ��x�����՟����� ���S�>�w�b��� ��'2A ��ʯܯ��� ���E�0�i�T���x� ��ÿտ翢����/� �?�e�1�/���/�� �Ϯ��������,�� P�>�`߆�tߪߘ��� ���������L�:� p�^��������� ��� �6�H�>/`�r� ���������������  0Vhz8� �����
. �R@vd��� ����//</*/ L/r/`/�/�/�/�/�/ �/�/�/?8?&?\?J? �?n?�?�?�?�?���? OO�?FO4OVOXOjO �O�O�O�O�O�O__ �OB_0_f_T_v_�_�_ �_z_�_�_�_oo>o ,oboPoroto�o�o�o �o�o�o(8^ L�p����� ��$��H�6�l�~� (O����f�d��؏� ��2� �B�D�V����� ��n����ԟ
���.� @�R�d����v����� ���Я���*��N� <�^�`�r�����̿�� �޿��$�J�8�n� \ϒπ϶Ϥ������� ߊ�(�:�L���|�j� �߲ߠ���������� 0�B�T��x�f��� �����������,�� P�>�t�b��������� ������:(J L^������  �6$ZH~ l��^���dߚ  //D/2/h/V/x/�/ �/�/�/�/�/�/?
? @?.?d?v?�?�?T?�? �?�?�?�?OO<O*O `ONO�OrO�O�O�O�O �O_�O&__6_8_J_ �_n_�_�_�_�_�_�_ �_"ooFo��po�o ,oZo�o�o�o�o�o 0Tfx�H� ������,�>� �b�P���t������� ��Ώ��(��L�:� p�^�������ʟ��� ܟ� �"�$�6�l�Z� ��~�����دꯔo� �&�ЯV�D�z�h��� ����Կ¿��
��.π�R�@�v�dϚτ� s ���� ��������$TBJO�P_GRP 2����� O ?������������x/JBЌ��9�� �< �zX���� @����	 �C�� >t�b  C����>��͘Րդ��>̚йѳ33=��CLj�ff�f?��?�ffB@G��ь�����t�ц��>�(�\)��ߖ�E噙�;���hCYj��  �@h��B�  A�����f��C� � Dhъ�1���O�4�N����
�:���Bl^���j�i�l�l����A�ϙ�A�"��D��֊=qH������p�h�Q�;��A�j�ٙ7�@L��D	2��������$�6�>B�\p��T���Q�tsx�@33@���C����y�1����>G��Dh�������<���<{�h�@i� ��t� �	���K&� j�n|���p��/�/:/k/�ԇ����!��	V3�.00J�m61cI�*� IԿ��/��' Eo��E��E���E�F���F!�F8���FT�Fqe\�F�NaF����F�^lF����F�:
F�)�F��3G��G��G���G,I�!CH`��C�dTDU��?D��D���DE(!/E\��E��E�h��E�ME���sF`F+'�\FD��F`�=F}'�F���F�[
F����F��M;��;WQ�T,8�4` *Q�ϴ?�2���3�\�X/O��ESTP?ARS  ��	����HR@ABLE� 1����0��D
H�7 8��9
G
H�
H����
G	
H
�
H
HYE��
H�
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_Ht_�^:BS _� �J GoYoko}o�o�o�o�o �o�o�o1CU gy����`#oRL �y�_�_�_�_�O�O�O��O�OX:B�rNUM�  ����P��� V@P:B_?CFG ˭�Z��h�@��IMEBF_TT%AU��2@�GVERS�q���R 1���
 (I�/����b� �� ��J�\���j�|���ǟ ��ȟ֟�����0� B�T���x�������2��_���@�
��M�I_CHAN�� �� ��DBGLV����������ET�HERAD ?*��O�������xh�����ROUT�!��!������?SNMASKD��>U�255.���#������OOLOF/S_DI%@�u.��ORQCTRL �����}ϛ3rϧ� ����������%�7� I�[�:���h�z߯�A�PE_DETAI�"�G�PON_SV�OFF=���P_M�ON �֍�2���STRTCHK� �^�����VTCOMPAT���O�����FPROG� %^�%MU�LTIROBOT�Tݱ���9�PLA�Y&H��_INST+_Mް �������US�q��LCK����QUICKM�E�=���SCRE�Z�G�tps� ���u�z�����_��@@n�.�SR_�GRP 1�^�/ �O���� 
��+O=sa�쀚�
m���� ��L/C1g U�y����� 	/�-//Q/?/a/�/�	123456�7�0�/�/@Xt�1����
 �}i�pnl/� gen.htm�? ?2?�D?V?`Pan�el setupZ<}P�?�?�?�?�?�? �??,O>OPO bOtO�O�?�O!O�O�O �O__(_�O�O^_p_ �_�_�_�_/_]_S_ o o$o6oHoZo�_~o�_ �o�o�o�o�o�oso�o 2DVhz�1 '���
��.�� R��v���������Џ|G���UALRM��oG ?9� � 1�#�5�f�Y���}��� ����џן���,���P��SEV  �����ECFG ��롽�}A��   BȽ�
 Q���^���� 	��-�?�Q�c�u���Й��������� P�����I��?����(%D�6� �$�]� Hρ�lϥϐ��ϴ��π����#��G���� ��߿U�I_Y�H�IST 1�� � (�� ���3/SOFTP�ART/GENL�INK?curr�ent=edit�page,��,1����!�3��� �����menu��962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V