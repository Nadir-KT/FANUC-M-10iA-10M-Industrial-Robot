��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY T� u3|4|H �RG_STR1� � $TIT�P$I��1��{�����5��6�7�8�9�0��z���T��1�1�1 '�1
'2"GSBN�_CFG1  �8 $CNV_�JNT_* |$�DATA_CMN�T�!$FLAG�S�*CHECK��!�AT_CEL�LSETUP � P $HO_ME_IO,G�}%�#MACRO�"�REPR�(-DR�UN� D|3S�M5H UTOBA�CKU0 � ?$ENAB��!oEVIC�TI� � D� DX�!2ST� ?0B�#$�INTERVAL�!2DISP_UNsIT!20_DOn6�ERR�9FR_F�!2IN,GRE5S�!0Q_;3!4C_WA�471�8G�W+0�$Y $D�B� 6COMW�!2MO� H.	� \rVE�1$qF�RA{$O��UDcB]CTMP1_5FtE2}G1_�3�BԎ2FXD�#
� d $CARD_EXIST4�$FSSB_T�YP!AHKBD�_SNB�1AGN G�n $SLO�T_NUM�AP�REV4DEBU�� g1G ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�U0LEToE_OK�BUS�oP_CR�A$;4xAV� 0LACIw�1�R�@k �1$@M{EN�@$D�V��Q`PvVA{�B�L� OU&R ,�A�0�!� B� L�M_O�
eR�"C�AM_;1 x�r$ATTR84�@� ANNN@5�IMG_HEIG�H�AXcWIDTH�4VT� �UU0F�_ASPEC�A;$M�0EXP�.@�AX�f�CF�D X $GR� �� S�!.@B�PNF�LI�`�d� UIR�E 3T!GITCH�+C�`N� S�d_LdZ`AC�"�`EDp*�dL� J�4S�0� �<za�!p;G0� � 
$WARNM�0f�!�@� -s�pNST� CORyN�"a1FLTR{u�TRAT� T}p  $ACCa1�p��|{�rORIضP�C�kRT0_S�~B\qHG,I1� [ T�`�"3I��pTYD�@*2 �3`#@� �!�B*HEDDcJ* Cd�2_�U3_�4_�5_�6_��7_�8_�94c'��CO�$ <�� �o�o�hK3 1#`O�_Mc@AC t e� E#6NGPvABA� �c1�Q8��`,��@nr1�� �d�P�0e�]p� cvnpUP&Pb26��4�p�"J�p_R�rPB�C��J�rĘߜJV �@U� B��s}�g1�"vYtP_*0OFS&Rw @� RO_K8�T��aIT�3T�NOM_�0�1p�3W >��D �� Ќ@�2�hPV��mEX�p� Ĝ0g0ۤ�p�r
$�TF�2C$MD3&i�TO�3�0U� F�/ ��Hw2tC%1(�Ez�g0#E{`"F�"F�40CP@��a2 �@$�PPqU�3N)ύLRևAX�!DU�v�AI�3BUF�F8=�@1 |pp��ցpPIT� PP��M�M�y��F>�SIMQSI�"�ܢVAڤT�F@�w T�`(zM��P�B^�qFACTb�@EW�P1�BTv?��MC� �$�*1JB`p�*1DEC��F�������� �H0CHN�S_EMP1�$G��8��@_4�3�p2|@P��3�TCc�(r /�0-sx��ܐ� MB0i��!����JR� i�_SEGFR��Iv *�aR�TpN�C���PVF4>�bx &��f{uJc!� Ja��� !28�ץ�AJ���SIZ�3S�c�B��TM���g��JaRSINFȑb���q�� ��н����L�3��B���CRC�e�3CCp����c��mc� �b�1J�cѿ�.����D$ICb�Cq�5r��`���@v�'���EV����zF��_��F,pN��ܫ�?�4�0A�! �r���h�� ���p�2�͕a�� ��د\qR�Dx Ϗ��o"27��!ARV�O`C�$L	G�pV�B�1�P��@��t�aA�0'�|�+0Ro�� MEp`"1 �CRA 3 AZ�V�g6p�O �FCCb�`�`F�`K������ADI��a�A �bA'�.p��p�`�c¢`S4PƑ�a�AMP$��-`Y�3P�M�]p�UR��QUA1  $.@TITO1/S@S��!����"0�DBP�XWO��B0!5�g$SK���FDBq��!"�"�PR��� 
� =����!# �S q1$2�$z���L�)$�/���R� %�/�$C�!&?��$ENE�q.'�*?�Ú RE�p2(�H ��O�07#$L|3$$�#�B�[�;���FO_D��ROSr�#�������3RIGGE�R�6PApS����E�TURN�2�cMR-_8�TUw��0�EWM��M�GN�P���BLAH�<E��y�P��&$P�" �'P@�Q3�CkD{��DQ���4�11��FGO_AWAY�B�MO�ѱQ#!��DCS_�)  �PIS� I gb @{s�C��A��[ �B�$�S��AbP�@�EW�-�TNTVճ�BV �Q[C�(c`�UWr�P��J��P�$0��SAF�E���V_SV�bEOXCLU��n'ONL2��SY�*a�&�OT�a'�HI_�V�'���B���_G *P0� 9�_z���p �!�@SG�� +nrr�@�6Acc*b��G�#@E�V�.iHb?fANNUNX$0.$fdID�U�2�SC@�`�i�a��jP�f��z��@I$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6�a�QM�SW�E. 8Q�KgEYI5���TM�100s�qA�vIN��#��b��/ D��H7OST_P!�rT���ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  A8	=ȳ�ј Tk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&Q�DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F�码df�J� �q��T�E�T+6 H�bLL_DUs�~a3@{�0�3:���OTX"����s	q��0NO�AUTO�!7�p!$)�$�*��c4�(��C� 8�C, �"�q&�L�� 8H *8�LH <6� ���c"�`, `Ĭ�k� ��q��q��sq��~q���7��8��9��0T����1��1̺1ٺU1�1�1 �1ʕ1�2(�2����2�̺2ٺ2�2�2� �2�2�3(�3R��3��̺3ٺ3�U3�3 �3�3��4(�a��?��!9 A<�9�&�z��I��01���M�O�FE@'@΂ : ,6��Q?3 �@P?9��
5�9�E�@A�q�A�� ;p$TP~�$VARI:��ፂ@P2�P< ���TDe���K`�Q���"���BAC��"= T�p��e$)�_,�bn�kp+ IFI@G�kp�H  ��P��Y�@`�!>t� ;E��sC�ST�D� D���c�<� 	C��{��_����l���R  ���F?ORCEUP?b���FLUS�`H�N�>�F ���RD_CM�@E������ ��@v\MP��REMr F�Q���1k@���7Q
Kr4	NJ�5EFFۓ�:�@IN2Q��OV�O�OVA�	TR3OV���DTՀ�DTMX� ��@ �
ے_PH"p��CL��_TpE�@�p2K	_(�Y_T��v*(��@A;QD� ������!0tܑ0RQ���_�a����M�7�CL�dρR�IV'�{��EAR6ۑIOHPC�@��2��B�B��CM9@����R �GCLF�e!DYk(M�ap#5TuDG��� ��%��FSSD �s?C P�a�!�1���PQ_�!�(�!1��E�3�!3�+5�&�GR)A��7�@��;�P�W��ONn��EBUG_SD2H`{�_E A �p|뀢0�TERM`5yBi5��ORI#�e0Ci5�p�SM_��P��e0D�7 �T�A�9Ei5 ��UP\�F� -��A{�AdPw3S@B�$SEG�:� EL�{UUSE�@NFIJ�B$�;1젎4�4�C$UFlP=�!$,�|QR@��_G�90Tk�D�~SNST��PAT����AP'THJ��E�p% B`�'EC���A�R$P�I�aSHFT�y�A�A�H_SHOQRР꣦6 �0$�7rPE��E�OVR=���aPI�@�U�b �QAYLOW����IE"�r�A��?���ERV��XQ�Y��mG�>@�BN��U\��Rz2!P.uASYMH��.uAWJ0G�ѡE q�A�Y�R�Ud>@ ��EC���EP;�uP�;�6WOR>@M`�]0SMT6�G3�cGR��13�aPAL@���`�q�uH � u���TOCA��`P	P�`$OP@����p�ѡ�`0YO��RE�`R4Cb�AO�p낎Be�`�R�Eu�h�A��e$7PWR�IMu�R�R_�cN��q=B �I&2H���p_AD�DR��H_LENAG�B�q�q�q$�R��S�JڢSS��SKN��u\��u̳�uٳ�SE�A�jrS��M-N�!K�����b����OLX��px����`ACRO3p J�@��X�+��Q��N6�OUP3�b_�IX��a�a1��}� ����(��H��D��`ٰ��氋�IO2ES�D�����N
�7�L $l��`Y!�_OFFr�PR�M_���aTT�P_+�H:�M (�|pOBJ]"�p��-$��LE~Cd����N � ��֑AKB_�TqᶔS�`lH�LVh�KR"~uHITCOU��[BG�LO�q����h�����`��`S9S� ���HW�#A�:�Oڠ<`INC�PU2VISIO W�͑��n��to��to�~ٲ �IOLN��P 8��R��p�$SLob PU�T_n�$p��P�& ¢��Y F_AS:�"Q��$L�������Q  U�0	P4A0��^���ZPHY��-�2�y��UOI �#R `�K����$�u�"pPpk�`��$�������UJ5��S-���NE6WJO9GKG̲DIS����1Kp���#T (�uAqVF�+`�CTR�C�
�FLAG2��LG�dU ���؜�~13LG_SIZ�����b�4�a��a�FDl�I`�w� m�_�{0 a�^��cg���4������Ǝ���{0��� SC#H_���a7�N�d�VW���E�"����D4��UM�Aљ`LJ�n@�DAUf�EAU�0p��d|�r�GH�ba����BOO��WL3 ?�6 IT���y0�REC��SCR ܓ�D
�\���MARGm�!��զ  ��d%�����S�����W���U� �JGM�[�MNCHJ���F�NKEY\�K��PRG��UF��7P��FWD��HL��STP��V��=@�����RS��HO`����C9T��b ��7�[�UL���6�(RD� ��2��Gt��@PO���������MD�FOCUޛ�RGEX��TU%I��I��4�@� L�����P�����`��P��NE��CA�NA��Bj�VAI�LI�CL !�UDCS_HII4��s�O�(!�S����S��D���BUFUF�!X�?PTH$m���v`�ě�*��AtrY�?P���j�3��`OS1Z2�Z3Z��� Z � ��[aEȤ��.ȤIDX�dPSRraO���zA�STL��R}�Y&�� Y$E�C���K��&&9�п![ LQ��+00�	P���`�#qdt
�U�dw<���_ \ �`4Г��\��Ѩ#\0C4�] =��CLDPL��UTRQLI��dڰ�)�$FLG&�� 1��#�D���'B�LD8�%�$�%ORGڰ5� 2�PVŇVY8�s�T�r�$}d^ ���$6��$�%S�`T� �B0��4�6RCLMC��4]?o?�9�9MI��p}d_ d=њR�Q(��DSTB��p� ;F�HHA�X�R JHdLEXWCESrEM!p
�a`�/B�Ta�B���`a�p=F_A@7Ji��KbOtH� K�d�b \Q���v$M�BC�LI|�)SREQUIR�R�a.\o��AXDEBUZ�AL
t M��c�b�{P��4��2ANDRѧ``d;�2�ȺSDC��N�INl�K�x`찄�X� N&��aZ���UPST� enzrLOC�RIrp�EX<fA�p�9A� ��`AQ��f� XY�OND�rMF,Łf�s"��}%��e/� �a�FX3@I�GG�� g ���t"��ܓs#N�s$R�a%��iL��hL�xv�@�DATA#?pE�%�E���Y��Nh t $+MD`qI}�)nv� ytq�ytHP`�Pxu��<(�zsANSW)�yt�@��yuD+�)AO����0o�i �@C�Uw�V�p 09AAR;R2��j Du�{Q���7Bd$CALI�A@��G��2��R�IN��"�<9INTE��Ck�r^�آX�]���_N�qlk����9�D���Bm��D3IV(�E�DH�@��:�qnI$V,��Sv�$��$Z��X�o�*����o�H �$BEL�T�u!ACCEL��.�~�=�IRC��� ���D�T�8��$PS�@�"L   Šp��#^�S�Eы T�PATH3���I���3x�p�A_W��ڐ����2nC��4�_M=G�$DD��T���$FW�Rp9���I�4��DE7�P�PABN��ROTSPEE�[g�� �J��[�C@4�x��$USE_+�VP�i��SYY���1 �qYN!@A�ǦOsFF�qǡMOU��3NG���OL����INC�tMa6��HBx��0HBENCS+��8q9Bp�4�FDm�IN��Ix�]��B��V�E��#�y�23_UyP񕋳LOWL�A��p� B���Du�@9B#P`�x ���BCv��r�MOSI��BM�OU��@�7PERC7H  ȳOV��â 
ǝ����D�Sc@F�@MP����� Vݡ�@y�j�LUk��GjĆp�UP=ó���ĶT�RK��AYLOA�Qe��A��x�����8N`�F�RTI�A$��MOUІ�HB�BS0�p7D5���ë�Z��DUM2ԓS_�BCKLSH_C x�k����ϣ����=���ޡ �	ACLA�L"q��1м@��C�HK� �S�RT�Y��^�%E1Qq_��޴_UM�@�C�#��SCL0�r�LMT_J1_L��"9@H�qU�EO�p��b�_�e�k�e�SPC`��u���N�PC�BN�Hz \P��C�0�~"XT��CN_b:�N9��I�SF!�?�V���U�/���x�dT���CB!�SH� :��E�E1T�T����0y���T��PA ��_P��_� =��Ơ���!����J6 L��@��OG�G�ToORQU��ONֹ���E�R��H�E�g_	W2���_郅T���I�I�I��	Ff`xJ�1�~1��VC3�0BD:B�1��@SBJRK�F9�0DBL_�SM��2M�P_D9L2GRV��0��fH_��d���COS���LNH���������!*,�aZ���fMY�_(��TH��)THET=0��NK23���"l��CB�&CB�CAA�B�"��!��!Ư&SB� 2�%GT	S�Ar�CIMa������,4#97#$DU���H\1� �:Bk6�2�:AQ(rSf$NE�D�`I��B+5��	$̀�!A�%�5�7���LPH�E�2���2SC%C%�2�-&FC0JM&̀V�8V��8߀LVJV!KV�/KV=KVKKVYKVgIH�8FRM��#X�!KH/KH=KHKKH�YKHgIO�<O�8OT�YNOJO!KO/KUO=KOKKOYKOM&�F�2�!+i%0d�7S�PBALANCE�_o![cLE0H_�%SPc� &�b&�b>&PFULC�h�b��g�b%p�1k%�U�TO_��T1T2�i/�2N��"�{� t#�Ѱ`�0�*�.��T��OÀ<�v IN�SEG"�ͱREV84vͰl�DIF�ŕ��1lzw��1mn`OaBpq�я?�MI{����nLCHWAR�Y�_�AB��!�$MECH�!o ��q�AX��P����7Ђ�`n 
�d(�nU�ROB��CRx��H���B'�MS�K_f`�p P �`_��R/�k�z�����1S�~�|�z�{�ؔ�z��qINUq�MTCOM_C� >�q  ���p~O�$NOREn�����pЂr 8fp GRe�uSD�0�AB�$XYZ�_DA�1a���DE�BUUq������s �z`$��COD��� L���p��$BUFINDX�|�  <�MOR^m�t $فUA� �֐���y��r�G��u � $SIMUL  S�*�xY�̑a�OBJE�`>̖ADJUS�ݐOAY_IS�D��3����_FI�=��Tu 7�~�6�'���p} =�C�}p�@b�DN��FRIr��T��RO@ \�E}�����OPWOYq�v}0Y�SYSBU/@v�$SOPġd����ϪUΫ}pPRUN,����PA��D���r\ɡL�_OUo��q�$)�IMA�G��w��0P_qIM��L�INv�K�?RGOVRDt�梄X�(�P*�J�|��0L�_�`]��0�RB�1�0��M��E�D}��p ��N�PMdֲ��1c�w�SL�`�q�w x $OwVSL4vSDI��DEX����#�$��-�V} *�N4�\@#�B�2�G�B�_�M��x� �q�E� �x Hw��p��AT+USW���C�0o��s���BTM�ǌ�I
�k�4��x�԰q�y Dw�E&���@E�r��7��жЗ�EXE��ἱ���8��f q�z @w���3UP'��$�pQ�XN����������� �PG΅{ h? $SUB�����0_���!�MPW�AIv�P7ã�LO�R���F\p˕$R�CVFAIL_C���BWD΁�v��DEFSP!p | Lw���Я�\���UNI+�����bH�R�+�}_L\pIP��t�P��p�}H��> �*�j�(�s`~�NN�`KETB�%�J�PE Ѓ~��J0SIZE\���X�'����S�OR��FORMAT�`��c ��WrEM�t��%�UqX��G��PLI��~p�  $ˀP_SWI�pq�J�_PL��AL_ S�����A��B���� C��D�$E���.�C_�U��� � � ���*�J3K0�����TIA4��5��6��MOM������h���ˀB��AD����������PU� NAR������H���m��� A$PI�6q��	��� ��K4�)6�U��w|`��SPEEDgPG��������Ի� 4T�� � @��SAMr`��\�]��MOV_�_$�@npt5��5���1���2��������'�2S�Hp�IN�'� @�+����4($<4+T+GAMMWf�1>'�$GET`�p����Da���

pLI�BR>�II2�$H�I=�_g�t��2�&E�;��(A�.� �&LW �-6<�)56�&]��v��p��V��$�PDCK���q��_?�����q�&����7��4���9+� ��$IM_SR��pD�s�rF��r�rL	E���Om0H]��0�	-�pq��P~JqUR_SCRN��FA���S_SAV�E_D��dE@�NOa�CAA�b�d@�$q� Z�Iǡs	�I� �J�K � ����H�L��> �"hq������ɢ �ɡ bW^US�A�
,M4���a��)q `��3�WW�I@v�_�=����MUAo�� � �$PY+�$W�P�vNG�{��P�:��RA��RH��RO�PL�����q� ��s'�%X;�OI�&�Zxe ���m�� p��ˀ�3s�O�O�O�O�O�a:a�_т� |��q� d@��.v��.v��d@���[wFv��E���% (��t;B�w�|�t�P���PMA�QU.a ��Q8��1��QTH�HOL�G�QHYS��ES���qUE�pZB��O.τ�  ـPܐ(��A����v�!�t�O`�q��u�"���FA�ÎIROG�����Q2����o�"��p��INFOҁ�׃V�����R�H�OI��� =(�0SLEQ������Y���O���Á���P0Ow0����!E0NU��A�UT�A�COPY��=�/�'��@Mg�N@��=�}1������ ���RG��Á���X_�P�$;ख�`��W��P��@��������EXT_CYC� btН�RpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�H�SdB����2�$��F�p���GPLeAdA
�TAR��Б@���P����裔d� ,�0F1L`�o@YN��K��M��Ck��PWR�+�9ᘐ��DELiA}�dY�pAD�a��QSKIPN4� �A�$�OB`�NT�FP��P_ $�M�ƷF@\bIpݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q�����q������ ���`���RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�d��REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"����+ ��2�Қ�߼ߠ��������3�қ�'�9�K�]�o���4�Ҝ�����������
�5�ҝ!�3�E�W�(i�{��6�Ҟ��������������7�ҟ�-?Qcu�8�Ҡ������^�SMSKÁ�lЩ�a��EkA�QR�EMOTE6������@�݂�q�IIO}5�IS�tR�9W@��� �pJ�"�������E�"�$DSB_SIG!N�1UQ�x�C\��p~ ��RS232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+��q��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�PHE#�0�����p_XP�C)�$FREEFROMS	pna��GET�0��UPD��A�2E#P� :���� !$U�SAN�na&����EcRI�0�RpRYq5*"_j@�Pm1�!�6'WRK9KD���6���QFRIEND��Q�RUFg�҃�0T�OOL�6MY�t�$LENGTH_;VT\�FIR�pC�@ˀE> +IUFI�N-RM��RGI<�1ÐAITI�$G�Xñ3IvFG2v7G�1���p3�B�GPR�p�1F�O_n 0��!RE��p�53҅U��TC��3A�A�F �QG(��":���e1 n!��J�8�%���%]�� �%�� 74��X O0�L��T�3H&��8���%b453%GE�W�0�WsR�TD����T��M����Q��T]�$V 2!����1�а91�8�0U2�;2k3�;3�: ifa�9-i�aQ��NSL��ZR$V��2BVwE�V�	V�B;���� �&�S�`��F�"�k�@��2a�PS�E ��$r1C��_$Aܠ6wPR��7vMU�c�S�t '�/89�� 0G�aV`��p�d`A���50�@��-�
25�S�� ��aRHW����B�&�N�SAX�!�A:@LA�h��rTHIC�1pI���X�d1TFEj�|�q�uIF_CH�3��qI܇7�Q�pG1@RxV���]��:�u�7_JF~�PRԀƱ��RVAT���� ��`���0RҦ�D9OfE��COUԱ���AXI���OFF{SE׆TRIGNS ���c����h������H�Y��IGMA�0PA�pJ�E�OR?G_UNEV�J���S�����d� �$CА�J�GgROU����TOށܒ!��DSP��JO1GӐ�#��_Pӱ�"�O�q����@�&KE�P�IR��ܔ�@ML}R��AP�Q^�Eh08��K�SYS�q"vK�PG2�BRK�B��߄�pY�=�d�����`AD������B�SOC���N��D?UMMY14�p�0�SV�PDE_OP��#SFSPD_O+VR-���C��ˢ&ΓOR٧3N]0ڦ�F�ڦ��OV��S!F��p���F+�|!����CC��1q"LCH�DL��RECOV(ʤc0��Wq@M����F��RO�#��Ȑ_+���� @0�e@VE}R�$OFSe@3CV/ �2WD�}�`�Z2���TR�!����E_FDO>�MB_CM���B��BL�bܒ#��adtVQR�$0p���G$�7�AM5��� eŤ��_M;��"'�<���8$CA��'�|E�8�8$HBK(1,���IO<�����QPPA������
���Ŋ����DVC_DBhC;��#"<Ѝ�D�S�1[ڤ�S�3[�^��ATIOq 1q�� ʡU�3���CABŐ�2�CvP��9P^��B���_� �SUB'CPU�ƐS�P  �M�)0NS�cM�"~r�$HW_C���U��S@��SA�A�pl_$UNITm�l_��AT���e�ƐCY{CLq�NECA����FLTR_2_�FIO�7(��)&B�L�Pқ/�.�_SCT�CF_`�Fb�l����|�FS(!E�e�CH�A�1��4�D°"3�RSD��$"}����;_Tb�PRO������ EMi_��a�8!�a !�a���DIR0�RAIL�ACI�)RMr�LO��C���Qq��#q��դ�PR=�S�A�C/�c 	��F�UNCq�0rRIN�P�Q�0��2�!RAC �B ��[����[WARn���BL�Aq�A�����DAk�\���L�D0���Q��qeq�TI"r��K��hPRIA�!r"AF��Pz!=�;��?,`(�RK���MǀI�!ÇDF_@B�%1n�L�M�FAq@HRDiY�4_�P@RS�A��0� �MULSE�@���a �8�ưt��  �1�$�1$1 �p����� x�*�EG00����!A1R���Ӧ�09�2,%ܲ 7�AXE��RO%B��WpA��_l-��CSY[�W!‎&S�'�WRU�/-1��@�SCTR������Eb� 	�%��J��AB�� ���&9�����OT�o0 	$��ARAY�s#2��Ԓ�	ё�FI@��$LI�NK|�qC1�a_��#���%kqj2XYZ��t;rq�3�C1)j2^8'0B��'��4����+ �3FI����7�q����'��_�Jˑ���O3�QOP�_�$;5���ATB�A�QBC��&�DU�β�&6��TURN ߁"r�E11:�p��9GFL�`_���* �@�5��*7��Ʊ 1�J� KŐM��&8��p�"r��ORQ�� a�(@#p=�j�g��#qXU�����mTOV	EtQ:�M��i���U��U��VW�Z�A�W b��T{�, ��@;�uQ ���P\�i��UuQ�We0�e�SERʑe�	��E� O���UdA as��4S�/7����AX��B�'q�� E1�e��i��irp�j J@�j�@�j�@�jP�j @ �j�!�f��i��i ��i��i��i�y �y�'y�7yTqHyoDEBU8�$3 2���qͲf2G + CAB����رnSVS�7� 
#�d��L� #�L��1W��1W�JAW� �AW��AW�QW�@!Ep@?D2�3LAB�2�9U4�Aӏ��C �  ERf�5� O� $�@_ A��!�PO��à�x0#�
�_MRAt�_� d � T���ٔERR����;T)Y&���I��V�0�cNz�TOQ�d�PL[ H�d�"��	��C!_ � pp`T)0���_V1Vr�aӔ����2ٛ2�E�����@�H�E���$W������V!��$�P��o�cI��aΣ�	 HELL_C�FG!� 5���B_BASq�SqR3��� a#QSb���1�%��U2��3��4��5���6��7��8���RaO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CO,. U�OUG�P~ ��`��m�������TPհ�_KAR�[@_�R�E*��P���|�Q�UE���uP����C�STOPI_AL 7�l�k0��h��]�l0GSEM�4�(�M4�66�TYN�SO���DIZ�~�A�����m�_TM�MANR�Q��k0E����$�KEYSWITCaH���m���HE��OBEAT��|�E- �LE~�����U��F�!Ĳ���B�O_HOuM=OGREFUP�PR&��y!� [�Cr��O��-ECOC�|�Ԯ0_IOCMWD<
�a�'k���� � Dh1���U�X���M�βgPgCFgORC��� ���m�OM.  � Q@�5(�U�#P, Q1��, 3��45�	�NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�Ѝ� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E��VP���UPDs� � �`NЦ�5�YS�LOt�� � �L��d���A�aTAp�0d��|�ALU:eLd�~�CUѰjgF!a�ID_L�ÑeHI��jI��$FILE1_���d��$2�f;SA>�� hO��`?E_BLCK��b|$��hD_CPUy�M�yA��c�o�d��Y�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA���J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP��_(�g����pr��{ `�`GROUw`���B��NFLI�C��f�REQUI;RE3�EBU��qB���w�2����p��x�q5�p�� \��/APPR��C}�Y��
ްEN٨CLO7��S_M��H����u�
�qu�� �`�MC�����9�_MG��C�Co��`M��в�N�BRKL�N�OL|�N�[�R��_CLINђ�|�=�J����Pܔ�����������������6ɵ�̲�8k�+��q����# ��
��q)��7�PATH3�L�BàL��H�wࡠ�J�CN�CA�Ғ�ڢB�IN�rUCV�4a��-C!�UM��Y,����aE�p����ʴ�~��PAYLOA���J2L`R_AN�q�Lpp���$��M�R_F2LSHR��N�LOԡ�R����`ׯ�ACRL_@G�ŒЛ� ��Hj`�߂$HM���FL[EXܣ�pJ�u� :���� ���������1�F1�V�j�@�R�d�v�������E����ȏ ڏ����"�4�q��� 6�M���~��U�g�y�$ယT��o�X��H� �����藕?����� ǟِݕ�ԕ�����%�7��JJ�� �� V�h�z���`A�T�採@�EL�� �S��J|�Ŝ�J�Ey�CTR��~�T�N��FQ��HAN/D_VB-���v`n�� $��F2M����ebSW�q�'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)�F�AW�Z`i�Aw�A���X X�'pi�Dw�Dʆ�Pf�G�p�)ST�k��!x��!N��DY �pנM�9$`%Ц�H� �H�c�׎���0� ��Pѵڵ���������PL���� ���1��R�6��QOASYMvř����v��J���cі�_SH>��ǺĤ�ED����������J�İ%�p�C�IDِ�_VI��!X�2PV_UN!IX�FThP�J��_R �5_Rc�cTz�pT�V�݀@���İ�߷��U $��������Hqpˢ3��aEN�3�DI����O4d�`NJ�� x g"IJAAȱz�aabp�coc�`pa�pdq�a� ��/OMME��� �b4�RqAT(`PT�@� S��a7�;�Ƞ�@�h��a�iT�@<� $DUMMY9Q��$PS_��RF�C�  S�v p�p���Pa� XƠ����STE���S�BRY�M21_V�F�8$SV_ER�F�O��LsdsCLR�JtA��Odb`O��p � D �$GLOBj�_LO���u�q�cAp�r�@�aSYS�qADR�``�`TCH  �� ,��ɩb�W7_NA���7���SR���l ���
*?�&Q� 0"?�;'?�I)?�Y)�� X���h���x������) ��Ռ�Ӷ�;��Ív��?��O�O�O�D�XS�CRE栘p��f��ST��s}y`����a/_HAΗq� TơgpTYP�b���G�aG�j��Od0IS_i䓀d�UEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI� m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��12�ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���>4�VSHIF��Nc�P�`ג�E�ȐyR����OSUR��=Wk`RADILѮ��_�a��:�9a��`a��r��LULQ$O�UTPUT_BM����IM�AB �@��rTILSC	O��C7��� ����&��3��A����q���m�I�2$G��V�pLe�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM���F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? �EaZABC%��  $�"R���
`�$$CLA}S������!�pE`� � VIRT8]��/ 0ABS�����1 5�� <  �!F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o �$6HZi{0-�A�XL�p��"�63  �{tIN��qztGPRE�����v�p��uLARMRECOV 9�rwt�NG�� .;	 A   �.�0�PPLIC��?�5�p�H�andlingT�ool o� 
�V7.50P/2�3-�  �Pfv��
��_SWt�w UP�!� x�#F0��t���A0v� 864��� �it�y� r�2 7wDA5�� �� ?Qf@��o��Noneisͅ�˰ ��T��~�!LAex>�E_l�V�uT��s9�UTO�"�Њt�y��?HGAPON
0g��1��Uh�D 1581����̟�ޟry����Q 1���p�,�蘦����;�@��q_��"{2 �c��.�H���D�HTTHKYX��"� -�?�Q���ɯۯ5��� �#�A�G�Y�k�}��� ����ſ׿1����� =�C�U�g�yϋϝϯ� ����-���	��9�?� Q�c�u߇ߙ߽߫��� )�����5�;�M�_� q�������%��� ��1�7�I�[�m�� ��������!���� -3EWi{�� ����)/ ASew���� /��/%/+/=/O/ a/s/�/�/�/�/?�/ �/?!?'?9?K?]?o? �?�?�?�?O�?�?�?0O#O]���TO�E��W�DO_CLEA�N��7��CNM  � �__�/_A_S_�DSPDgRYR�O��HIc��M@�O�_�_�_�_o o+o=oOoaoso�o�o0���pB��v �u����aX�t������9�PLUGG���G��U�WPRCvPB�@��_�orOr_7�/SEGF}�K[mw xq�O�O�����?rqLAP�_�~q� [�m��������Ǐُ�����!�3�x�TO�TAL�f yx�USWENU�p�� �H����B��RG_STRING 1u��
�Mn�S�5�
ȑ_ITE;M1Җ  n5��  ��$�6�H�Z�l�~� ������Ưد����� �2�D�I/O SIGNAL̕�Tryout� ModeӕI�np��Simul�atedבOu�t��OVER�R�P = 100�֒In cyc�l��בProg� Abor��ב~��StatusՓ�	Heartbe�atїMH F�aul��Aler'�W�E�W�i�{ύ���ϱ�������  �CΛ�A����8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|���WOR{pΛ��(� ������ ��$�6�H� Z�l�~���������������� 2PO ̛�X ��A{�� �����/ ASew�����SDEV[�o �#/5/G/Y/k/}/�/ �/�/�/�/�/�/??�1?C?U?g?y?PALTݠ1��z?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O_�?GRI�`ΛDQ �?_l_~_�_�_�_�_ �_�_�_o o2oDoVo�hozo�o�o�o2_l�R ��a\_�o"4F Xj|����� ����0�B�T��oPREG�>�� f� ��Ə؏���� �2� D�V�h�z��������ԟ���Z��$AR�G_��D ?	����;���  	$�Z�	[O�]O���Z�p�.�SBN_C�ONFIG �;�������CI�I_SAVE  �Z�����.�TC�ELLSETUP� ;�%HO�ME_IOZ�Z�%MOV_��
��REP�lU�(�UT�OBACKܠ���FRA:\z� \�z�Ǡ'`�z���ǡi�WINI�0z����n�MESSAG༠�ǡC���ODEC_D������%�O��4�n�PAUSX!��;� ((O >��ϞˈϾϬ����� �����*�`�N߄��rߨ߶�g�l TSK�  wͥ�_�q�UgPDT+��d!�~A�WSM_CF���;���'�-�G�RP 2:�?� �N�BŰA��%�XS�CRD1�1
7� �ĥĢ������ ����*�������r� ����������7���[� &8J\n��|*�t�GROUN�|UϩUP_NA��:�	t��_E�D�17�
 ��%-BCKED�T-�2�'K�`����-t�z��q�q�z���2 t1�����q�kp�(/��ED3/ ��/�.a/�/;/M/ED4�/t/)?�/.p?p?�/�/ED5`? ?�?<?.�?O�?�?ED6O�?qO�?.pMO�O'O9OED7�O `O_�O.�O\_�O�O�ED8L_,�_�^�-�_ oo_�_ED!9�_�_]o�_	-9o�oo%oCR_  9]�oF�o�k� � ?NO_DEL���GE_UNUSE���LAL_OU�T ����W?D_ABORﰨ~���pITR_RT�N��|NONS�k���˥CAM�_PARAM 1�;�!�
 8
�SONY XC-�56 23456�7890 �~��@���?��( А\�
����{����^�HR5pq�̹��ŏR57ڏ��Aff��K�OWA SC31�0M
�x�̆�d @<�
��� e�^��П\�����*�<��`�r�g�CE�_RIA_I�j!�=�F��}�vz� ��_LIU�Y]�����<���FB�GP 1��Ǯ�M�_�q��0�C*  ����CU1��9��@��G��Z�CR�C]��d��l��s��R�����U[Դm��v����}����� C���ő(�����=�HE�`ONFIǰ�B��G_PRI 1�{V���ߖϨϺ�����������CHK�PAUS�� 1K� ,!uD�V�@� z�dߞ߈ߚ��߾��� ���.��R�<�b���O��������_MOR�� =�^Biq-���� 	 �����*�@�N�`�������$?��q?;�;����)K��9�P���ça�-:���	�

��M���pU��ð��<��,~��D�B���튒)
m�c:cpmidb�g�f�:�0��0��¥�p�/��  ��p۰��� �s>_�  ���UX�?��p(�p�)Ug�/����Uf�M/w�O/�
D�EF l��s)��< buf.t�xts/�t/��ާ��)�	`�����=�L���*MC��1�����?43��1���t�īCz � BHH�CPUe�B�_B�y�;��>C����CnY
K�E?�{hD]^Dٿ�?r���1D���^�=G	���F��F���Cm	fF�O�OF�ΫY	���&�w�1���s�J��.�p��ዐ�BDLw�M@x8��1Ҩ�����g@D�p@�0E�Y�1X�E�Q�EJP F��E�F� G���=F^F E��� FB� H�,- Ge��H�3Y��:�  >�33 ���N~  n8�~@��#5Y�E>�ðA��Yo<#�
"Q ����+_�'RSMOF�S�p�.8��)T1>��DE ��F� 
Q��;�(P � B_<_��R��X��	op6C4P�Y
�s@ ]AQ�2s@CR�0B3�MaC{@@*c�w��UT�pFPROG %�z�o�o�igI�q���v��ldK�EY_TBL  ��&S�#� �	
��� !"#�$%&'()*+�,-./01i�:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������vq���͓���������������������������������耇���������������������p`LCK�l4�p`�`�STAT ��S_A�UTO_DO����5�INDT_ENB!���R�Q?�1��T2}�^�STOP�b���TRLr`LE�TE��Ċ_SCREEN �Z�kcsc��U���MMENU 1� �Y  < �l�oR�Y1�[���v� m���̟�����ٟ� 8��!�G���W�i��� �����ïկ��4�� �j�A�S���w����� 迿�ѿ����T�+� =�cϜ�sυ��ϩϻ� ������P�'�9߆� ]�o߼ߓߥ������ ��:��#�p�G�Y�� ����������$��� �3�l�C�U���y��� �������� ��	V�Y)�_MANUAyL��t�DBCO[��RIGڇ
�DBN�UM� ��B1 e
��PXWORK 1!�[�_U/�4FX�_AWA�Y�i�GCP r b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�(!mc�(&/~&lMZ�IdPx�@P@#ONTIM6ه� d�`&��
�e�MOTNE�ND�o�RECO_RD 1(�[g2�/{�O��!�/k y"?4?F?X?�(`?�? �/�??�?�?�?�?�? )O�?MO�?qO�O�O�O BO�O:O�O^O_%_7_ I_�Om_�O�_ _�_�_ �_�_Z_o~_3o�_Wo io{o�o�_�o o�oDo �o/�oS�oL �o����@�� �+�yV,�c�u�� ������Ϗ>�P��� ��;�&���q���򏧟 ��P�ȟ�^������ I�[����� ���$��6�������jTO�LERENCwB����L�͖ C�S_CFG )��/'dMC:�\U�L%04d.'CSV�� c��/#[A ��CH��z� �//.ɿ��(S�R�C_OUT *����SGN �+��"��#��09-MAY-20 11:330�15-JANp�0�:51+ P/Vt�ɞ�/.��f��pa�m��P�JPѲ��VE�RSION �Y�V2.0.�84,EFLOGI�C 1,� 	:ޠ=�ޠL���PROG_ENB���"p�ULSk' �����_WRST�JNK ��"fEM�O_OPT_SL� ?	�#
 ?	R575/#=ـ����0�B����TO  �ݵϗ��[V_F EX�d�%���PATH AY�A\������5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAU���z�^"MSWX�.D��4,#�Y�/�
!J�6%ZI�~m��$SBL_/FAUL(�0�9'/TDIA[�1<��� ���12�34567890
��P��HZl ~������� / /2/D/V/h/�� -P� ѩ�y� �/��6�/�/�/?? /?A?S?e?w?�?�?�?��?�?�?�?�,/�UM�P���� �AT�R���1OC@PME�l�OOY_TEMP?�È�3F���G��|DUNI��.�YN_BRK 2_��/�EMGDI_S�TA��]��ENC2_SCR 3�K7(_:_L_^_l&_��_�_�_�_)��C�A14_�/oo/oAoԢt�B�T5�K�� �o~ol�{_�o�o�o '9K]o�� �������#� 5��/V�h�z��л`~� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T���x���������ү �����,�>�P�b� t���������ο�� ��(�f�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������:� �2� D�V�h�z������ ������
��.�@�R� d�v������������ ��*<N`r ������� &8J\n�� ��������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?��?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O�__NoETMODoE 16�5�QW �d�X
X_�j_|Q�PRROR_PROG %GZ�%�@��_  �UTABLE  G[��?oo)oRjRR�SEV_NUM � �`WP��QQY`�Q_AUTO_ENB  �e�OS�T_NOna �7G[�QXb  �*��`��`��`��`d`+�`�o�o�o�d�HISUc�QOP�k_�ALM 18G[� �A��l�P+ �ok}�����o�_Nb�`  G[�a�R
�:PTCP_�VER !GZ!��_�$EXTLO�G_REQv蜁i\�SIZe�W�T�OL  �QDz�r�A W�_B�WD�p��xf́t�_�DI�� 9�5��d�T�QsRֆST�EP��:P�OP�_DOv�f�PF�ACTORY_T�UNwdM�EAT?URE :�5̀�rQHan�dlingToo�l �� \sfm�Englis�h Dictio�nary��rod�uAA Vi�s�� Masteyr����
EN̐�nalog I/yO����g.fd̐�uto Soft�ware Upd�ate  F O�R�matic �Backup��H�596,�gr�ound Edi�tޒ  1 H5�Cameraz�F��OPLGX��ell𜩐II)� X�ommՐsh�w���com��co����\tp���p�ane��  op�l��tyle s�elect��al� C��nJ�Ցon�itor��RDE���tr��Rel�iab𠧒6U�D?iagnos(��^��5528�u���heck Safety UIF���Enhanced� Rob Ser}v%�q ) "S��r�User Fr�[�����a��xt.� DIO �fi�G� sŢ��end�x�Err�LF� IpȐĳr됮� ��  !��FCT�N Menu`�v�-�ݡ���TP I�nېfac�  ER JGC�}pבk Exct��g��H558��i�gh-Spex�S�ki1�  2
�P��?���mmun;ic'�ons��&��l�ur�ې��ST� Ǡ��connz��2��TXPL���ncr�stru�����"FAT�KAREL Cmod. LE�uaG��545\��Runw-Ti��Env���d
!���ؠ+:+�s)�S/W��[��Licens�eZ��� 4T�0�o�gBook(Syvڐm)��H54O�MACROs,\¿/Offse��Loa�MH�������r, k�Mech�Stop Proyt���� lic/�{MiвShif����ɒMixx��)�xStS�Mod�e Switchn�� R5W�Mo�z:�.�� 74 ����g��K�2h�ulti-T=�M����LN (Po=s�Regiڑ�������d�ݐt Fu�n�ǩ�.�����N�um~����� ln�e��ᝰ Adj�up�����  -{ W��tatuw����T�RDM�z�ot��scove U�9����3Ѓ�uest 4�92�*�o�����6�2;�SNPX b< ���8 J7`����Libr��J�48����ӗ� �Ԅ�
�6�O�� Parts� in VCCMt�32���	�{Ѥ�oJ990��/I�� 2 P��TMI�LIB��H���P��AccD�L�
�TE$TX�ۨ�a�p1S�Te����p�key��wգ�d���Unexc�eptx�motn`Z��������єƉ� O���� 9�0J�єSP CS�XC<�f��Ҟ� �Py�We}���PR�I�>vr�t�m�en�� ��i�Pɰa�����vG�rid�play`��v��0�)�H1��M-10iA(B�201 �2\� �0\k/�Asci�i�l�Т�ɐ/�C�ol��ԑGuar&� 
�� /P-�ޠ�"K��st{Pa�t ��!S�Cyc8�҂�orie�⑻IF8�ata- q�uҐ�� ƶ��mH�574��RL��a�m���Pb�HMI De3�(b�����PCϺ�Passswo+!��"PE? cSp$�[���tp��.� ven��Tw�N��p�YELLOW� BOE	k$ArcN��vis��3*��n0WeldW�ci�al�7�V#t�O�p����1y� 2zF�a�portN�(�p�T1�T� ��� ��xy]�&TX��tw�igj�1� �b� ct\�JP�N ARCPSU� PR��oݲOL�� Sup�2fil� &PAɰאcro�� "PM(�����O$SS� eвte�x�� r���=�t��ssagT��P��P@�Ȱ�锱��rtW��H'>r�dspn��n1
t��!� z ��asc�bin4psyn���+Aj�M HE�L�NCL VI�S PKGS PwLOA`�MB ��,�4VW�RIP�E GET_VA�R FIE 3\�t��FL[�OOL�: ADD R7�29.FD \j�8'�CsQ�QE��D�VvQ�sQNO W�TWTE��}PD � �^��biRFO;R ��ECTn�`���ALSE AL�AfPCPMO-1�30  M" #�h�D: HANG FROMmP�AQ�fr��R709 �DRAM AVA�ILCHECKS�O!��sQVPCS �SU�@LIMCH�K Q +P~dFF �POS��F�Q R�5938-1?2 CHARY�0�PROGRA �W�SAVEN`AM]E�P.SV��7��$En*��p?FU�{��TRC|� SHA�DV0UPDAT �KCJўRSTAT�I�`�P MUCH� y�1��IMQ �MOTN-003���}�ROBOGU�IDE DAUG�H�a���*�tou�����I� Šhd�A�TH�PepMOVE�T�ǔVMXPA�CK MAY A�SSERT�D��Y�CLfqTA�rBE COR vr*Q�3rAN�pRC O�PTIONSJ1v�r̐PSH-17�1Z@x�tcǠS�U1�1Hp^9R!�Q�`_�T�P��'�j�d�{tby app �wa 5I�~d�PHqI���p�aTEL��MXSPD TB$5bLu 1��UB6@�q�ENJ`CE2�61ꏠp��s	�mayc n�0� R6{��R� �Rtraff\)�� 40*�p���fr��sysva�r scr J78��cj`DJU��b�H V��Q/�PSE�T ERR`J` �68��PNDAN�T SCREEN? UNREA��'�J`D�pPA���pR�`IO 1���PF�I�pB�pGROUN�PD��G��R�P�Q>nRSVIP !p�a��PDIGIT VgERS�r}BLo�U�EWϕ P06 9 �!��MAGp�abZV�DI�`� �SSUE�ܰ�EPLAN JOT`O DEL�pݡ#Zz�@D͐CALLOb��Q ph��R�QIwPND��IMG��R719��MNT]/�PES �pVL�c��Hol�0Cq��N�tPG:�`C�M��canΠ��pg.�v�S: 3D m~K�view d�`� �p��ea7У�b�� of �Py���A�NNOT ACCESS M��Ɓ*��t4s a��lo�k��Flex/:ڈRw!mo?�PA�?�-�����`n�pa� SNBPJ AUTO-�06f�����TB��PIABLE�1q 636��PLgN: RG$�pl;p�NWFMDB�VI|���tWIT 9x�:0@o��Qui#0�Ҿ�PN RRS?pU�SB�� t & _remov�@ )��_��&AxEPFT_f=� 7<`�pP:�OS-144 ���h s�g��@OS�T� � CRAS�H DU 9���$P�pW� .$���LOGIN��8�&�J��6b046 �issue 6 �Jg��: Slo�w �st��c (Hos`�c���`�IL`IMPRWtS?POT:Wh:0�T�STYW ./�V�MGR�h�T0CA]T��hos��E�q���� �O�S:N+pRTU' k�-S�Y ����E:��pv@8�2�� t\hߐ��9m ��all��0�s  $�H� WA͐���3 CNT0 �T�� WroU�a�larm���0s�d � �0SE1���r R{�OMEBp���nK� 55��REà�SEst��g   �  �KANJ�I�no���IN�ISITALIZ-p�dn1weρ<���dr�� lx`�S�CII L�fa_ils w�� ��`�YSTEa���o���Pv� IIH���1�W�Gro>Pm ol\wpSh@�P��~Ϡn cflxL@�АWRI �OF �Lq��p?�F�up���de-rela��d "APo S�Y�ch�Abetw}e:0IND t0�$gbDO���r� �`�GigE�#operabilf  PAbHi�H`��c��lead�\et�f�Ps�r�OS p030�&: fig��GLA )P ��i����7Np tpswZx�B��If�g�������5aE�a E�XCE#dU�_�tPC�LOS��"robV�NTdpFaU�c��!���PNIO /V750�Q1��Q�a��DB ��P �M�+P�QED�DEyT��-� \rk���ONLINEhSBUGIQ ߔĠi`Z��IB�S apABC JARKYFqr� ���0MIL�`*� R�pNД �p0WGAR��D*pRМ�P�"! jK�0cT��P�Hl#n�a�ZE� V�� TASK�$VP2(�4`
�!p�$�P�`WIBPKk05�!FȐB/���BUSY RUNN�� "�򁐈���R-p�LO�N�D;IVY�CUL��gfsfoaBW� p���30	V��ˠ�IT`�a505.��@OF�UNEXH�P1b�af�@�E���SVEMG� NM�Lq� D0pCC_�SAFEX 0c�08�"qD �PET�`N�@�#J87����RPsP�A'�M�K�`�K�H GUNC{HG۔MECH�p�Mc� T�  y,� g@�$ ORY LEAKA�;�ޢGSPEm�Ja��V�t�GRIܱ�@�C7TLN�TRk�Fp�epR�j50�ENF-`IN�����p �`0�Ǒk!��T3/dq.o�STO�0A�#�L�p �0�@�Q�АaY�&�;pb1TO8pP�s���FB�@Yp`&�`DU��aO�sup$k�t4 � P�F� B�nf�Q�PSVGN�-1��V�SRSR)J�UP�a2�Q�#<D�q l O��Q?BRKCTR5Ұ��|"-�r�<pc�j!I{NVP�D ZO� ���T`h#�Q�cHse�t,|D��"DUA�L� w�2*BRVO_117 A]�TN�p�t�+bTa2473�0�q.?��sAUz�i��B�complet�e��604.�{ -�`hanc�U� F��e8��  ��npJtPd!q�ܱ`��� 5h59	6p�!5d�� "p�P�P�Q�0�P2�p�A� HxP��R(}\xPe� %aʰI���E��1���p� j  �� xStO�^t �A�AxP��q 5 sig��a��"AC;a��
��bCexPb_p��.�pc]l<bHbcb_�circ~h<n�`tl1�~`xP`o�dxP�b,]o2�� �cb�c�i|xP�jupfrm�d8xP�o�`exe�a�o<FdxPtped}o��|u`�cptlibxzxP�lcr�xrxP\blsazEdxP_fm�}gcxP�x���o|�sp�o�mc(��ob_�jzop�u6�wf(��t��wms�1q��csld�)��jmc�o�\�n��nuhЕ��|s1t�e��>�pl�qp��iwck���uvf�0uߒ��lvisn��CgaculwQ
}E F  ! Fc�.fd�Qv�� q�w���Data A�cquisi��nxF�|1�RR631`���TR�QDMCM Z�2�P75H�1�P�583xP1��71֫�59`�5�P57@<PxP�Q����(����Q��o pxP!daq\�oA��@��� ge/�etdm~s�"DMER"؟�,�pgdD���.�mp���-��qaq.<ጡ�xPmo��h���f�{�u�`13��MACROs, SksaCff�@z����03�SQR�Q(��Q6��1�Q9ӡ�R�ZSh��PxP�J643�@7ؠ6X�P�@�PRS�@����e �Q�UС PIK��Q52 PTLC��W��xP3 (��p/O��!�Pn ��xP5��03\sf�mnmc "MNCMCq�<��Q��\$AcX�FM���ci,� ��X����cdpq+�
�sk�SK�xP�SH560,P��,��y�refp "R#EFp�d�A�jxP	�of�OFc�<gy�to�TO_���������+je�u>��caxis2�xP�E�\�e�q"ISD�Tc��]�prax ��MN��u�b�isde܃h�\�w��xP! isbaskic��B� P]�ޔQAxes�R6p������.�(Ba�Q�ess��xP����2�D�@�z�atis���(�{�����4~��m��FMc�u�x{�
ѩ�MNIS�� ݝ����x����ٺ���x� j75��D�evic�� In?terfac�R��QJ754��� xP�Ne`��xP����2�б����dn� "DNE���
�tpdnui5U1I��ݝ	bd�bP|�q_rsofO�b
dv_aro���u�����stchkc��z	 �(}onl��G!ffL+H�J(��"l"/�n�b��z�Ohamp��T�C�!i�a"�59��S�q��0 (�+P�o�u��!2��xpc_2pc�chm��CHMP8_�|8бpevws��8�2쳌pcsF��#�C SenxPac�ro�U·�-�R6 �Pd�xPk�����p��qgT�L��1d M�2 `��8�1c4ԡ�3 q;em��GEM,\i|(��Dgesnd�5����H{�}Ha�@sy���c�Isu�xD��Fmd��I��7�4����u���AccuCaAl�P�4� ��ɢ7ޠ�B0��6+6f�6���99\aFF q�S( �U��2�
X�p�!�Bd��cb_�SaUL��  �� ?�ܖ�to��otplu?s\tsrnغ�qb�Wp��t���1���Tool (N. A.)�[K�7�Z�(P�m����b�fcls� k94�"�K4p��qtpap� "PS9H�stpswo��p�L7��t\�q����D� yt5�4�q��w�q���� �M�uk��rkey����s��}t�s�featu6�EA��� cf)t\Xq������d�h5���LaRC0�md�!�587���aR�(����2V���8c?u3l\�pa3}H�&r-�Xu���1t,�� �q "�q�O t��~,���{�/��1c�}����y�p�r�� 5���S�XAg�-�y��ށWj874�- �iRVis���Queu�� Ƒ�-�6�1���(����u����tӑ����
�t�pvtsn "V�TSN�3C�+�� v�\pRDV����*�p�rdq\�Q�&�vstk=P�������nm&_�դ�clrqqν���get� TX��Bd���aoQϿ�0qstr�D[� ¡�t�p'Z����np8v��@�enlIP0���D!x�'�|���sc ߸��tvo/��2�q���vb���� q���!���h]��(�� Contro�l�PRAX�P5ξ�556�A@59��P56.@56@5�A�J69$@98�2 J552 IDVR7�hqA���16��H���La��� ��Xe�frlp�arm.f�FRL�am��C9�@(F�����w6{��x�A��QJ643��� 50�0LSE�
_pVAR $S�GSYSC��RS_UNITS �P�2�4tA�TX.$�VNUM_OLD� 5�1�xP{�5�0+�"�` Funct���5tA� }��`#@�`3�a0�cڂ��19���@H5נ� �P���(�A���� ۶}����ֻ}��bcPRb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`d���1���96������%C�� Aف��J�bIncr�	�����\���1o5qn=i4�MNINp	xP��`���!��Hour  �� 2�21 �AAVM����0 ��TUP ���J545 ���6162�VCAM  (�CLIO ��R6�N2�MgSC "P �?STYL�C��28~ 13\�N�RE "FHRM� SCH^�D�CSU%ORSR� {b�04 ��EIOC�1 j� 542 � os�| � egistP�����7�1��MASK�9�34"7 ��OCSO ��"3�8�b�2���� 0 HBh��� 4�"39N�� Re�� �LC{HK
%OPLG%z��3"%MHCR.%�MC  ; 4? ��6m dPI�54�sn� DSW%MD� 9pQ�K!637�0�0dp"�1�Р"4 ��6<27 CTN �K � 5 ���"7���<25�%/�T�%F'RDM� �Sg!��930 FB( N�BA�P� ( HLB�  Men�SMx$@jB( PVC ���20v��2HTC��CTMIL���\@PAC 16�U�hAJ`SAI \@E�LN��<29s��UECK �b�@FgRM �b�OR����IPL��Rk0C�SXC ���VV�FnaTg@HTTP9 �!26 ���G�@obIGU=I"%IPGS�r� H863 qb�!�0�7r�!34 �r�84 \so`! Qx`&CC3 Fb�21�!�96 rb!51 L���!53R% 1!Qs3!��~�.p"9js� VATFUJ77Q5"��pLR6^RP�wWSMjUCTO�@bxT58 F!80����1XY ta3!77s0 ��885�UOL  GTSo
�{`� LCM �r| T3SS�EfP6 W�\@�CPE `��0V1R� l�QNL"��@�001 imrb�c3 =�b�0���0ƒ`6 w�b-P- �R-�b8n@5EW�b9 �Ґa� ���b��`ׁ�b2 200I0��`3��`4*5��`5!�c�#$�`7�.%�`8 h605v? U0�@B6E"a�Rp7� !Pr8 �t�a@�tr2 i�B/�1vp3�vp5I Ȃtr9Σ�a4@9-p�r3 F��r�5&�re`u��r7 ���r8�U�p9 \�h738�a�R2�D7"�1f��2�&�7� �3 7iC��4>w5Ip�Or'60 C�L�1bEN�4 I�pyL�uPИ�@N�-PJ8�N�8NeN�9 H�r`�EE�b7]�|���8���ࠂ9 2��a`�0�qЂ5�%U09'7 0��@1�0����1 (�q�3 5R���0���mp U��0�0�7*��H@(q�\P"RB6�q124�b;��@����@06� x�3 �pB/x�u ��x�6_ H606�a1� <��7 6 ��x�p�b155 �����7jUU162 L�3 g��4*�65 2e "_���P�4U1`���B1����`0'�174 �q��P�E186 3R ��P�7 ��P��8&�3 (�907 B/�s191���Θ@202��6 a3���A�RU2� <d��2 b2h`���4�᪂2�4���1I9v Q�2��u2d��Tpt2� ��H�a2�hP�$�5���!U2��p�p
�2�p��@5��0-@��8 @�9F��TX@�� �e5�`'rb26Af�2^R�a@�2Kp��1y�b5Hp�`
�5�0@�gqGA����a52ѐ�Ḳ6��60ہ5� ׁ2Ҹ�8�E��9�EU5@ٰ\�q5hQ`S�2ޖ5�p\w�۲�p�J �-P��5�p1\�t�H�4��PCH�7j��phiw�@��P��x��559 ld u� P�D���Q�@������� �`.��P>�8�581�"�q5�8�!AM۲T�A ;iC�a589��@�x����5 �a��1�2׀0.�1���,�2p����,�!P\h8��RLp ��,�7��6�0�840\� ANRS 0C}A��p���{��ran��FRA��Д�е���A %���ѹ�Ҍ����� (����Ќ���З� ��������ь����B$�G��1��ը���������� x9S�`q�  ������`64��M��iC?/50T-H����0��*��)p46��� �C��N����m75s֐� Sp��b�46��v����ГM-71?�7�З����42������C��-�а�70�r�	E��/h����O�$��rD���c7c7�C�q��Ѕ���L���/��2\imm7c7�g������`���(��e��� ��"�������a �r��c�T,�Ѿ�" ��,�� ��x�Ex�m77t����k����5�����)�iC��-HS-� B
�_�>���+�Т�7@U�]���Mh7��s��7������-�9?�/260L_@������Q����h���]�9pA/@����q�S�хx���h621��c��92������.�)92c0�g$ �@�����)$��5$���pylH"O"
�2�1���t?�350 ����p��$�
�� �350!����0��9�U/0\m=9��M9A3��(4%� s��3M$���X%u���"him9@8J3����� i d�"m4~�103p�� ����h794̂�&R���H�0����\��� g�5AU��՜��0���*2��00��#06��АՃ�է!07{r ��������k�@�@����EP�# ������?��#!��;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?�ҽCD�25L����0:�"l�2BL
#��B��\20�2_�r�r e���X��1��N���H�A@��z��`C�p`U��`��04��$DyA�\�`fQ���sU���\�5  ���� p�3^t��<$85����+P=�ab1l��1#LT��lA8�!uD�nE(�20T��J8�1 e�bH85���b4�Ռ�5[�16Bs ��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3�  ��b�s��-`�_W8�_����6Id	$�X5�1�U85��R�p6S����/�/ +q�!�q��`�6o��q5m[o)�m6sW���Q�?��set0�6p ��3%H�5��10p$����g/�Jr�H��  ��A�856����F2�� ���p/2��h� ��܅�✐)�5��̑`v��(��m6��BY�H�ѝ̑m�6�Ҕ���a6�DM����-S�+��H2���� �Ҽ�� �r̑���`����l���p1����F���2�\t6h T6H����Ҝ� 'Vl���ᜐ�V7᠜�/����;3A7���p~S��������4��`圐�V���!3
��2�PM[��%ܖnO�chn��vel5�����Vq���_ar�p#��̑�.���2l_hemq$�.�'�6415���5���?�@���F�����5g�L�ј[���1����1����M7NU��М��eʾ����u"q$D;��-�4��3&H�f�c�Ĝ�h���� ��u���㜐���ZS�!ܑ4���M-����S�$̑�ք �� 0��<�����07shJ�H�v�À� sF��S*󜐳���̑@���vl�3�A�T�#���QȚ�Te��q�prX����T@75j�5�d d�̑1�(UL�&�(�,����0�\�?���̑�a�� xSt���a�e�w�2��(�	�2�C��A/���\��+p�����21 (ܱ�CL S���� B̺��7F���?�<�lơ1L����c� Č��u9�0����e/q��O���9�K��r9 (��,�Rs����5�G�m20c ��i��w�2��:�0`�$��2�2l�0�k� X�S� ,�ι2��O�4��1!41w���y2T@� _std��G�y� �ң�H� jdgm����w0\�  �1L���	�P�~�W*�b��t 5�����J�3�,���E{�������L��5	\L��3�L�|#~���~!���4�#��O����h�L6A��������2璥���4�4�����[6\j4s��·���#��ol�E"w�8Pk����� ?0xj�H1�1Rr�>�l�]�2a�2Aw�$P ��2��|41�8�� ˡ��{� �%�A<��� +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K� R��ˑb�W���Fs� ��)�ѐ�!���a�1�����5��16�1�6C��C����0\imBQ��d����b���\B5�-���DiL���O�_�<ѠPEtL�E�RH�ZǠPg���am1l��u��� ̑�b�<����<�$�T�̑�F����Ȋ�Dpb��X"�ᒢ���p� ���^t��9�0\� j97�1\kckrcf�J�F�s�����c��e? "CTME�r������!�a�`main�.[��g�`run}�_vc�#0�w�1�Oܕ_u����bct�me��Ӧ�`ܑ�j�735�- KA�REL Use {�U���J��1���p� Ȗ�9�B@@��L�9��7j[��atk208 "�K��Kя��\��9���a��̹����cK�RC�a�o ��kc �qJ�&s�����Grſ �fsD��:y��s��Af1X\j|хrdtB�2, ��`.v�q��� �sǑIf�Wfj5�2�TKQuto �Set��J� H�5K536(�93�2���91�58(�94�BA�1(�74O,A~$�(TCP Ak����/�)Y� �\�tpqtool.�v��v���! c�onre;a#�Co�ntrol Re�ble��CNRE(�T�<�4�2���D�8)���S�552��q(g�� (򭂯4X��cOux�\sfuts�UTS`�i������t�棂��? q6�T�!�SA OO+D6���������,!��6c+� i\gt�t6i��I0�TW8 ���la��vo58�o�bFå��i�Xh��!Xk�0Y�!8\m6e�!6#EC���v��6���� �����<16�A���A�6s����U�g˰T|ώ���r1�qR��˔Z4�T�����,#�eZp)g����@<ONO0���uJ��tCR�;��F�a� xSt��f��prdsuc#hk �1��2&&?���t��*D%$�r(��✑�娟:r��'�sp�qO��<scrc�xC�\At�trldJ�"o�\�V����P�aylo�nficrm�l�!�87��@7��A�3ad� ! �?ވI�?plQ��3��3"�q��x pl�`���d7��l�calC�uDu���;��mov�����OinitX�:s8O���a�r4 ��r67�A4|�e Gene�ratiڲ���7�g2q$��g R� G(Sh��c ,|�"bE��$Ԓ\�(:�"��4��4�4�. sg��5�F$d�6"e�!p "S�HAP�TQ ngcr pGC�a(�&x"� ��"GDA¶&��r6�"aW�/�$dataX:s�"�tpad��[q�%tput;a__O7;a�Po8�1�yl+s�r�?��:�#�?�5x�?�:c O�:y O�:�IO�	s`O%g�qǒ�?�@p0\��"o�j92;!��Ppl.Coll{is�QSkip#� �@5��@J��D��@\�ވ�C@X�7��7��|s2��ptcl�s�LS�DU�k<?�\_ ets�`�< \�Q��@���`2dcKqQ�FC;��1J,�n��` (��"4eN����T�{�� �'j(�c�q���/I��aȁ��̠H������зa�e\m�cclmt "C�LM�/��� mat�e\��lmpALaM�?>p7qmc?����2vm�q��%�3s���_sv90�_x_Gmsu�2L^v_� K�o�{in�8(3r><�c_logr���rtrcW� "�v_3�~yc���d�<�te��de�r$cCe� Fiρ�R��Q�?�>l�enter߄|���(Sd��1�TXj�+fK�r�a99sQ�9+�5�r\tq~\� "FNDR�}��STDn$�LANG�Pgui��D⠓�S�������sp�!ğ֙uf�ҝ�s����$�����e+�=����������������w�H�r\�fn_�ϣ��$`x�t�cpma��- T�CP�����R63�8 R�Ҡ��38��M7p,���Ӡ� $Ӡ�8p0Р�VS,�>�tk��99�a��B3 ���PզԠ��D�2�����UI��t���hqB� ��8��������p����re�ȿ��exe @4φ�B���e38�ԡ�G�rmpWXφ�var@�φ�3N��ψ��vx�!ҡ��q��RBT $c�OPTN ask� E0��1�R M{AS0�H593/՟96 H50�i�480�5�H0��mԢQ�K��7�0�g�P�l�h0ԧ�2�OR�DP��@"��t\mas��0�a��"��������k�գR�����ӹ`m��b��7�.If��u�d��r��splayD�E���|1w�UPDT Ub���887 (��D	i{���v�Ӛ�Ԛ‧���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q`�䗣�#��К�`2�� vlv������$�>�b���! <S��Easy/К�Util��룙�5�11 J�����R�7 ��Nor֠��i�nc),<6Q�� ��`c��"4�[���9�86FVRx So����q�nd6����P ��4�a\ (��
  ��������d��K�bd�Z���men7���-7 Me`tyFњ�Fb�0�TUa�577?i3R��\�5�u?��!� �n���f������l\mh�Ц�űE|�hmn�	��<\�O���e�1�� �l!��y��Ù�\|p����B���Ћmh�@��:.a G!���/�t�55�6�0�!X�l�.us��Y/>k)ensubL���eK�h�� �B\1 ;5g?y?�?�?D��?*�rm�p�?Ktbox O2K|?�G��C?�A%ds���?1ӛ#� �TR��/��P�4B �`�U�P�V�P"�Q�P�0�U�PO��P�"�T3��U�P�f�Pk"�2}�4��T�P�f�P2�"�Q5 �S�Q���R?Ă�Q3t.�P׀al��P+�OP517��IN0a��Q(}g��P'ESTf3ua�PB�l�ig�h�6�aq��P � xS�΅`  n�0mbusmpP�Q969g�C69�Qq��P0�ba�Ap�@Q� BOX8��,>vche�s��>vetu㒣=wffse�3���]�`;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q<twaNǂ tp�Q҄Ta�ror Reco�v�b�O�P�642����a�q��a�f�QErǃ�Qry���`�P'�T�`�aar�������	{'�pak971��71��m���>�pjot��PXch��C�1�adb -�a;il��nag���b�QR629�a�Q����b�P  �
�  �P��$$�CL[q ����������$��PS_DIGIT\���"� !�4�F�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv�����@��*璬1�:PRODUCT��Q0\PGSTK�bV,n�99��\���$F�EAT_INDE�X��~��� 搠ILEC�OMP ;���)��"��SET�UP2 <����  N �!�_AP2BC�K 1=� G �)}6/E+%,/i/��W/�/~+/ �/O/�/s/�/?�/>? �/b?t??�?'?�?�? ]?�?�?O(O�?LO�? pO�?}O�O5O�OYO�O  _�O$_�OH_Z_�O~_ _�_�_C_�_g_�_�_ 	o2o�_Vo�_zo�oo �o?o�o�ouo
�o. @�od�o��� M�q���<�� `�r����%���̏[� ������!�J�ُn� ������3�ȟW���� ��"���F�X��|�� ��/���֯e������ 0���T��x������ =�ҿ�s�ϗ�,ϻ��9�b�� P/ }2) *.VRi���!�*����������PC�7�!��FR6:"�c��χ��T��߽�L�����ܮx���*#.F��>� �	N�,��k��ߏ��STM� �����Qа����!�iPenda�nt Panel���H��F���4���8���GIF��������u����JPG&P��<�����	PANEL1'.DT��������2�Y� G��
3w�@����//�
4��a/�O///�/�
�TPEINS.XSML�/���\�/��/�!Custom� Toolbar�?�PASSW�ORD/�FR�S:\R?? %�Password Config�? ��?k?�?OH�6O�? ZOlO�?�OO�O�OUO �OyO_�O�OD_�Oh_ �Oa_�_-_�_Q_�_�_ �_o�_@oRo�_voo �o)o;o�o_o�o�o�o *�oN�or�� 7��m��&�� �\�����y���E� ڏi������4�ÏX� j��������A�S�� w�����B�џf��� ����+���O������ ���>�ͯ߯t���� '���ο]�򿁿�(� ��L�ۿpς�Ϧ�5� ��Y�k� ߏ�$߳�� Z���~�ߢߴ�C��� g�����2���V��� �ߌ���?����u� 
���.�@���d���� ��)���M���q��� ��<��5r�% ��[�&� J�n��3� W���"/�F/X/ �|//�/�/A/�/e/ �/�/�/0?�/T?�/M? �??�?=?�?�?s?O �?,O>O�?bO�?�OO 'O�OKO�OoO�O_�O :_�O^_p_�O�_#_�_ �_Y_�_}_o�_�_Ho�)f�$FILE_�DGBCK 1=���5`��� ( �)�
SUMMARY�.DGRo�\MD�:�o�o
`Di�ag Summa�ry�o�Z
CONSLOG�o�o�a
�J�aConso?le logK�[��`MEMCHECCK@'�o�^q�Memory D�ata��W��)�qHADOW����P��sSh�adow Cha�ngesS�-c-��)	FTP=Ъ�9����w`qmment TBD׏��W0<�)ET?HERNET̏�^��q�Z��aEth�ernet bpf�iguratio�n[��P��DCSV�RFˏ��Ïܟ�q�%�� veri?fy allߟ-c�1PY���DIF�Fԟ��̟a��p%=��diffc����q��1X�?�Q��c ����X��CHGD��¯ԯi�B�px��� ���2`�8G�Y�� ��� �GD��ʿܿq��pq���Ϥ�FY3h�8O�a��� ��(�GD������y��p��ϡ�0�UPDATES.�Ц��[?FRS:\������aUpdate?s List���k�PSRBWLD.CM.��\��B���_pPS_ROBOWEL���_����o ��,o!�3���W���{� 
�t���@���d��� ��/��Se��� ��N�r�  =�a�r�&� J���/�9/K/ �o/��/"/�/�/X/ �/|/�/#?�/G?�/k? }??�?0?�?�?f?�? �?O�?OUO�?yOO �O�O>O�ObO�O	_�O -_�OQ_c_�O�__�_ :_�_�_p_o�_o;o �__o�_�o�o$o�oHo �o�o~o�o7�o0 m�o� ��V� z�!��E��i�{� 
���.�ÏR������� ���.�S��w���� ��<�џ`������+� ��O�ޟH������8�ຯ߯n����$FoILE_��PR����������� �MDO?NLY 1=4��? 
 ���w� į��诨�ѿ������ �+Ϻ�O�޿sυ�� ��8�����n�ߒ�'� ��4�]��ρ�ߥ߷� F���j�����5��� Y�k��ߏ���B��� ��x����1�C���g� �����,���P����� ����?��Lu�?VISBCKR�<�>a�*.VD|�>4 FR:\���4 Visio�n VD file� :LbpZ �#��Y�}/ $/�H/�l/�/�/ 1/�/�/�/�/�/ ?�/ 1?V?�/z?	?�?�??? �?c?�?�?�?.O�?RO dOO�OO�O;O�O�O qO_�O*_<_�O`_�O��__%_�_�MR_�GRP 1>4��L�UC4  B�P	 ]�ol�`�*u����RHB ���2 ��� ��� ���He�Y�Q `orkbIh�oJd�o�S�c�o�oL:R��LE��Jr�I�F�5U�aS'�Q�o�o F
��F8_�E����.���9���>���}A'��A}�lq�?�o�A}�q�xq}E�� F�@ �r�d�a}J���NJk�H9��Hu��F!���IP�s}?��`�.9�<9��896�C'6<,6�\b�}B���Bǥ�Casd�B�n;B���B��{-�&W�A��B�-�A��VAƯ�A�e���,fp�PA�����|�ݏx����%���p�A6Β@U��{ �v�a�������П�� ��ߟ��<���i{~BH�P>p�``�Q��QA@(�K���ï��T
6�P=��P��\�˯�o�oB��P5���@�33�@���4�m�,�@U�UU��U�~w�>u?.�?!x�^���ֿ���3��=[�z�=�̽=�V6<�=�=��=$q��~���@8�i7G���8�D�8?@9!�7ϥ��@Ϣ���cD�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p���������^��� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__>���  DE_�Hly_�\@@m_B�=��vR/��I�O�SMT
�G�SUoo&o�RHOSTC�19H�I� ��zM�SM�l[�bo�	127.�0�`1�o  e �o�o�o#z�oF�Xj|�l60s	a�nonymous�������)2(ao�&�&��o� x��o������ҏ�3 ��,�>�a�O���� ������Ο�U%�7�I� �]����f�x����� ���ү����+�i� {�P�b�t�������� ����S�(�:�L� ^ϭ�oϔϦϸ���� ��=��$�6�H�Zߩ� ��Ϳs���������� � �2���V�h�z�� �߰���������
�� k�}ߏߡߣ���߬� ��������C�*< Nq�_����� �-�?�Q�c�eJ�� n������ �/"/E�X/j/|/ �/�/�%'/? [0?B?T?f?x?��? �?�?�?�??E/W/,O�>OPObO�KDaENT� 1I�K P!\�?�O  �P�O �O�O�O�O#_�OG_
_ S_._|_�_d_�_�_�_ �_o�_1o�_ogo*o �oNo�oro�o�o�o	 �o-�oQu8n �������� #��L�q�4���X��� |�ݏ���ď֏7����[���B�QUICC0��h�z�۟��A1ܟ��ʟ+���2,����{�!ROU�TER|�X�j�˯!?PCJOG̯���!192.168.0.10���}GNAME !��J!ROBOT��vNS_CFG �1H�I ��Auto-s�tarted�$FTP�/���/�? ޿#?��&�8�JϏ? nπϒϤ�ǿ��[��� ���"�4ߵ&������ ����濜�������� ��'�9�K�]�o��� �����������/�/ �/G���k��ߏ����� ��������1T� ��Py����� "�4�	H-|�Qc u�VD���� /�;/M/_/q/�/ ����/
/�/>? %?7?I?[?*/?�?�? �?�/�?l?�?O!O3O EO�/�/�/�/�?�O ? �O�O�O__�?A_S_ e_w_�O4_._�_�_�_ �_oVOhOzO�O�_so �O�o�o�o�o�o�_ '9Kno�o�� ���o*o<oNoP 5��oY�k�}�����p ŏ׏����0���C��U�g�y���_�T_ERR J;������PDUSIZ  ���^P����>~ٕWRD ?z����  guest���+��=�O�a�s�*�SCD�MNGRP 2K�z�Ð���۠\��K�� 	�P01.14 �8�q   y���B  �  ;����{ �����������������������~ �`ǟI�4�m�X�|���  i  _�  
���� �����+��������
���lZ�.x����"�!l�ڲ۰s�d��������_GROU���L�� ��	웡۠07K�QUPOD  ���P�V��TYg������TTP_AUTH� 1M�� <!�iPendan����<�_�!KAREL:*�����KC%�5�G���VISION SETZ���|��Ҽߪ�������� �
�W�.�@��d�v����CTRL Nи������
 �.FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@oG %j%@�_MOV�u����MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�5�
�4-�8��"�۵M�O~q_DCd~�1P�L_NAME �!<u� �!D�efault P�ersonali�ty (from� FD) �4RR�2k! 1j)TE�X)TH��!�AX d�?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�Ox2-?�O�O�O__@0_B_T_f_x_�b<�O �_�_�_�_�_�_o o�2oDoVoho&xRj" �1o�)&0\�b,� �9��b�a �@D�  �a?�ľc�a?�`�a�aA'�6�ew;�	�l�b	 ��xJp���`�`	p �<w �(p� �.r�� K�K ���K=*�J����J���JV�`�kq`q�P�x��|� @j�@T;;f�r�f�q�a�crs�I�� چ�p���p�r�ph}��3��´  Æ�>��ph�`z���꜖"�3Jm�q� H�N���ac��$�dw�� ~ �  P� �Q� �� |  �а�m�Əi}	'�� � �I�� �  ��ވ�:�È�È�=���(��#�a	����I  �n @H�i~�ab�ӋB�b�$w���"N0��  'Ж�q�p�@2��@���X�r�q5�C�pC0C�@ C���=�`
�A1q   @B�UV~X�
nwB0"h�A��p�ӊ�p�`���aDz���֏����Я	�pv�( �� -���I��-�=��A�a��we_q�`�p �?�ff ��m��>� ����ƼЇ!1!ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`�� <
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC��������#/*/c/N/�wi�����v/C�`� CHs/`
=$�p��<!�!��ܼ�'��3A�A�AR�1AO�^?�$��?���±�
=ç>�����3�W
=�#��]�;e�׬a@�����{�����<�>(��B�u���=B0�������	R��zH�F��G���G���H�U`E����C�+��}I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*O ONO9OrO]O�O�O�O �O�O�O�O_�O8_#_ \_G_�_�_}_�_�_�_ �_�_�_"oooXoCo |ogo�o�o�o�o�o�o �o	B-fQ� u������� ,��P�b�M���q��� ��Ώ���ݏ�(�� L�7�p�[������ʟ ���ٟ���6�!�Z��E�W���#1( �ٙ9�K���ĥ ������Ư!3��8���!4Mgqs��,�IB+8��J��a���{�d�d�����ȿ��쿔ڼ%P8�P�= :GϚ�S�6�h�z���R�Ϯ����������  %�� ��h� Vߌ�z߰�&�g�/9�$�������7�����A�S�e�w�   ������������̿2 F�$�&Gb��������!C���@���8������F� Dz�N�� F�P �D�������)#�B�'9K]o#?_���@@v
4$�8�8��8�.
 v��� !3EWi{�����:� ���ۨ�1��$M�SKCFMAP � ���� ���(.�ONREL  ��!9��EXC/FENBE'
#7%�^!FNCe/W$JO�GOVLIME'dtO S"d�KEYE'u�%�RUN�,��%�SFSP�DTY0g&P%9#S�IGNE/W$T1M�OT�/T!�_C�E_GRP 1p��#\x��?p� �?�?�?�?�?O�? OBO�?fOO[O�OSO �O�O�O�O�O_,_�O P__I_�_=_�_�_�_ �_�_oo�_:o��TCOM_CFG 1q	-�vo�o��o
Va_ARC_�b"�p)UAP_�CPL�ot$NOCHECK ?	+ �x�% 7I[m���������!�.+N�O_WAIT_L� 7%S2NT^ar�	+�s�_ERR�_12s	)9��  ,ȍޏ��x����&��dT_MO��t>��, ��*oq��9�PARAM��u	+��a�ß'g�{�� =?�345?678901�� ,��K�]�9�i�����`��ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDS�P�c#6p(OFFSET_CART�oη�DISƿ��PE?N_FILE尨!��ai��`OPTIO�N_IO�/��PW�ORK ve7s# ��V�ؤ!!p�p�4�p�	 ����p��<���RG_DSBL  ���P#��ϸ�RIE�NTTOD ?�Cᴭ !l�UT__SIM_D$�"����V��LCT w}�h�iĜa[�1ԟ_PEXE�j�R�ATvШ&p%� ��2�^3j)TEX)T�H�)�X d 3�������%�7�I� [�m��������������!�3�E���2 ��u���������������c�<d�AS ew������`��Ǎ�^0OUa0�o(��(�����u2, ����O H @D��  [?�aG?��cc�D][�Z��;�	ls��xJ��������<� ��� ���2�H(��H3�k7HSM5G��22G���Gpc
͜�'f�/,-,2�CR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t3�!�/ �/�"�t32����/6 W ��P%�Q%��%�|T��S62�q?�'e	'� � ��2I� � � ��+==�̡ͳ?�;	�h	�0��I  �n �@�2�.��Ov;���ٟ?&gN�]O  �''�uD@!� C�C��@F#H!�/�O�O Nsb
���@�@E��@�e`0B��QA�0Yv: �13Uwz$oV_�/z_�e_�_�_	��( �� -�2@�1�1ta�Ua�c����:Ar���.  �?�ff���[o"o�_!U�`oXÜQ8���o:�j>�1  Po�V(���eF0�f�Y����L�?����x�b�P<
6b<�߈;܍�<��ê<� <�#&�,/aA�;r��@Ov0P?fff?��0?&ip�T@�.�{r�J<?�`�u#	�Bdqt�Yc �a�Mw�Bo�� 7�"�[�F��j����� ��ُ����3�����,���(�E��� E��3G+� F��a��ҟ������,��P�;���B�pAZ�>��B��6�<O ίD���P��t�=����a�s�����6j�h�y�7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�<%?��?������(���#	Ę��P �N�||CH���Ŀx������@I�_��'�3A�A�A�R1AO�^??�$�?��� ��±
=ç>�����3�W
=�#� U��e����B��@��{�����<����(�B�u���=B0�������	�b�H��F�G���G���H�U`E����C�+��I�#�I��H�D�F��E��RC�j=[��
I��@H��!H�( E?<YD0߻� �������� �9�$� ]�H�Z���~������� ������#5 YD }h������ �
C.gR� ������	/� -//*/c/N/�/r/�/ �/�/�/�/?�/)?? M?8?q?\?�?�?�?�? �?�?�?O�?7O"O[O mOXO�O|O�O�O�O�O��O�O�O3_Q(���3���b��gUU���W_i_2�3ǭ8��_�_2�4M�gs�_�_�RIB+��_�_�a���{�miGo5okoYo(�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�u�,��  �p���o ��/��S��z
uү ܠ�������ڱ������������  /�M�w�e�������~�l2 F�$��'Gb��t��a�`�,p�S�C�y�@p�5��G�Y�۠F� D�z�� F�P D��]����پ��ʯܯ� ��~ÿ?���@@�J?�K�K���K���
 �|��� ����Ŀֿ������0�B�T�fϽ�V� ����{��1��$�PARAM_ME�NU ?3���  �DEFPULS�Er�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L��	�OPT���PTB4�.�C��R_DECSN ���e��ߑߣ����� ������!�3�\�W��i�{���USE_PROG %��q%�����CCR����e����_HOSoT !��!��:���T�`�V��/��X����_TIMqE��^��  ��?GDEBUG\�����GINP_FL'MSK����Tfp�����PGA  ��̹�)CH����TY+PE������� ����� - ?hcu���� ���//@/;/M/ _/�/�/�/�/�/�/�/��/??%?7?`?��W�ORD ?	=�	RSfu	P�NSUԜ2JO�K�DRTEy�]T�RACECTL �1x3��� }�`F G&�`��`�>�6DT Q�y3�%@�0D �  #T�Q2@�8B%6D&6DU'6D(6D)6D*6DT`8B,6D-6D.6D�/6D06D16A�c'�a8@U��BTR��H�D�D�C�2@M 8BJ�8BF�8B�6D6D	6D
6D�6D6D6D6D�6D^�8B6D6D�6D6D6D�8B*6D6D6D6DV�(8Bj�8B6D6DҀ(8B�8B!6D"6D5O GOYOkO}O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo�O�O�Oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՊ .AZev���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p ��Zer����� ,>Pbt� ������// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ����������� �*��$�PGTRACEL�EN  )�  ��(���>�_UP z/���m�u�Y��n�>�_CFG7 {m�W�(�En���PЬ� ���DEFSPD e|���aP��>��IN��TRL �}��(�8��IPE_CONFI��}~m��m����Ԛ�>�LID����=�GRP� 1��W���)�A ���&f�f(�A+33D��� D]� C�O� A@1��Ѭ(��d�Ԭ��0�0�� 	 1��1���G ´�����B� 9����O�9�s�(��>�T?�
5�������� =��=#�
���� P;t_��������  Dz (�
H�X ~i������ /�/D///h/S/�/���
V7.10�beta1��  A�E�"�ӻ�A (�� ?�!G��!>��r�"����!���!oBQ��!A\� P�!���!2p����Ț/8?J?\?n?};� ���/��/�?}/ �?�?OO:O%O7OpO [O�OO�O�O�O�O�O _�O6_!_Z_E_~_i_ �_�_�_�_�_�_'o 2o�_VoAoSo�owo�o �o�o�o�o�o.�R=v1�/�#F@ �y�}��{m��y =��1�'�O�a��? �?�?������ߏʏ� �'��K�6�H���l� ����ɟ���؟�#� �G�2�k�V���z��� �����o��ίC� .�g�R�d��������� �п	���-�?�*�c� ����Ϯ���� ��B�;�f�x����� ��DϹ��߶������ ��7�"�[�F�X��|� �����������!�3� �W�B�{�f������� �� �����/S >wbt���� ��=Ozό� �ψ����ϼ� / .�'/R�d�v߈߁/0 �/�/�/�/�/�/�/#? ?G?2?k?V?h?�?�? �?�?�?�?O�?1OCO .OgORO�OvO�O�O�� �O�O�O__?_*_c_ N_�_r_�_�_�_�_�_ o�_)oTfx�to ���/�o/ >/P/b/t/mo�| �������3� �W�B�{�f�x����� Տ�������A�S� >�w�b����O��џ�� ����+��O�:�s� ^�������ͯ���ܯ �@oRodo�o`��o�o �o��ƿ�o���*< N�Y��}�hϡό� �ϰ��������
�C� .�g�Rߋ�v߈��߬� ����	���-��Q�c� N�ﲟ���l����� ���;�&�_�J��� n�����������,� >�P�:L������� �����(�:�3 ��0iT�x�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?a?s? ��?�?X?�?�?�?�? O'OOKO6OoOZO�O ~O�O�O�O�O*\ &_8_r���_�_���$PLID_K�NOW_M  ~�� Q��TSV ��]�P��? o"o4o�OXoCoUo�o� R�SM_GRP� 1��Z'0{`J�@�`uf�e�`
�5� �gpk 'Pe]o�� ��������S+MR�c��mT�EyQ}? yR�������� ��폯���ӏ�G�!� �-������������ ����ϟ�C���)� ����������寧����QST�a1 1�j�)���P0� A 4��E2�D�V� h�������߿¿Կ� ��9��.�o�R�d�v�@���ϬϾ����2�90� Q�<3��A3�/�A�S��4l�~ߐߢ��5���������6
��.�@��A7Y�k�}���8���������MAD � )��P�ARNUM  �!�}o+��SCH
E� S�
��f���S��UPDf�x�|�_CMP_�`�H�� �'�UE�R_CHK-�a��ZE*<RSr��_�Q_MOG����_�X�_RES_G��!���D� >1bU�y�� ���/�	/����+/�k�H/g/ l/��Ї/�/�/�	� �/�/�/�X�?$?)? ���D?c?h?����?x�?�?�V 1��U��ax�@c]�@t�@(@c\�@��@D@c[�*@���THR_INR�r�J�b�Ud2FMA�SS?O ZSGMN�>OqCMON_QU?EUE ��U�V� P~P X�N$ U�hN�FV�@END8�A��IEXE�O�E���BE�@�O�COP�TIO�G��@PR�OGRAM %��J%�@�?���BT�ASK_IG�6^O?CFG ��Oz���_�PDATA�c�.�[@Ц2=�Do Vohozo�j2o�o�o�o �o�o);M j�INFO[��m� �D������ ��1�C�U�g�y��� ������ӏ���	�dwpt�l )�QE ?DIT ��_i�>�^WERFLX	C��RGADJ M�tZA�����?נ�ʕFA��IORIT�Y�GW���MPD�SPNQ����U�G�D��OTOE@1��X� (!A�F:@E� c�Ч!�tcpn���!�ud����!i�cm���?<�XY_��Q�X���Q)�� *�1�5��P��]�@�L���p��� �����ʿ��+�=Ϡ$�a�Hυϗ�*��P�ORT)QH��P��E��_CART�REPPX��SK�STA�H�
SSA�V�@�tZ	25?00H863���_�x�
�'��X�@�swPtS�ߕߧ���/URGE�@B��x	WF��DO�F"[�W\�������WRU�P_DELAY ��X���R_HO�TqX	B%�c���R_NORMALq^xR��v�SEMI�������9�QSKIP�'��tUr�x 	7�1�1��X�j�|� ?�tU������������ ��$J\n4 ������� �4FX|j� ������/0/ B//R/x/f/�/�/�/�tU�$RCVTM�$��D�� DCR�'���Ў!Cq��C�3�C����?�A!>��Q�<|�{:���p�� �����Š���Ҿ���|��:��o?�� <
6b�<߈;܍��>u.�?!<�&�?h?�?�? �@>��?O O2ODOVO hOzO�O�O�O�O�O�? �O�O__@_+_=_v_ Y_�_�_�?�_�_�_o o*o<oNo`oro�o�o �o�_�o�o�o�o�o 8J-n��_�� �����"�4�F� X�j�U������ď�� �ӏ���B�T�� x���������ҟ��� ��,�>�)�b�M��� ���������ïկ� Y�:�L�^�p������� ��ʿܿ� ����6� !�Z�E�~ϐ�{ϴϗ� ����-�� �2�D�V� h�zߌߞ߰������� ��
���.��R�=�v� ��k��������� �*�<�N�`�r����� �����������& J\?���� ����"4F�Xj|��!GN_�ATC 1�	;� AT&F�V0E0�A�TDP/6/9/�2/9�ATA��,AT%G1%B960�_+++�,��H/,�!IO_T?YPE  �%�#�t�REFPO�S1 1�V+ 'x�u/�n�/ j�/
=�/�/�/Q?<? u??�?4?�?X?�?�?^�+2 1�V+�/��?�?\O�?�O�?�!3 1�O*O<OvO�O��O_�OS4 1� �O�O�O_�_t_�_+_S5 1�B_T_f_�_o	oBo�_S6 1��_�_�_5o�o�o|�oUoS7 1�lo�~o�o�oH3l�oS8 1�%_����SMAS�K 1�V/  
8?�M��XNOS/�r�������!MOT�E  n��$��_CFG ����q����"PL_RANG������POWER� �����S�M_DRYPRG %o�%�P��TART ���^�UME_PRO�-�?����$_EXE�C_ENB  <���GSPD��Ր8ݘ��TDB��
�sRM�
�MT_'��T����OBO�T_NAME �o����OB_�ORD_NUM �?�b!H863  ��կ���PC�_TIMEOUT��� x�S232�Ă1�� L�TEACH PENDAN��w���-��Ma�intenanc?e Cons����s�"���KCLC/Cm��

���t��ҿ No U�se-��Ϝ�0�N�PO�򁋁z��.�CH_L��3����q	��s�?MAVAIL����糅��SPAC�E1 2��, j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��� ���ߚ� �2�D��� hߊ�|��`������ ����� �2�D�� h��|���`�������(��y���2���� 0�B���f�����{ ���3) ;M_����@��/� /44 FXj|*/���/��/�/?(??=?5 Q/c/u/�/�/G?�/�/ �?O�?$OEO,OZO6n?�?�?�?�?dO�? �?_,_�OA_b_I_w_7�O�O�O�O�O�_ �O_(oIoo^oofo�o8�_�_�_�_�_ �oo6oEf){�x��G �o�� ���
M� ���*�<�N�`� r�������w���o�収���d.��%� S�e�w����������� Ǐَ���Θ8�+�=� k�}�������ůׯ͟ ����%�'�X�K�]� ��������ӿ�������#�E�W� `� @�������x�����\�e����� ������R�d߂�8� j߬߾߈ߒߤ���� ������0�r���X� ������������8�����
�ύ�_M?ODE  �{��/S ��{|�2ς0�����3�	�S|)CWORK�_AD��t�L^+R  �{�`�� �� _INTV�AL���d���R_�OPTION� ���H VAT_�GRP 2��u;p(N�k|��_� ����/0/B/�� h�u/T� }/�/�/�/ �/�/�/?!?�/E?W? i?{?�?�?5?�?�?�? �?�?O/OAOOeOwO �O�O�O�OUO�O�O_ _�O=_O_a_s_5_�_ �_�_�_�_�_�_o'o 9o�_Iooo�o�oUo�o �o�o�o�o�o5G Yk-���u� ����1�C��g� y���M�����ӏ叧� 	��-�?�Q�c����� ����������ǟ��;�M�_����$SCAN_TIM���_%}�R ��(�#((�<0�4d d 
!D�ʣ���u�/�����U��25���@��d5�P�g��]	 ���������dd�x��  P����; ��  8� ҿx�!���D��$� M�_�qσϕϧϹ���������ƿv���F�X��/� ;G�ob��pm���t�_Di�Q̡  � l �|�̡ĥ������� !�3�E�W�i�{��� ������������/� A�S�e�]�Ӈ����� ��������); M_q����� ��r���j�T fx������ �//,/>/P/b/t/��/�/�/�/�/�%�/  0��6��!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O*�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo�O�OJ�o�o �o�o�o�o�o 2 DVhz��������
�7?   ;�>�P�b�t������� ��Ǐُ����!�3� E�W�i�{�������ß �ş3�ܟ�� &�8�J�\�n�������������ɯ�����,� �+�	�1234567�8�� 	� =5���f�x�������������
��.� @�R�d�vψϚ�៾� ��������*�<�N� `�r߄߳Ϩߺ����� ����&�8�J�\�n� �ߒ����������� �"�4�F�u�j�|��� ������������ 0_�Tfx��� ����I> Pbt����� ��!/(/:/L/^/ p/�/�/�/�/�/�/�2�/?�#/9?K?�]?�iCz  B}p˚   ��h�2��*�$SCR�_GRP 1�(��U8(�\x�d�@} � ��'�	 �3�1�2�4(1*�&��I3�F1OOXO}m��D�@�0ʛ�)���HUK�LM�-10iA 89�0?�90;��F;�M61C D�:�CTP��1
\&V�1 	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^�o OUO>oPo#G�/����o'o�o�o�o�oB��0�rtAA�0*  @�Bu&"Xw?��ju�bH0{�UzAF@ F�`�r��o���� �+��O�:�s��mBq�rr����������B� ͏b����7�"�[�F� X���|�����ٟğ�� �N���AO�0�B�CU�
L���E�jqBq>m3󵔯$G@�@pϯ7 B���G�I�
E�0EL_DEFAULT  �T���E���MIPOWERFL  
E*���7�WFDO� �*��1ERVENT? 1���`(��� L!DUM�_EIP��>��j�!AF_INEx�¿C�!FT�������!o:� ���a�!RP?C_MAINb�D�q�Pϭ�t�VIS}��Cɻ����!TP&��PU�ϫ�d��E��!
PMON_POROXYF߮�e4ߐ���_ߧ�f����!�RDM_SRV��߫�g��)�!R��Iﰴh�u�!
�v�M�ߨ�id���!RLSYNC���>�8���!R3OS��4��4��Y� (�}���J�\������� ������7��[" 4F�j|�����!�Eio�I�CE_KL ?%�� (%SVCPRG1n>����3��3���4�//�5./3/�6V/[/�7~/�/��D$�/�9�/�+�@� �/��#?��K?� �s?� /�?�H/�? �p/�?��/O��/ ;O��/cO�?�O� 9?�O�a?�O��?_ ��?+_��?S_�O {_�)O�_�QO�_� yO�_��Os��� �>o�o}1�o�o�o�o �o�o�o;M8 q\������ ���7�"�[�F�� j�������ُď��� !��E�0�W�{�f��� ��ß���ҟ��� A�,�e�P���t�����࿯�ί�y_DE�V ���MC:��_.!�OUT��2�~�REC 1�`e��j� �� 	 �����ȿ೿�׿��!�
 ��PJ�%6 (�޷&�!�a�}���u,��0�  Z�+ 3��3��Ge3�c���V��˒��� � ��$��H�6�l�~�`� �ߐ��ߴ������� � ��V�D�z�h��� ����������
�� R�@�v���j������� ������*N< ^�r����� �&J8Z� b������� "/4//X/F/|/j/�/ �/�/�/��2��/�/�/ ?:?(?^?L?�?�?v? �?�?�?�?�?�? O6O OFOlOZO�O~O�O�O �O�O�O_�O2_ _B_ h_V_�_n_�_�_�_�_ �_
o�_.o@o"odoRo tovo�o�o�o�o�o�o <*`Np� x������� 8�J�,�n�\������� ��Ə�Ώ�����F��4�j�X���`�p�V [1�}� P������ܺ.  K ����TYPE�\��HELL_CFG �.�F��Ϗ  	�����RSR������ӯ�� �����?�*�<�u� `�����������ο�  ��!%@�3�E��Q�\�Ӑ1M�o�p������2Ӑd]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&���!1�OW_REG�_UI��8�IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he���� ��������ж��) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������o���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( ��}3copy f�rs:order�fil.dat �virt:\tm�pback\=>�inspiron:3304��r��o�}*.mdb:*.*CU
Y����	.x.:\ �8R�n���/.a6HZ_� //�-?Qb/t/ �/�/�F/��/�/? ?)�M�/p?�?�? �8?J?��? OO�%�
xyzrate 61 �?�?�?nOȀO�O�%.GR(6368 HOZO�O�O_ "/4/�/�Ga_s_�_�_ �/E_�HY_�_�_o!? 3?FO�C�_no�o�o�? 6oHo�@^o�o&_ 8_�_�_m��_�_ �_Z���"o4o�o Xoi�{����o�oC��o ����O0Oԏe��w����O�O� 2112�OY�����!�3� ��˟ݟn���������400G�Y����� !3���a�s����� �E���Y�����!� 3�F�£ݿnπϒϥ� 6�H�Š^�����&� 8���ܿm�ߑߤ��� ȿZ������"�4��� X�i�{��ϲ�C��� ������0�B�T�e� w����߮�I������� ,��P�as� ���;��`� (����o��&�� ��deskto�p-mbmd4ji 208�Z�� /"4����o/�/x�/��4084N/ `/�/??(�:.�@�@�/�"h?z?�?�1���I?�+`?�?OO$���$SNPX_AS�G 1�����9A� P� 0 '%�R[1]@1.1,O �?�$�%dO�O sO�O�O�O�O�O�O _ _D_'_9_z_]_�_�_ �_�_�_�_
o�_o@o #odoGoYo�o}o�o�o �o�o�o�o*4` C�gy���� ���	�J�-�T��� c�������ڏ���� �4��)�j�M�t��� ��ğ������ݟ�0� �T�7�I���m����� ���ǯٯ���$�P� 3�t�W�i�������� ÿ����:��D�p� Sϔ�wω��ϭ��� � ��$���Z�=�dߐ� sߴߗߩ������� � �D�'�9�z�]��� �������
����@� #�d�G�Y���}����� ��������*4` C�gy���� ��	J-T� c������/ �4//)/j/M/t/�/ �/�/�/�/�/�/?0?�4,DPARAM ��9ECA W�	��:P�4�0�$HOFT_KB_CFG  q3�?E�4PIN_SI/M  9K�6�?��?�?�0,@RVQS�TP_DSB�>��21On8J0SR ���;� & M�ULTIROBO�TTASK=Oq3��6TOP_ON_ERR  �F��8�APTN z�5�@A�B�RING_PRM��O J0VDT_?GRP 1�Y9�@  	�7n8_(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2Dkh z������� 
�1�.�@�R�d�v��� ������Џ����� *�<�N�`�r������� ��̟ޟ���&�8� J�\�����������ȯ گ����"�I�F�X� j�|�������Ŀֿ� ���0�B�T�f�x� �ϜϮ���������� �,�>�P�b�tߛߘ� �߼���������(� :�a�^�p����� ������ �'�$�6�H� Z�l�~���������������3VPRG_CoOUNT�6��A��5ENB�OM�=�4J_UPD �1��;8  
 q2������  )$6Hql~ �����/�/  /I/D/V/h/�/�/�/ �/�/�/�/�/!??.? @?i?d?v?�?�?�?�? �?�?�?OOAO<ONO `O�O�O�O�O�O�O�O �O__&_8_a_\_n_��_�_�_YSDE�BUG" � �Pd�k	�PSP_PAS�S"B?�[LOoG ��m��P�X�_  ��g�Q
MC:\xd�_b_MPCm���o�o�Qa�o ��vfSAV �bm:dUb�U\g�SV�\TEM_T�IME 1��k (�`.�S,�o�	T1SVGUNYS} #'k�sp�ASK_OPTICON" �gosp�BCCFG ���| �b�{�}`����a&��#� \�G���k�����ȏ�� ����"��F�1�j� U���y���ğ���ӟ����0��T�f��U R���S���ƯA����� � ��D��nd��t9� l���������ڿȿ�� ���"�X�F�|�j� �ώ��ϲ�������� �B�0�f�T�v�xߊ� �ߦؑ�������(� ��L�:�\��p��� �������� �6�$� F�H�Z���~������� ������2 VD zh������ ���4Fdv� �����// */�N/</r/`/�/�/ �/�/�/�/�/??8? &?\?J?l?�?�?�?�? �?�?�?�?OO"OXO FO|O2�O�O�O�O�O fO_�O_B_0_f_x_ �_X_�_�_�_�_�_�_ oooPo>otobo�o �o�o�o�o�o�o :(^Lnp�� ���O��$�6�H� �l�Z�|�����Ə؏ ꏸ����2� �V�D� f�h�z�����ԟ�� ��
�,�R�@�v�d� ��������ίЯ�� �<��T�f������� &�̿��ܿ��&�8� J��n�\ϒπ϶Ϥ� ���������4�"�X� F�|�jߌ߲ߠ����� ������.�0�B�x� f��R���������� ��,��<�b�P����� ��x��������� &(:p^��� ���� 6$ ZH~l���� ����/&/D/V/h/ ��/z/�/�/�/�/�&�0�$TBCSG_GRP 2��%��  ��1 
 ?�  /?A?+?e?O?�? s?�?�?�?�?�;23��<d, ��$A?1	 HC�=��6>��@E�5?CL  B�'2^O�jH4J��B\})LFY  A�jOf�MB��?�IBl�O��O�@�JG_�@�  D	�15_ __$YAC-P{_F_`_j\��_�]@0�>�X�Uo�_ �_6oSoo0o~o�o�k��h�0	V3�.00'2	m6;1c�c	*�`�d�2�o�e>�JC0(��a�i ,p�m- ; �0����om�vu1JCFG -��% 1 #0vz+��rBrv�x����z� � %��I�4�m�X���|� �������֏���3� �W�B�g���x����� ՟��������S� >�w�b�����'2A �� ʯܯ������E�0� i�T���x���ÿտ� �����/��?�e�1 �/���/�ϜϮ����� ���,��P�>�`߆� tߪߘ��߼������ ��L�:�p�^��� ���������� �6� H�>/`�r�������� �������� 0V hz8����� �
.�R@v d������� //</*/L/r/`/�/ �/�/�/�/�/�/�/? 8?&?\?J?�?n?�?�? �?�?���?OO�?FO 4OVOXOjO�O�O�O�O �O�O__�OB_0_f_ T_v_�_�_�_z_�_�_ �_oo>o,oboPoro to�o�o�o�o�o�o (8^L�p� ������$�� H�6�l�~�(O����f� d��؏���2� �B� D�V�������n���� ԟ
���.�@�R�d�� ��v��������Я� ��*��N�<�^�`�r� ����̿���޿�� $�J�8�n�\ϒπ϶� ��������ߊ�(�:� L���|�jߌ߲ߠ��� �������0�B�T�� x�f���������� ����,��P�>�t�b� �������������� :(JL^�� ���� �6 $ZH~l��^� ��dߚ //D/2/ h/V/x/�/�/�/�/�/ �/�/?
?@?.?d?v? �?�?T?�?�?�?�?�? OO<O*O`ONO�OrO �O�O�O�O�O_�O&_ _6_8_J_�_n_�_�_ �_�_�_�_�_"ooFo ��po�o,oZo�o�o �o�o�o0Tf x�H����� ��,�>��b�P��� t���������Ώ�� (��L�:�p�^����� ��ʟ���ܟ� �"� $�6�l�Z���~����� دꯔo��&�ЯV� D�z�h�������Կ¿ ��
��.��R�@�v�8dϚτ�  ����� �������$�TBJOP_GR�P 2ǌ���  ?�������������xJ�BЌ��9� �<� �X����� @���	 ��C�� t�b  �C����>��1͘Րդ�>̚й���33=�C�Lj�fff?��?�ffBG��ь������t�ц�>��(�\)�ߖ�E����;��hCY�j��  @h��B�  A����f�~��C�  Dh�8��1��O�4�N�����
:���Bl^��j�i�l�l�����Aə�A��"��D��֊=qqH���нp�h���Q�;�A}�j�ٙ�@L��D	2�������$�6�>B�\��T���Q��tsx�@33@���C���y�x1����>��Dh�����������<{�h�@i�  ��t��	��� K&�j�n| ���p�/�/(:/k/�ԇ���!��	V3.00J��m61cI�*� IԿ��/�' �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I��!CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;��;Q�T,8�4` *�ϴ?�2���3\�X/O���ESTPARS c ��	���HR@ABLE 1���I�0��
H�7 8��9
G
H
H����*
G	
H

H
HYE���
H
H
HN6FRDIAO�XO@jO|O�O�O�ETO"_�4[>_P_b_t_�^:BS _� �JGoYoko}o �o�o�o�o�o�o�o 1CUgy�� ��`#oRL�y�_�_�_ �_�O�O�O�O�OX:B~�rNUM  �ū�P��� �V@P:B_CFG �˭�Z�h�@��IMEBF_TT%ApU��2@�VERS��q��R 1̞��
 (�/����b� ����J�\��� j�|���ǟ��ȟ֟� ����0�B�T���x��������2�_���@��
��MI_CH�AN�� � ��DOBGLV����������ETHERA�D ?��O��������h�����R�OUT�!��!�������SNMA�SKD��U�25�5.���#�����O�OLOFS_DI�%@�u.�ORQC?TRL ����� }ϛ3rϧϹ������� ��%�7�I�[�:����h�z߯�APE_D�ETAI"�G�PON_SVOFF=����P_MON ��֍�2��STRTCHK �^������VTCOM�PAT��O�����FPROG %^��%MULTIROBOTTݱ��֞9�PLAY&H��_�INST_Mް 2������US�q�΃�LCK���QUICKME�=���oSCREZ�G�tps� ���u�z����_��@@n��.�SR_GRP �1�^� �O����
��+O=sa�쀚�
 m������L/ C1gU�y� ����	/�-//�Q/?/a/�/	1234567�0�/�/�@Xt�1���
 ��}ipnl/�� gen.htm��? ?2?D?V?`�Panel s/etupZ<}P�?`�?�?�?�?�? �? ?,O>OPObOtO�O�? �O!O�O�O�O__(_ �O�O^_p_�_�_�_�_ /_]_S_ oo$o6oHo Zo�_~o�_�o�o�o�o �o�oso�o2DVh z�1'��� 
��.��R��v����������ЏG���UA�LRM��G ?9� �1�#�5�f� Y���}�������џן����,��P��SEoV  �����ECFG ���롽�A��  w BȽ�
 Q� ��^����	��-�?� Q�c�u������������� �����eI��?���(%D� 6� �$�]�Hρ�lϥ� ���ϴ�������#��G���� �߿U��I_Y�HIST �1��  (��� ��3/S�OFTPART/�GENLINK?�current=�editpage,��,1���!�3�ν�� ����me;nu��962�߆������K�]�o�36 u�
��.�@���W�i� {���������R����� /A��ew� ���N�� +=O�s��������f��f/ /'/9/K/]/`�/�/ �/�/�/�/j/�/?#? 5?G?Y?�/�/�?�?�? �?�?�?x?OO1OCO UOgO�?�O�O�O�O�O �OtO�O_-_?_Q_c_ u__�_�_�_�_�_�_ ��)o;oMo_oqo�o �_�o�o�o�o�o�o %7I[m�  �������3� E�W�i�{������Ï Տ�������A�S� e�w�����*���џ� ����ooO�a�s� ��������ͯ߯�� �'���K�]�o����� ����F�ۿ����#� 5�ĿY�k�}Ϗϡϳ� B���������1�C� ��g�yߋߝ߯���P� ����	��-�?�*�<� u����������� ��)�;�M������ ����������l� %7I[���� ���hz!3 EWi����� ��v////A/S/�e/P���$UI_�PANEDATA 1�����!�  	�}w/�/�/�/�/?? )?>?��/i? {?�?�?�?�?*?�?�? OOOAO(OeOLO�O �O�O�O�O�O�O�O_.&Y� b�>RQ? V_h_z_�_�_�__�_ G?�_
oo.o@oRodo �_�ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_ ��!�3�E�W��{� �_����ÏՏ���`� �/��S�:�w���p� ����џ������+� �O�a��������� ͯ߯�D����9�K� ]�o��������ɿ�� �Կ�#�
�G�.�k� }�dϡψ����Ͼ��� n���1�C�U�g�yߋ� �ϯ���4�����	�� -�?��c�J���� ������������;� M�4�q�X������� ����%7��[ �������@ ��3WiP �t�����/ �//A/����w/�/�/ �/�/�/$/�/h?+? =?O?a?s?�?�/�?�? �?�?�?O�?'OOKO ]ODO�OhO�O�O�O�O N/`/_#_5_G_Y_k_ �O�_�_?�_�_�_�_ oo�_Co*ogoyo`o �o�o�o�o�o�o�o�-Q8u�O�O}��������)�>��U-�j�|��� ����ď+��Ϗ�� �B�)�f�M������� �������ݟ�&�S��K�$UI_PA�NELINK 1��U  ��  ���}1234567890s��������� ͯդ�Rq����!�3� E�W��{�������ÿ�տm�m�&����Qo�  �0�B�T�f� x��v�&ϲ������� ��ߤ�0�B�T�f�x� ��"ߘ���������� �߲�>�P�b�t��� 0������������ $�L�^�p�����,�>�������� $�0,&�[gI�m� ������> P3t�i��� �� -n��'/9/K/ ]/o/�/t�/�/�/�/ �/�/?�/)?;?M?_? q?�?�UQ�=�2"� �?�?�?OO%O7O�� OOaOsO�O�O�O�OJO �O�O__'_9_�O]_ o_�_�_�_�_F_�_�_ �_o#o5oGo�_ko}o �o�o�o�oTo�o�o 1C�ogy�� ���B�	��-� �Q�c�F�����|��� ����֏�)��M� ��=�?��?/ȟڟ ����"�?F�X�j� |�����/�į֯��� ��0��?�?�?x��� ������ҿY���� ,�>�P�b��ϘϪ� ������o���(�:� L�^��ςߔߦ߸��� ����}��$�6�H�Z� l��ߐ��������� y�� �2�D�V�h�z� ���-���������
 ��.RdG�� }����c��� <��`r���� ����//&/8/J/ �n/�/�/�/�/�/7� I�[�	�"?4?F?X?j? |?��?�?�?�?�?�? �?O0OBOTOfOxO�O O�O�O�O�O�O_�O ,_>_P_b_t_�__�_ �_�_�_�_oo�_:o Lo^opo�o�o#o�o�o �o�o ��6H� l~a����� ���2��V�h�K� ������1�U
� �.�@�R�d�W/���� ����П������*� <�N�`�r��/�/?�� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��+������:� L�/�p���e������� ���� ��6����ۏ��$UI_�QUICKMEN�  ����}��REST�ORE 1٩��  �A
�8m3 \n���G�� ��/�4/F/X/j/ |/'�/�/�//�/�/ ??0?�/T?f?x?�? �?�?Q?�?�?�?OO �/'O9OKO�?�O�O�O �O�OqO�O__(_:_ �O^_p_�_�_�_QO[_ �_�_I_�_$o6oHoZo loo�o�o�o�o�o{o �o 2D�_Qc u�o������ �.�@�R�d�v����ଏ��Џ⏜SCR�E� ?��u1sc� u2��3�4�5�6��7�8��US#ER����T���Sks'���4��5���6��7��8��� N�DO_CFG mڱ  �  � PDATE h���None��SEUFRAM/E  ϖ���RTOL_ABRqT����ENB(�~�GRP 1��	��Cz  A� ~�|�%|�������įB֦��X�� UH��X�7�MSK  hK�S�7�N�%u�T�%�����VIS�CAND_MAX�I�I�3���FA?IL_IMGI�z ��% #S���IMR_EGNUMI�
����SIZI�� ��ϔ,�ONTM�OU'�K�Ε��&����a��a���s�FR�:\�� � �MC:\(�\L�OGh�B@Ԕ �!{��Ϡ�����z MCV�����UD1 �EX�	�z ��PO6�4_�Q��nm6��PO!�LI��Oڞ�e�V�N�fy@`�I�� =	_�wSZVmޘ��`��WAImߠ�STAOT �k�% @��4�F�T�$#�x ��2DWP  ���P G��=���͎���_J�MPERR 1��
  �p2345678901�� ��	�:�-�?�]�c� ��������������<��$�MLOW�ޘ������_TI/�˘'���MPHASE'  k�ԓ� ���SHIFT%�1 Ǚ��<z�� _����F /|Se���� ���0///?/x/ O/a/�/�/�/�/�/�����k�	VSF�T1\�	V��MN+3 �5�Ք p�����A�  B8*[0[0�Πpg3a1bY2�_3Y�7ME���K�͗	6e���&%���M���b���	��$��TDINGEND3�4��4OH�+�G1�OS2OIV �I���]LREL�EvI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�Y?BOX �ǝf_V\��b�2�TI�190.0.��P83p\�V2�54p^�Ԓ	 ��S�_�[b��?robot84q_   p�<9o\�pc�PZo Mh�]Hm�_Jk@1�o�ZABCd��k�, ���P\�Xo}�o0 );M�q���������>��aZ�b��_V