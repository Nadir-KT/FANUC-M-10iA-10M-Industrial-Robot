��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�   � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1���GPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|~GRG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"GSB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6*_�7_�8_�94F;CO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"YtP_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0��1p�34 >��DC �� Ќ@��hPV���mEX�p� �0g0xۤ�p�r
$TF��2C$MD3i�TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F�"F��?�@�a2 6�@$�PPU�3N�)ύRևA�X�!DU��AI�3BUF�F=�@1� |pp���pPIZT� PP�M��M�y��F�SIMQSI�"ܢVAڤrT�=�w T�`�(zM��P�B�qFAkCTb�@EW�`P1�BTv?�MC�� �$*1JB8`p�*1DEC��F�x�ŏ�� �H0�CHNS_EMP�1�$G��8��@_�4�3�p|@P��3�TCc�(r/�0-sx���ܐ� MBi��!����J�R� i�SEGFRR��Iv �aR�Tp9N�C��PVF4>�>bx &��f {uJc!�Ja��� !28�pץ�AJ���SIZ�3S�c�B�TM���g��>JaRSINFȑb� ��q�۽�н�����L�3�B���CRC�e�3CCp���� c��mcҞb�1J�cѿ��.����D$ICb�C q�5r�ե��@v�'���SEV���zF��_�եF,pN��ܫ�p?�4�0A�! �r ���h�Ϩ��p�2��@�a�� �د�R�Dx Ϗ��oH"27�!ARV�O`C�'$LG�pV�B�1�P��@�t�aA�0'�|�b+0Ro�� MEp`0"1 CRA 3 CAZV�g6p�O �#FCCb�`�`F�`K�8������ADI��a �A�bA'�.p��p�`�c�`S4PƑ�a�A�MP��-`Y�3P�M��s�UR��QUA1 � $@TITO1�/S@S�!����"0�D�BPXWO��B0!5�$SK���2ѓDBq�!"�"�PR�� 
� =���΁!# S q1$�2�$z���L�)$��/���� %�/�$Cr�!&?�$ENE�q�.'*?�Ú RE|�p2(H ���O�0#$L|3$�$�#�B[�;���FO�_D��ROS�r�#������3RIoGGER�6PApS|����ETURN�2n�cMR_8�TUw���0EWM���M�GN�P���BLA�H�<E���P��&$P� �'P@�Q3�CkD{��DQ���4��11��FGO_AWAY�BMO�ѱQ#!�� CS_�)  �PIS� I g�b {s�C��A��[  �B$�S��AbP�@�E9W-�TNTVճ�BV�Q[C�(c`�UWr��P�J��P�$0��SAsFE���V_SV�b�EXCLU��NnONL2��SY��*a&�OT�a'�HI�_V�4��B���_G *P0� 9�_z���p �TSG�� +nrr�@6A@cc*b��G�#@E�V.i|Hb?fANNUN$0,.$fdID�U�2�SC@�`�i�a��j�f���z��@I$2,O�c$FibW$}�OT9@��1 $DUM�MYT��da��dn��� � �E- ` ͑HE4(sg�*b�S|AB��SUFFIW�[�@CA=�c�5�g6�a��!MS�W�E. 8Q�KE3YI5���TM�10s�qA�vIN��#�p��D��/ D��H7OST_P!�rT���ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  A8	=ȳ�ј Tk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&Q�DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F��df�J� �q�aC1+�6 H�bLL_DUs�~a3@{��3:���OTX"���s�o��0NOAUTO�!7�p$)�$�*�R�c4�(�C� 8�IC, �"�!&�L�� 8H *8�LH <6����c"�` , `Ĭ�kª�q��q���sq��~q��7��8J��9��0����1��U1̺1ٺ1�1�U1 �1�1�2(ʩ2����2̺2ٺ2��2�2 �2�2*�3(�3��3��̺U3ٺ3�3�3 ��3�3�4(�3%����?��!9 < �9�&�z��I��1���M��QFE@'@� �: ,6��Q? �@P?9��5�9�E�@A�!�A�z� ;p$TP�?$VARI:�Z�n��UP2�P< ���TDe���K`Q�p���"���BAC�"G= T�p��e$)_,p�bn�kp+ IFIG� kp�H  ��P��"�F@`�!>t �;E��sC�ST �D� D���c�<�� 	C��{��_����l���R  ���FO�RCEUP?b��FWLUS�`H�N>�xF ���RD_CM�@E������ ��@vMP.��REMr F�Q��@1k@���7Q
K4	9NJ�5EFFۓ:f�@IN2Q��OVO�OVA�	TRO�V���DTՀ�DTMX� ��@�
�ے_PH"p��CL��_TpE�@�pK	_(�Y_T��v(���@A;QD� �������!0tܑ0R�Q���_�a����M̝7�CL�dρRIqV'�{��EARۑIOHPC�@����B�B��CM9@���R{ �GCLF��e!DYk(M�ap#5TuDG��� �%���FSSD �s? �P�a�!�1���P_(�!�(�!1��E�3�!�3�+5�&�GRA���7�@��;�PW泅ONn��EBU�G_SD2H�P{�_?E A �p�Z �TERM`59Bi5x�ORI#e0yCi5p�SM_�P�e0Di5�����TA�9E�6 ��UP\�F� -��A{�AdPw3S@B�$SEG�:� EL�{UUSE�@NFIJ�B$�;1젎4�4�C$UFlP=�!$,�|QR@��_G�90Tk�D�~SNST��PAT����AP'THJ3Q�E�p% B`�'EC���A�R$P�I�aSHFT�y�A�A�H_SHOQRР꣦6 �0$�7rPE��E�OVR=���aPI�@�U�b �QAYLOW����IE"�r�A��?���ERV��XQ�Y��mG�>@�BN��U\��Rz2!P.uASYMH��.uAWJ0G�ѡE q�A�Y�R�Ud>@ ��EC���EP;�uP�;�6WOR>@M`�]0SMT6�G3�cGR��13�aPAL@���`�q�uH � u���TOCA��`P	P�`$OP@����p�ѡ�`0YO��RE�`R4Cb�AO�p낎Be�`�R�Eu�h�A��e$7PWR�IMu�R�R_�cN��q=B �I&2H���p_AD�DR��H_LENAG�B�q�q�q$�R��S�JڢSS��SKN��u\��u̳�uٳ�SE�A�jrS��M-N�!K�����b����OLX��px����`ACRO3p J�@��X�+��Q��N6�OUP3�b_�IX��a�a1��}� ����(��H��D��`ٰ��氋�IO2S�D�����	�7�L $l��`Y!_�OFFr�PRM�_��"�HTTPu_+�H:�M (|p�OBJ]"�p��$���LE~Cd���N� � ��֑AB%_�TqᶔS�`6H�LVh�KR"u�HITCOU��B-G�LO�q����h�����`��`SS� ���HW�#A:��Oڠ<`INCP}U2VISIOW� ͑��n��to��to�ٲ� �IOLN��P� 8��R��p$�SLob PUTM_n�$p��P& x¢��Y F_AS�"Q��$L������DQ  U�0	P4A��50��ZPHY��-���x��UOI �#R `�K����$�u�"pPpk���$�������UJ5�S�-���NE6WJOG�KG̲DIS���K�p���#T (�uAV8F�+`�CTR�C
��FLAG2�LG�dU ���؜�13?LG_SIZ����`b�4�a��a�FDl�I`�w� m�_�{0a� ^��cg���4�����������{0��� SCH�_���a7�N�d�V
W���E�"����4�"�UM�Aљ`LJ�@�7DAUf�EAU�p��d|�r�GH�b�����BOO��WL ?�6 IT��y0��REC��SCR� ܓ�D
�\���MARGm�!��զ ���d%�����S����Wp���U� �JGM[��MNCHJ���FN�KEY\�K��PR�G��UF��7P��F�WD��HL��STP��V��=@��А�RS��HO`����C�9T��b ��7�[�U L���6�(RD� ����Gt��@PO������z��MD�FOCU���RGEX��TUI��I��4�@� L�����P����`���P��NE��CAN�A��Bj�VAIL�I�CL !�UDCS�_HII4��s�O��(!�S���S��1� ��BUFUF�!X�?PTH$m���v`�ě�*��AtrY�?P���j�3��`OS1Z2�Z3Z�1�� � Z � ��[aEȤ\��ȤIDX�dPSR�rO���zA�ST�L�R}�Y&�� /Y$E�C����K�&&�����![ LQ��+00�	P���`�#qdt
�U�dw<���_ \ �`4Г��\��Ѩ#\0C4�] =��CLDPL��UTRQLI��dڰ�)�$FLG&�� 1��#�D���'B�LD8�%�$�%ORGڰ5� 2�PVŇVY8�s�T�r�$}d^ ���$6��$�%S�`T� �B0��4�6RCLMC��4]?o?�9세�MI��p}d_ d=њR�Q��DSTB��p� ;F�HHA�X�R JHdLEXGCESr��BM!p
�a`�/B�T��B���`a�p=F_A@7Ji��KbOtH� K�d�b \Q���v$M�BC�LI|�)SREQUIR�R�a.\o��AXDEBUZ�AL
t M��c�b�{P����2�BNDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��XB� N&��aZ���UwPST� ezr7LOC�RIrp�EX<fA�p�9AA�ODAQ��f XfY�OND�rMF,� �Łf�s"��}%�e/�� ����FX3@IG}G�� g ��@t"��ܓs#N�s$R�a%��iL��hL�v<�@�DATA#?pAE�%�tR��Y�N�h t $MD
`qI}�)nv� ytq�ytHP`�Pxu��(�zsANSW)�yt@��
yuD+�)\b���0o��i �@CUw�V��p 0XeRR2��j� Du�{Q��7Bd$OCALIA@��G�:�2��RIN��"��<E�NTE��Ck��r^�آXb]���_N�qlk���9�D���B�m��DIVFDH�@���qnI$V�,��S�$��$AZ�X�o�*�����oH �$B�ELT�u!ACC�EL�.�~�=�ICRC�� ���D�T��8�$PS�@�"Ly�r��#^�S�E�<� T�PATH3���DI���3x�p�A_W ��ڐ���2nC��4��_MG�$DDx��T���$FW��Rp9��I�4��DE�7�PPABN��R?OTSPEE�[g�� J��[�C@4�~y$USE_+�2VPi��SYY��Z�1 qYN!@A��ǦOFF�qǡMO�U��NG���OL����INC�tMa6���HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]��BƉ�VE��#�y�23�_UP񕋳LOWL���p� B���Du�9B�``�x ���ByCv�r�MOSI���BMOU��@�7PE�RCH  ȳOV ��â
ǝ����D �ScF�@MP����� !Vݡ�@y�j�LUk��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A��x������N`�F�RTI�A$��MOUІ�HB@�BS0�p7D5����x��Z�DUM2ԓ�S_BCKLSH_Cx�k����ϣ����=���ޡ �	ACLAL"q��1м@N��CHK� �S�RTY��^�%E1rQq_�޴_UM�@r�C#��SCL0��r�LMT_J1_�L��9@H�qU�E�O�p�b�_�e�k�e�S�PC��u���N�P	C�N�Hz \P��C�0~"XT��C�N_:�N9��I�S	F!�?�V���U�/����x�T���CB!�SH�:��E�E1T�T�����y���T��PAL ��_P��_� �=������!����Jb6 L�@��OG��G�TORQU��ONֹ��E�R��H�E�&g_W2���_郅P���I�I�%I��Ff`xJ�1�,~1�VC3�0BD:B��1�@SBJ�RKF9�0DBOL_SM��2M�P�_DL2GRV�����fH_p��d���COS���LNH�� ������!*,�baZ���fMY��_(�TH��)TH�ET0��NK23����"��CB�&CB�CAA�B�"��!��!�&SB� 2�%'GTS�Ar�CIMa������,4#97#$DU���H\1� ��:Bk62�:AQ(rSf$NE�D�`I��B$+5��$̀�!A�%�5p�7���LPH�E�2���2SC%C�%�2-&FC0JM&̀V��8V�8߀LVJV�!KV/KV=KVKKV
YKVgIH�8FRM���#X!KH/KH=KH�KKHYKHgIO�<OR�8O�YNOJO!KUO/KO=KOKKOYKOM&F�2�!+i%0d��7SPBALANgCE_o![cLE0H_�%SPc� &�b�&�b&PFULC��h�b�g�b%p�1k�%�UTO_��Tg1T2�i/�2N�� "�{�t#�Ѱ`�0�*�.�T��OÀ<�v �INSEG"�ͱR�EV4vͰl�DIF��ŕ�1lzw��1m��0OBpq�я?�M�I{���nLCHW3ARY�_�AB��!�?$MECH�!o X��q�AX��P��p��7Ђ�`n 
��d(�U�ROB��C�Rr�H���-%��MSK_f`�p WP �`_��R/�k�z�����1S�~�|�`z�{���z��qINUq��MTCOM_�C� �q  ����pO�$NOR�En����pЂr� 8p GRe�uS�D�0AB�$XYZ_DA�1a���DEBUUq�������s z`$��COD��� L���p��$BUFIN�DX|�  <�M{ORm�t $ف�UA��֐����y��rG��u � $SIMUL  �S�*�Y�̑a�OBJ�E�`̖ADJUS<�ݐAY_IS��D�3����_FI�=��Tu 7�~� 6�'��p} =�C�}p�@:b�D��FRIr��MT��RO@ \�E}z���y�OPWOY�q�v0Y�SYS�BU/@v�$SOP�ġd���ϪUΫ}pPgRUN����PA���D���rɡL�_OUbo顢q�$)�/IMAG��w��0�P_qIM��L�IN�v�K�RGOVR!Dt��X�(�P*�J�|��0L_�`]��0�RB1�0��ML��ED}��p ��%N�PMֲ��c�w��SL�`q�w x �$OVSL4vS;DI��DEX�� ��#���-�V} *�N4�\#�B�2�G�B�_�M��y�q�>E� x Hw��p^��ATUSW����C�0o�s���BTMT�ǌ�I�k�4��x�԰q�y Dw�E&���@E�r��7�8�жЗ�EXE�����������f q�z �@w���UP'��$�pQ�XN�����x����� �PG΅�{ h $SUB����0_���!�_MPWAIv�P7�&��LOR�٠F\p˕�$RCVFAI�L_C��٠BWD�΁�v�DEFSP>!p | Lw����Я�\���UNI+�����H�R�+�}�_L\pP����P��p�}H�> �*�j��(�s`~�N�`KET�B�%�J�PE Ѓ~z��J0SIZE�����X�'���S�OR~��FORMAT�``��c ��WrEM�t��%�UX��G���PLI��p� � $ˀP_SWqI�pq�J_PL��?AL_ ����ХA��B��� C��Dn�$E��.��C_�U�� �� � ���*�J�3K0����TIA4��5��6��MOM���������ˀB��AD����������PU� NR�������G��m��� A$PI�6q��	 �����K4�)6��U��w`��SPEEDgPG������ ��Ի�4T�� �p @��SAMr`���\�]��MOV _�_$�npt5��5���1���2���������'�S�Hp�IN�'�@�+�����4($4+T+GAM�MWf�1'�$GE�T`�p���Da���
�
pLIBR>�II.2�$HI=�_g�t�$�2�&E;��(A�.� �&LW�-6<�)56��&]��v�p��V��$PDCK��D�q��_?����� q�&���7��4���9�+� �$IM_SR�pD�s�rF�L�r�rLE���Om0H]��0��-�pq���PJqUR_S�CRN�FA���S_?SAVE_D��dE@�NOa�CAA�b� d@�$q�Z�Iǡs	�I � �J�K� ����H� L��>�"hq��� ���ɢ�� bW^U�S�A�u��M4� ��a��)q`��3�WW� I@v�_�q�.MUAo��� � $PY�+�$W�P�vNG�{��P:��RA��RH��RO�PL�����qP� ��s'�X;�OI��&�Zxe ���m�� p��ˀ�3s�O�O��O�O�O�aa�_т� |��q�d@��.v��.v��d@��[wFv��E����%s�t;B�w�t|�tP���PMA��QUa ��Q�8��1٠QTH�H{OLW�QHYS��3ES��qUE�pZB���Oτ�  ��P�ܐ(�A����v�!�t�O`�q��u�"���8FA��IROG�����Q2���o�"��p�^�INFOҁ�׃hV����R�H�OI���� (�0SLEQ ������Y�3����Á��P0Ow0��5�!E0NU���AUT�A�COPAY�=�/�'��@Mg��N��=�}1������ ���RG��Á���X_�P�$;ख�`
��W��P��@��������EXT_CY�C bHᝡRpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�H�SdB����2�$��F�p���GPLeAdA
�TAR��Б@���P����裔d� ,�0F1L`�o@YN��K��M��Ck��PWR�+�9ᘐ��DELiA}�dY�pAD�a�� �QSKIPN4� �A�$�OB`�NT����P_ $�M�ƷF@\bIpݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q����TQ������ ���`���RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�d��REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"�������2�Қ�߼���P������3�қ'��9�K�]�o�� 
��4�Ҝ�������(�����5�ҝ!�3�@E�W�i�{�|@��6����������������7�ҟ-?Qcu�8�Ҡ��������SMSKJÁ�l��a��EkAޘ�MOTE6������@�݂TQ�IIO}5�ISTP���POW@��� ��pJ����p�����E�"$DSB_S�IGN�1UQ�x�C�\��S232����R�iDEVICE�US�XRSRPAR�IT��4!OPBI�T�QI�OWCONTR+�TQ��?SR�CU� MpSUXTASK�3N�p�0p$�TATU�PP�OG!�0�����p_�XPC)�$FRE?EFROMS	pna��GET�0��UPeD�A�2��SP� �:��� !$USAN�na&�����ERI�0�RpRIYq5*"_j@�Pm1��!�6WRK9KD����6��QFRIE3ND�Q�RUFg�҃��0TOOL�6MY��t$LENGT�H_VT\�FIR��pC�@ˀE> +IU�FIN-RM��R�GI�1ÐAITI��$GXñ3IvFG2v7G1���p3�B�GcPR�p�1F�O_n 0��!RE��p�53҅U�TC��3A�A�FG�G(��":���e1n!��J�8�%����%]��%�� 74��X O0�L��T�3H&��8���%b453%GE�W�0�WsR�TD����T��M����Q��T]�$V 2!����1�а91�8�0U2�;2k3�;3�: ifa�9-i�aQ��NSL��ZR$V��2BVwE�V�2A Q�B;�����&�S�`��F�"��k�@�2a�PS�E���$r1C��_3$Aܠ6wPR��7vMU�cS�t '�D$61�9�� 0G�aV`��p�d`���50�@���-�
25S�� E��aRW����B��&�N�AX�!�A�:@LAh��rTHI�C�1I���X�d1T�FEj��q�uIF_CH�3�qI܇7�Q�pG1RxV���]�岺:�u�_JF~�P�RԀƱ�RVAT��� ��`���0�RҦ�DOfE��CO9UԱ��AXI����OFFSE׆TRIGNS���c����h����H�Y��IGGMA0PA�pJ��E�ORG_UNE9V�J� �S����?�d �$CА�=J�GROU�����TOށ�!��DSP���JOGӐ�#��_	Pӱ�"O�q����@n�&KEP�IR��dܔ�@M}R��AP�Q�^�Eh0��K�SY�S�q"K�PG2�B�RK�B��߄�p`Y�=�d����`AD_�<����BSOC����N��DUMMY1�4�p@SV�PDE�_OP�#SFSP_D_OVR-���1C��ˢΓOR٧3�N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1q"�LCHDL��REGCOVʤc0��Wq@1M������RO�#��rȐ_+��� @0��e@VER�$O�FSe@CV/ �2WD�}��Z2����TR�!���E_�FDO�MB_CiM���B��BL�bܒ#��adtVQR�$0�p���G$�7�AM�5��� eŤ��_M�;��"'����8$C�A��'�E�8�8$HcBK(1���IO<�q����QPPA�ʀ����
��Ŋ����DVC_DBhC;�� #"<Ѝ�r!S�1[ڤ��S�3[֪�ATIO"q 1q� ʡU�3���CABŐ�2�CvP ��9P^�B���_� �?SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW�_C��U��S@��SA��A�pl$UNITm�l_�AT���e��ƐCYCLq�NE�CA���FLTR_2_FIO�7(�ӌ)&B�LPқ/�.�_�SCT�CF_`�F0b�l���|�FS(!E�e�CHA�1��4�D��"3�RSD��$"}�����_Tb�PR�O����� EMi_䙰a�8!�a �!�a��DIR0�R�AILACI�)RM�r�LO��C���Q`q��#q�դ�PR=�%S�A�pC/�� =	��FUNCq�0rRINP�Q�0��2f�!RAC �B ��p[���[WARn�F��BL�Aq�A����DAk�\���LD0���Q�d�qeq�TI"rp��K�hPRIA�!r"AF��Pz!=�;@��?,`�RK���Mǀ9I�!�DF_@B�l%1n�LM�FAq@OHRDY�4_�P@�RS�A�0� �MU�LSE@���aG ��ưt��m��$�1$�1$�1o����� x*�EG00�����!AR���Ӧ�09p�2,%� 7�AXE���ROB��WpA��_l-��SY[�W!‎&MS�'WRU�/-1��@�STR������Eb� 	�%��J��AB� ���&9�����kOTo0 	$��ARY�s#2��Ԓ��	ёFI@��$�LINK|�qC1��a_�#���%kqj2XYZ��t;rq�3��C1j2^8'0B��'�4����+ �3FI���7�q����'��_Jˑ���O3�Q'OP_�$;5���A#TBA�QBC��&��DUβ�&6��TURN߁"r�E11:�p��9GFL�`_���* Ȩ@�5�*7��Ʊ +1�� KŐM��&�8���"r��ORQ��a�(@#p=� j�g�#qXU�����mT'OVEtQ:�M��i�@��U��U��VW�Z �A�Wb��T{�, ��@ ;�uQ���P\�i��UuQ��We�e�SERʑe	��E� O���UdAas��4S�/7����AX��B� 'q��E1�e��i��i rp�jJ@�j�@�j�@�j P�j@ �j�!�f��i ��i��i��i��i �y�y�'y�7y�TqHyDEBU8�$32���qͲf2G + AB����رnS9VS�7� 
#�d� �L�#�L��1W��1W� JAW��AW��AW�QW��@!E@?D2�3LAB�29U4�Aӏ��Co s o�ERf�>5� � $�@_ mA��!�PO���à�0#�
�_MR}At�� d � 9T��ٔERR����;TY&���I��V8�0�cz�TOQ�d�PL[ �d�"�� ?�w��! � pp`T8)0���_V1Vr�a(Ӕ����2ٛ2�E�ĺ��@�H�E���$QW�����V!��$�P��o�cI��a�Σ	 HELL_�CFG!� }5��B_BASq��SR3��� �a#Sb���1�%���2��3��4��5*��6��7��8����RO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CYO. U�OUG�P~ �����m�������TPհ_KAR�l�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h��]��l0SEM�4�(�Ml4�6�TYN�SO���DIZ�~�A������m_TM�MAN�RQ��k0E�����$KEYSWIT�CH�ӵ�m���HE���BEAT��EF- LE~�����U���F!Ĳ���B�O_H�OM=OGREFUPPR&��y!� [��C��O��-ECO�C��Ԯ0_IOCMWD
�a���m���� � Dh1���U�X���M�βgPgCF�ORC��� ����OM.  � Q@�5(�U�#P, Q1��, 3��45���NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�� �� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E��VP���UPDs� � �`NЦ�5�YS�LOt�� � �L��d���A�aTAp�0d��|�ALU:eLd�~�CUѰjgF!a�ID_L�ÑeHI��jI��$FILE�_���d��$2�OveSA>�� hO�~�`E_BLCK���b$��hD_CPU yM�yA��c�o�db�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA�i�J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP�9_(�g�%�qr��� `�`GRO�Uw`��B��NF�LIC��f�REQ�UIRE3�EBU`��qB���w�2�����p���q5�p�� �\��APPR��C�}�Y�
ްEN٨CsLO7��S_M���H���u�
�qu�� ���MC�����N9�_MG��C�Co���`M�в�N�BRK�L�NOL|�N�[�R��_LINђ�|�=�	J����Pܔ������@�����������6ɵ��̲8k�+��q��ď� ��
��qx)��7�PATH3ǀL�B�L��H�wࡠ�6J�CN�CA�Ғ�lڢB�IN�rUCV��4a��C!�UM��Y,���aE�p�����ʴ���PAYLO�A��J2L`R_AN�q�Lpp����$�M�R_F2LgSHR��N�LO���Rׯ�`ׯ�ACRL_G�ŒЛ� ��9Hj`߂$HM��үFLEXܣ�qJ>�u� :�� �����������1�F1�V�j�@�R� d�v�������E���� ȏڏ����"�4�q� ��6�M���~��U�g�Hy�ယT��o�X�� H������藕?��� ��ǟِݕ�ԕ�����%�7��JJ�� � V�h�z���`cAT�採@�EL��S S��J|�Ŝ�;JEy�CTR��~��TN��FQ��HA_ND_VB-����v`�� $��F20M����ebSW��q�'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aDM)F�AW�Z`i�Aw�AA��X X�'pi�Dw��D��Pf�G�p�)S�Tk��!x��!N��DY�pנM�9$`%Ц� H��H�c�׎���0� ��Pѵڵ������������� ����1��R�6��QA'SYMvř���v���J���cі�_SH >��ǺĤ�ED����������J�İ%��C��IDِ�_VI��!X�2PV_UNIX�FThP�J��_R�5 _Rc�cTz�pT�V��@�@��İ�߷��U �Ԓ��	D���Hqpˢ���aEN�3�D	I����O4d�`J��� x g"IJAA �az�aabp�coc�`a��pdq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a��iT�@<� $�DUMMY9Q�o$PS_��RFC�v�$v �p8���Pa� XƠ����STE���SB}RY�M21_VF�8$SV_ERF�qO��LsdsCLRJtEA��Odb`O�p� � D $�GLOBj�_LO ���u�q�cAp�r�@awSYS�qADR`�`�`TCH  �� ,��ɩb�W_NA���7���SR���l ���
*?�&Q�0" ?�;'?�I)?�Y)��X� ��h���x������)�� Ռ�Ӷ�;��Ív�?���O�O�O�D�XSCSRE栘p����3ST��s}y`��R��/_HA�q�� TơgpTYP �b���G�aG�蕵�Od0IS_�䓀daUEMd� �����ppS�qaR�SM_�q*eUNE�XCEP)fW�`S_}pM�x���g�z�����ӑCOU��S�Ԕo 1�!�UE&���Ubwr��PROG�M�FL@$C�UgpPO�Q���U�I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp��OUS�� �� @6p�v$BU�TTp�RpR�CO�LUMq�e��SE�RV5�PANE|H�q� � �@'GEU���Fy��?)$HELPõ)B/ETERv�)ෆ� ��A � ��0`��0��0ҰIN簊�c�@N��IH�1��_� �v��LN�r� �qprձ_ò=�$H���TEXl����F�LA@��RELVB��D`��������M��?,�ű�m�����"�USRVwIEW�q� <6p�`U�`�NFI<@;�FOCU��;�7PRI� m�`�Q�Y�TRIP�qm��UN<`Md� x#@p�*eWARN)e��SRTOL%���g��ᴰONCOR�N��RAU����T����w�VIN�Le�� $גPA�TH9�גCACH���LOG�!�LI�MKR����v���HwOST�!�bz�R��OBOT��d�IM>� �� ����Zq�Zq;�V�CPU_AVAIYL�!�EX	�!AN���q��1r��1r���1 �ѡ�p� � #`C����@$�TOOL�$��_wJMP� ���e$SS���g ?�VSHIF��Nc�P�`ג�E�ȐyR����OSUR��=Wk`RADILѮ��_�a��:�9a��`a��r��LULQ$O�UTPUT_BM����IM�AB �@��rTILSC	O��C7��� ����&��3��A����q���m�I�2JG�АV�pLe�}���yDJU��N�/WAIT֖�}���{�%! NE�u�Y�BO�� ��� $`�t�SB�@TPE��NEC�p�J^FY�nB_T��R�І�a$�[$YĭcB��dM���F� m�CH$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"�`�"��[���P?� ]АZAB�C%��  $��"R��
�  ��$$CLAS������!ϐ� � � VIRT]��/ 0gABS����1 5�� < �!F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6HpZi{0-�AXL�pt��"�63  �{t�IN��qztPRE������v�p�uLA�RMRECOV c9�rwtNG��� .;	 A �  �.�0PPL�IC��?5�p��Hand�lingTool� o� 
V7.�50P/23-� � �Pz��
���_SWt� UPn�!� x�F0���t�QzA� v�� 864�� �it�y�2��2 7D�A5�� �� �d��@ϐo�Non�eisͅ˰ ���T���!�A�yx>�_l�V��uT��s9�UTO��"�Њt�y��HGA�PON
0g�1��U�h�D 1581����̟ޟry��^��Q 1��� �p�,�蘦���;�p@��q_��"�"� �c�.�H����D�HTTHKYX��"�-�?�Q� ��ɯۯ5����#�A� G�Y�k�}�������ſ ׿1�����=�C�U� g�yϋϝϯ�����-� ��	��9�?�Q�c�u� �ߙ߽߫���)���� �5�;�M�_�q��� �����%�����1� 7�I�[�m�������� ��!����-3E Wi{���� ��)/ASe w����/�� /%/+/=/O/a/s/�/ �/�/�/?�/�/?!? '?9?K?]?o?�?�?�? �?O�?�?�?O#O]����TO�E�W�DO?_CLEAN��7���CNM  � �__/_A_S_��DSPDRYRL�O��HIc��M@�O �_�_�_�_oo+o=o Ooaoso�o�o���pB�F�v �u���aX�t�������9�PLUG�G���G��U�PRC*vPB�@��_�o�rOr_7�SEGF}�K[mwxq�O�O������?rqLAP�_�~q�[�m�� ������Ǐُ�����!�3�x�TOTAL��f yx�USENU
�p�� �H���B���RG_STRIN�G 1u�
��Mn�S5�
~ȑ_ITEM1Җ  n5�� ��$� 6�H�Z�l�~������� Ưد���� �2�D��I/O SI�GNAL̕T�ryout Mo{deӕInp���Simulate�dבOut���OVERR�P �= 100֒I?n cycl��ב�Prog Ab�or��ב��St�atusՓ	Heartbeatї�MH Faul<��Aler'�W� E�W�i�{ύϟϱ������� �CΛ�A ����8�J�\�n߀ߒ� �߶����������"��4�F�X�j�|���WOR{pΛ��(ߎ�����  ��$�6�H�Z�l�~� �������������� 2PƠ�X  ��A{����� ��/ASe�w�����SDEV[�o�#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U?|g?y?PALT� �1��z?�?�?�?�?O "O4OFOXOjO|O�O�O��O�O�O�O�O_�?GRI�`ΛDQ�?_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o�o�o2_l�R��a\_ �o"4FXj| ����������0�B�T��oPREG�>�� f���Ə؏ ���� �2�D�V�h� z�������ԟ���~Z��$ARG_���D ?	����;�� � 	$Z�	[O�]O��Z�p�.��SBN_CONF�IG ;��������CII_S�AVE  Z������.�TCELL�SETUP �;�%HOME_�IOZ�Z�%MO�V_��
�REP��lU�(�UTOBA�CKܠ���FRA:\z�c \�z�Ǡ'`�qz���n�INI�0�z���n�MESSAG���ǡC�>��ODE_D����ą�%�O�4�n�PA�USX!�;� ((O>��Ϟˈ� �Ϭ���������� *�`�N߄�rߨ߶�g�~l TSK  w�xԿ׿q�UPDT+���d!�A�WSM�_CF��;����'�-�GRP 2�:�?� N�BŰA|��%�XSCRD1�;1
7� �ĥĢ����������*� ������r��������� ��7���[�&8J�\n��*�t�GR�OUN�UϩUP�_NA�:�	�t��_ED�1�7�
 �%-B?CKEDT-�2��'K�`���-(t�z�q�q�z���2t1�����q�k�(/��ED3/��/�.pa/�/;/M/ED4�/ t/)?�/.?p?�/�/ED5`??�?<?.p�?O�?�?ED6O �?qO�?.MO�O'O9OED7�O`O_�O.p�O\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o��_	-9o�oo%oCR_ 9]�oF�o�k� � NO_D�EL��GE_U�NUSE��LA�L_OUT �����WD_AB�ORﰨ~��pIT_R_RTN��|ONONSk����˥CAM_PAR�AM 1;�!�
� 8
SONY� XC-56 2�34567890� ਡ@����?��( С�\�
���{����^�HR5q�̹��ŏ�R57ڏ�Af�f��KOWA �SC310M
��x�̆�d @ <�
���e�^��П \����*�<��`��r�g�CE_RIA�_I�!�=�Ff��}�z� ���_LIU�]������<��FB�GP� 1��Ǯ��M�_�q�0�C* Y ����C1��9���@��G���CR�CU]��d��l��s��QR�����[Դm���v���������W C����(���숁=�HE�`ONF�Iǰ�B�G_PR/I 1�{V�� �ߖϨϺ�����������CHKPAUS��� 1K� , !uD�V�@�z�dߞ߈� ���߾������.��R�<�b���O���������_MOR��� �6��� 	 �����*�� N�<�������?Ғ�q?;�;����K���9�P���ça�-:���	�

��M���pU�ðț�<��,~��DB��튒)
mc�:cpmidbg��f�:�  &Ӱ^¥�p�/��  �(�Z(��� �s>܌���+�W��?�>��XgX�/�w�pxU�f�M/w�O/�
DE�F l��s)��< buf.txAts/�t/��ާ��)�	`�����=L����*MC��1�����?43��1���t�īCz  �BHH�B��_C�A��}2���BE��Y
�K�D6��CФ�B�s���D��9�D
}ʥ=F�6�*E��D�S����Fǔ_F7bY	���'w�K1���s���U.�p������BD�w�M@,!J�C�2�����g@D��0�0�EYK�EX��EQ�EJP �F�E�F� �G��>^F �E�� FB� �H,- Ge���H3Y��:���?33 ���~�  n8�~@��5�Y�E>�ðA��Y<7#�
"Q ����+_�'RSMOFSb�p�.8��)T1���DE ��F 
Q��;�(PB_<_��R����	op6�C4P�;s@ ,!(Q�2s@C�0B3�Ma�C{@@�3w��UT��pFPROG !%�z�o�oigI�q����v��ldKEY_TOBL  �&S�#�� �	
��� !"#$%&'�()*+,-./�01i�:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�����������������������p`LCK�l4�p`�`STAT� ��S_AUTO_�DO���5�IN?DT_ENB!���1R�Q?�1�T2}�^��STOPb���TR�Lr`LETE���Ċ_SCREEN� �Zkc�sc��U��MME�NU 1 �Y  <�l�oR�Y 1�[���v�m���̟�� ���ٟ�8��!�G� ��W�i��������ï կ��4���j�A�S� ��w�����迿�ѿ� ���T�+�=�cϜ�s� ���ϩϻ������� P�'�9߆�]�o߼ߓ� ���������:��#� p�G�Y������� ����$����3�l�C� U���y������������ ��	VY)�_M�ANUAL��t�DwBCO[�RIGڇ>
�DBNUM� ����1d e
�PXW�ORK 1!�[ �_U/4FX�__AWAY�i�/GCP  b=�Pj�_AL� #�j�Yи�܅ `�_�  1}"�[ , 
�@mg�&/~&lMZ��IdPx@P@#ON�TIMه� dɼ`&�
�e�MO�TNEND�o�R�ECORD 1(��[g2�/{�O� �!�/ky"?4?F?X? �(`?�?�/�??�?�? �?�?�?)O�?MO�?qO �O�O�OBO�O:O�O^O _%_7_I_�Om_�O�_  _�_�_�_�_Z_o~_ 3o�_Woio{o�o�_�o  o�oDo�o/�o S�oL�o���� @���+�yV,� c�u��������Ϗ>� P�����;�&���q� ��򏧟��P�ȟ�^� �����I�[�����  ���$�6��������jTOLEREN�CwB���L��͖ CS_CFG� )�/'d�MC:\U�L%0?4d.CSV�� �c��/#A ��CH
��z� //.ɿ���(S�RC_OUT *��1/V�?SGN +��"���#�17-F�EB-20 19�:090j�( PQ�8�ɞ�/.���f�pa�m�?�PJPѲ���VERSION �Y�V2.�0.84,EFLO�GIC 1,� 	:ޠ=�ޠ�L��PROG_E�NB��"p�ULS�k' ����_WRSTJNK ��"f�EMO_OPT_�SL ?	�#
� 	R575 /#=�����0�B��>��TO  �ݵ�l���V_F EX��d�%��PATHw AY�A\�����5+ICT�F�u-�j�#�egS�,�ST?BF_TTS�(�	�d���l#!w�� M�AU��z�^"MSWX�.�<�4,#�Y�/�
!J�6%�ZI~m��$SB�L_FAUL(�0��9'TDIA[�1�<�<� ����12345678#90
��P��H Zl~����� ��/ /2/D/V/h/��� P� ѩ �yƽ/��6�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�,/�gUMP���� ��ATR���1OC@P�MEl�OOY_TE{MP?�È�3F�8��G�|DUNI��.��YN_BRK �2_�/�EMGDI�_STA��]��EN�C2_SCR 3�K7(_:_L_^_ l&_�_�_�_�_)��C�A14_�/oo/o�AoԢ�B�T5�K�ϋo~ol�{_�o�o �o'9K]o �������� �#�5��/V�h�z��� �`~�����ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T���x������� ��ү�����,�>� P�b�t���������ο ����(�f�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ���������:�  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� �����*<N `r������ �&8J\n ���������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?��? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O��O�O__NoETM�ODE 16�5]�Q �d�X�
X_j_|Q�PRRO�R_PROG �%GZ%�@��_  ��UTABLE  G[�?oo)oRj�RRSEV_NU�M  �`WP��QQY`�Q_AU�TO_ENB  q�eOS�T_NOna� 7G[�QXb�  *��`��`��`��`d`+�`�o�o�o�dHISUc�aOP��k_ALM 18.G[ �A��l�P+�ok}������o_Nb�`  �G[�a�R
�:PTC�P_VER !�GZ!�_�$EXTLOG_REQvs�i\�SIZe�~W�TOL  �a{Dzr�A W�_BWD�p��xf́�t�_DI�� 9�5�d�T�asRֆSTEP��:P�_OP_DOv�f��PFACTORY�_TUNwdM�E�ATURE :��5̀rQH�andlingT�ool �� \s�fmEngl�ish Dict�ionary��r�oduAA �Vis�� Mas�ter����
E�N̐nalog �I/O����g.f�d̐uto So�ftware U�pdate  F� OR�mati�c Backup~��H596,��ground E�ditޒ  1 �H5Came�ra�F��OPL�GX�ell𜩐IwI) X�ommՐsshw���com��sco���\tp����pane��  �opl��tyle select��/al C��nJ�Ց�onitor��R�DE��tr��R�eliab𠧒6�U�Diagnosx(�푥�5528��u��heck S�afety UI�F��Enhanc�ed Rob S�erv%�q ) �"S�r�User �Fr[�����a��xt. DIO ��fiG� sŢ��e�ndx�Err�L&F� pȐĳr됮�� ����  !��F�CTN Menu�`�v-�ݡ���TPw Inېfac��  ER J�GC�pבk Ex�ct�g��H558���igh-Spe�x�Ski1�  2�
P��?���mm�unic'�ons��&�l�ur�ې���ST Ǡ��co�nn��2��TXP�L��ncr�st�ru����"FAT�KAREL �Cmd. LE�u�aG�545\��R�un-Ti��En=v��d
!����ؠ++�s)�S/W���[�LicegnseZ��� 4T��0�ogBook(�Syڐm)��H5�4O�MACROs�,\�/Offsen��Loa�MH��ܽ���r, k�Me�chStop P�rot���� li�c/�MiвShiqf����ɒMixx���)���,e�S�M�ode Swit�ch�� R5W�M�o�:�.�� 74� ���g��K�2~h�ulti-T=��M���LN (�Pos�Regi�ڑ������d�ݐt 'Fun�ǩ�.�����Num~����� �lne��ᝰ A�djup����� � - W��tat�uw᧒T�R�DMz�ot��scWove U�9����3Ѓ�uest' 492�*�o������62;�SNPX� b ���8 J7<`���Libr��J�#48���ӗ� �Ԅ��
�6O�� Par�ts in VCCMt�32���	��{Ѥ�J990��/�I� 2 P��T_MILIB��H�:��P�AccD�L�o
TE$TX��n��ap1S�Te����pkey��w����d��Une�xceptx�mo�tnZ��������є�� O����� 90J�єSP CSXC<�f���6�� Py�We}���gPRI�>vrЮt�men�� ��iPɰa������vGrid�pl�ay��v��0�)�H�1�M-10iA�(B201 �2�\� 0\k/�Ascii�l�Т�ɐ�/�Col��ԑGu�ar� 
�� /Pl-�ޠ"K��st{�Pat ��!S�C�yc�҂�ori�e��IF8�ata- quҐ�� ƶ���mH574��RL���am���Pb�H_MI De3�(b�����PCϺ�Pa�sswo+!��"P�E? Sp$�[���t�p��� ven��T�w�N�p�YELL�OW BOE	k$A;rc��vis��y3*�n0WeldW��cial�7�V#t&�Op����1y�� 2F�a�por1tN�(�p�T1�T�0 �� ��xy]�&kTX��tw�igjx�1� b� ct\��JPN ARCPSU PR��oݲ�OL� Sup�2f�il� &PAɰאc{ro�� "PM(�X���O$SS� eв7tex�� r���z=�t�ssagT��P��P@�Ȱ�����rtW��H'>�r�dpn��n1�
t�!� z ��a�scbin4ps�yn��+Aj�M �HEL�NCL �VIS PKGS� PLOA`�MB� �,�4VW�R�IPE GET_�VAR FIE �3\t��FL[�O�OL: ADD �R729.FD �\j8'�CsQ�QE���DVvQ�sQNO? WTWTE��}PD  Dp��biR�FOR ��ECT�n�`��ALSE �ALAfPCPMO�-130  M"� #h�D: HANG FROMmP��AQfr��R70�9 DRAM A�VAILCHEC�KSO!��sQVPC�S SU�@LIM�CHK Q +P~dF_F POS��F�Q� R5938�-12 CHAR�Y�0�PROGRAy W�SAVEN`wAME�P.SV��7��$En*��p?F�U�{�TRC|� S�HADV0UPDA�T KCJўRST�ATI�`�P MU�CH y�1��IM�Q MOTN-0�03��}�ROBO�GUIDE DA�UGH�a���*�t�ou����I� Šh�d�ATH�PepMO�VET�ǔVMX�PACK MAY ASSERT�Dn��YCLfqTA�r�BE COR v�r*Q3rAN�pRC� OPTIONS�J1vr̐PSH-�171Z@x�tcǠSU1�1Hp^9R!�Q��`_T�P��'�j��d{tby ap?p wa 5I�~d��PHI���p�aTE�L�MXSPD �TB5bLu 1��UBl6@�qENJ`CE2��61��p��s	�m�ay n�0� R�6{�R� �Rtrasff)�� 40*��p��fr��sys�var scr �J7��cj`DJUD��bH V��Q/�PSET ERR`�J` 68��PND�ANT SCRE�EN UNREAh��'�J`D�pPA��z�pR`IO 1����PFI�pB�pGROUN�PD��G��R��P�QnRSVIP �!p�a�PDIGIT� VERS�r}BL�o�UEWϕ P0�6  �!��MAG`p�abZV�DI<�`� SSUE�ܰ��EPLAN J=OT` DEL�pݡ�#Z�@D͐CAL9LOb�Q ph��RޫQIPND��IM�G�R719��MwNT/�PES �puVL�c��Hol�08Cq���tPG:�`C��M�canΠ��p�g.v�S: 3D� mK�view ed�` �p��ea7�:��b� of �Py����ANNOT ACCESS M��tƁ*�t4s a���lok��Flexj/:�Rw!mo?�PA?�-�����`n�pa SNBPJ? AUTO-�06f�����TB��PIAB{LE1q 636���PLN: RG$�pul;pNWFMDB��VI���tWIT �9x�0@o��Qui�#0�ҺPN RRS�?pUSB�� t & remov�@� )�_��&AxEPF�T_=� 7<`�pP�:�OS-144 ��h s�g��@�OST� � CR�ASH DU 9^��$P�pW� �.$��LOGIN���8&�J��6b04�6 issue �6 Jg��: Solow �st��?c (Hos`�c����`IL`IMPR�WtSPOT:Wh�:0�T�STYW ./�VMGR�h�T0wCAT��hos���E�q��� �O:�S:+pRTU' k�e-S� ����E:���pv@�2�� t\h�ߐ��m ��alļ�0�  $�H� W�A͐��3 CNT�0 T�� Wro>U�alarm���0s�d � �0SE1���t�r R{�OMEBp����K� 55��R�EàSEst��g �    �KA7NJI�no����INISITALcIZ-p�dn1weρl<��dr�� lx`~�SCII L�fails w��y ��`�YSTEa�p��o��Pv� IIH����1W�Gro>Pmo ol\wpSh@��P��Ϡn cfl�xL@АWRI �OGF Lq��p?�F��up��de-re�la�d "AP�o SY�ch�Abe�twe:0IND 1t0$gbDO����r� `�GigE��#operabi-lf  PAbHi�H`���c�lead�\�etf�Ps�r�O�S 030�&: fi=g��GLA )P ���i��7Np tpkswx�B��If�Ag������5aE�a EXCE#dU�_��tPCLOS��"r[ob�NTdpFa�U�c�!���PNI�O V750�Q1p��Qa��DB ��b�P M�+P�QED��DET��-� \r�k��ONLINEhSBUGIQ ߔĠ,i`Z�IB�S ap�ABC JARK�YFq� ���0MI�L�`� R�pNД \�p0GAR��D*pqR��P�"! jK�0cT�P�Hl#n�a��ZE V�� TA;SK�$VP2(�4`�
�!�$�P�`WIB�PK05�!FȐB�/��BUSY R7UNN�� "��d���R-p�LO��N�DIVY�CUL���fsfoaBW�p���30	V���ˠIT`�a50�5.�@OF�UN#EX�P1b�af�@�}E��SVEMG� �NMLq� D0pC?C_SAFEX 0c��08"qD �PETr�`N@�#J87��B��RsP�A'�M��K�`K�H GU�NCHG۔MEC�H�pMc� T�  �y, g@�$ OR?Y LEAKA�;�ޢSPEm�Ja��V�tGRIܱ�@އCTLN�TRpk�FpepR�j50�EN-`IN�����p� �`�Ǒk!��T3�/dqo�STO�0A�#�L�p �0�@�Q��АY�&�;pb1T!O8pP�s���FB�@�Yp`�`DU��aO��supk�t4 � P�F�� Bnf�Q�PSV�GN-1��V�SRSR)J�UP�a2�Q�#D�q l O���QBRKCTR 5Ұ�|"-�r�<pc��j!INVP�D ZO� ��T`h#�Q�cH�set,|D��"D�UAL� w�2*BRVO117 A]��TNѫt�+bTa24A73��q.?��r�{1} 009.fd8��y`j604.\P-^�`hanc�U�� F��e8��  ��npJtPd!q��`��w� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� \P��R�R(}\\Pe� aʰ�I���E��1��p�� j  �� ,e�Dp� �A�A\P�q �5 sig��a��"AC;a��
�bCe�\Pb_p��.pc�]l<bHbcb_cicrc~h<n�`tl1� ~`\P`o�d\P�b]o2�� �cb�c�i\P�jupfrm�d\P�o�`exe�a�oFd\Ptped}o��u`�cptlibxz\P�l�cr�xr\P\�blpsazEd\P_fm�} gc\P�x���o|sp�or�mc(��ob_jzo"p�u6�wf��t���wms�1q��sld�)��jmc�o\�n�b�nuhЕ��|st�e���>�pl�qp�iwc1k���uvf0uߒ<��lvisn�CgoaculwQ
E �`RFciV\PqiP��D�ata Acqu�isi��nZU�SR�631`��TR�QD�MCM �2�P7u5H�1�P583\Pm1��71��59`�5�P57<P\P�Q�����(���Q��o yp\P!daq\�1oA��@�� ge/��etdms�"DM�ER"؟,�pgdD���.�m���-��q�aq.<᡾\Pmoȷ�h���f{�oR50�3��MACROso, Sksaff�@(lR���03�SR�Q(�*�Q6��1�Q9ӡ�R�ZSh��P\PJ643�@7ؠ6�P�@�PRS�@���e �Q�U�С PIK�Q52 PTLC�W��\Pw3 (��p/O� �!�Pn �\P5���03\sfmnmc "MNMCq�<��Q��\$AcX�FM���ci,Ҥ�X���`�cdpq+�
�sk��SK�\P�SH56�0,P��,�y�refp "REFp�dd�A�j\P	�of�cOFc�<gy�to��TO_����ٺ����+je�u��ca�xis2�\PE�\�e>�q"ISDTc���]�prax ��M�N��u�b�isd�e܃h�\�iR\P! isbasic���B� P]��QAxes�R6�������.�(Ba�Q�ess��\P���2�D�8@�z�atis���(�{�����~��m��FMc�u�{�
ѩ�MNIS��ݝ�����x����ٺ��jW7}5��Devic��� Interfa�c�RȔQJ7540��� \P�Ne`� �\P�ϐ2�б�����dn� "DNE����
tpdnu�i5UI��ݝ	b�d�bP�q_rs�ofOb
dv_aro��u����>�stchkc���z	 �(}onl��G!ffL+H�@J(��"l"/�n�bx��z�hamp���T�C�!i�a"�59`��S�q��0 (�+�P�o�u�!2��xpc�_2pcchm��C�HMP_�|8бpe�vws��2쳌pc�sF��#C Sen\Pacro�U·�-�R6�Pd�\Pk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GE�M,\i(��Dgesnd�5���H{�}Ha��@sy���c�Isu�xD��Fmd��I��7��4���u���AccuCal�P�4t@��Rɢ7ޠB0��6+56f�6��99\aFF q�S(�U��2�
X�ap�!Bd��cb_��SaUL��  ��t@?�ܖto��ot�plus\tsr�nغ�qb�Wp��t����1��Tool (N. A.)�[K�7�Z�(P�m�����bfclst@k94�"K4p��qt�pap� "PS�9H�stpswo`��p�L7��t\�q ����D�yt5�4�q��@w�q��t@�M�uk��rkey����s���}t�sfeatu�6�EA��t@cf)t\�Xq�����d�h5���LRC0�md�!�C587���aR�(�����2V��8c?u3l\�pa3}H�&r-��Xu���t,�t@�q "�q�Ot��~,���{@�/��1c�}����y�p �r��5���S�XAg��-�y���Wj874��- iRVis<���Queu�t@�Ƒ�-�6�1���(����u���tӑ�����
�tpvtsn? "VTSN�3C�t+�t@v\pRDV����*�prdq\�Q<�&�vstk=P�������nm&_�դ��clrqν���get�TX��Bd����aoQϿ�0qstr�D[t@��t�p'Z��Ɵ�npv��@�enlIP0��D!x�'�|����sc ߸��tv�o/��2�q���v b����q���!���h�]��(� Con�trol�PRAuX�P5��556�A�@59�P56.@5�6@5A�J69�$@982 J55?2 IDVR7�hq A���16�H���La��� ��Xe�f�rlparm.fn�FRL�am��C9�@(F������w6{���A��QJ6�43�t@50�0L�SE
_pVAR� $SGSYSC���RS_UNIT�S �P�2�4tA�T�X.$VNUM_OLD 5�1�| �{�50+�"�` Funct���5tA�� }��`#@�`3�a0��cڂ��9���@HA5נt@�P���(�A ����۶}����ֻ}��bPRb�߶~p{pr4�TPSPI0�3�}�r�10�#;A � t�
`���1���96�����%C�� A�ف��J�bIncr �	����\���1o�5qni4�MNINp	�t@���!���Hour  �� 2�21� �AAVM����0 ��T�UP ��J5�45 ��616�2�VCAM � (�CLI{O ��R6�<N2�MSC "�P �STY�L�C�28~ 13�\�NRE "FwHRM SCH^��DCSU%O�RSR {b�04� �EIOC��1 j 542 �� os| � eg�ist�����7��1�MASmK�934"7 ���OCO ��"3�8��2���� C0 HB��� 4�";39N� Re�� ��LCHK
%OP�LG%��3"%MH�CR.%MC  ; 4l? ��6 dPI�s54�s� DSW%�MD� pQ�K!63!7�0�0p"�1�Р"�4 �6<27 CgTN K � 5 ��%�"7��<25�%/�=T�%FRDM� ��Sg!��930 FB( NBA�P� ( �HLB  Men��SM$@jB( PV3C ��20v��2�HTC�CT�MIL��\@PAC� 16U�hAJ`SA�I \@ELN��<29�s�UECK <�b�@FRM �b�sOR���IPL��}Rk0CSXC ���VVFnaTg@H�TTP �!26� ��G�@ob�IGUI"%IPG�S�r� H863 �qb�!�07r�!34 |�r�84 \so`0! Qx`CC3 Fb�291�!96 rb!g51 ���!53R%� 1!s3!��~�.rp"9js VATFU�J775"��pLR6�^RP�WSMjUCTO�@xT58 F!s80���1XY ta�3!770 ��8�85�UOL  GTS�o
�{` LCM ��r| TSS�EfP6� W�\@CPE �`��0VR� l�QN�L"��@001 i7mrb�c3 =�b0�0���0�`6 w�b^-P- R-�b8n@75EW�b9 �Ґa�� ���b�`ׁ�b2 O2000��`3��`4*5�`5!�c��#$�`7.%�`8 h�605? U0�@B�6E"aRp7� !Pr8 t�a@�tr�2 iB/�1vp3L�vp5 Ȃtr9Σʐa4@-p�r3 	F��r5&�re`u�&�r7 ��r8�U�p9 \h738�a��R2D7"�1�f��2&�7� �3� 7iC��4>w58Ip�Or60 C�L��1bEN�4 I�py�L�uP��@N�-PJ8d�N�8NeN�9 H�(r`�E�b7]�|�⠂8�Вࠂ9 2H��a`0�qЂ5�%?U097 0��@q1�0���1 (�q�3 5R���0 ���mpU��0�0��7*�H@(q�\P"wRB6�q124�b`;��@���@06� 6x�3 pB/x�u ���x�6 H606�a1� ��7 6� ���p�b15�5 ����7jUU1g62 �3 g���4*�65 2ec "_��P�4U1`����B1���`0'�1�74 �q��P�E1�86 R ��P�7� ��P�8&�3 (��90 B/�s1q91����@202��6 3���A�R�U2� d��2 bI2h`��4�᪂2�L4���19v Q�2�*�u2d�Tpt2� ��EH�a2hP�$�5��F�!U2�p�p
�2�p���@5�0-@��84 @�9��TX@�� :�e5�`rb26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0`@�gqGA���a52ѐ��Ḳ6�60ہ5�� ׁ2��8�E��9��EU5@ٰ\�q5�hQ`S�2ޖ5�p\�w�۲�pJ �-P��5��p1\t�H�4��PeCH�7j��phiw��@��P�x��559 ldu� P�D���Q �@������� �`.���P>��8�581l�"�q58�!AM۲�T�A iC�a58�9��@�x����5 �a��12׀0.�1����,�2����,�!P\�h8��Lp ��,�7���6�0840\t}� "T20C}A`��p��{��ran���FRA��Д�� ����A%���ѹ�� ������(����Ѐ� ��З���������������$�G��1���⨂��������� ,e�`q� � �����`64��M���iC/50T-�H������*��)p46��� C��N�����m75s֐� Sp�ѯb46��v��ༀГM-71?�70�З����42����Ȁ�C��-�а�70H�r�E��/h����O$��rD���c7c7C�q���ą���L��/��2\?imm7c7�g� ������`���(� ��e�����"��������a r��c�T,�Ѿ�"��,�� ��xx�Ex�m77t����k���5�����v)�iC��-HS -� B
_�>���+�Т�7U�]���M*h7�s��7������-9?�/260L_������QB�������]�9p�A/@���q�S��х���h6k21��c��92�������.�)92c 0�g$�@�����)$p��5$���pylH"O"
�21���t?�350����p���$�
�� �350!���0��9�U/�0\m9��M9AA3��4%� sё3M$��X%u���"him98J3����� �i d�"m4~�103�p�� �Ӏ�h794̂�&R���H�0���� \���g�5A���Ԝ� �0���*2��00��#06�АՃ���!07{r ����� ���kЙ@����EP�#������?�p�#!�;&07\;!�B1P�߀A��/��CBׂ2�!�:/��?8�ҽCD25L�����0�"l�2BAL
#��B��\20�2 _�r�re���X��1@��N����A@��z��`C�pU��`�#04��DyA�\�`fQ��sU���\��5  ���� p�Dp���<$8�5���+P=�ab1l�1LT��lA�8�!uDnE(�20�T��J�1 e�bH8�5���b�Հ�5[�16Bs��������d�2��x��m6t !`Q����bˀ���b#�(�6iB;S�p�! ��3� ��b�s��-`�_�W8�_���&�6I	$�X5�1�Uc85��R�p6S� ���/�/+q�!�q��`񈓃6o��5m[o)�m�6sW��Q�?��set06p ��3%H�5��10p$����g�/�JrH�� � ��A�856�����F�� ���p/2��� ��܅�✐)�5��̑v��(��m6��Y�H�ѝ̑�m�6�Ҝ��a6�DM�����-S�+��H 2�����Ҽ�� �r ̑��✐��l����p1���F���2�\wt6h T6H�� ��Ҝ�'Vl���� ���V7ᜐ/����;3A7��p~S��������4�`圐�V�T��!3��2�PM[�p�%ܖO�chn��vel5����Vq���_arp#��̑�.�~��2l_hemq$8�.�'�6415��� 5���?����F������5g�L�ј[���1���𙋹1����M7NU�М��eʾ����uq$D;��-�!4��3&H�f�c�Ĝ� h������u�� �㜐��ZS�!ܑ4�&��M-����S�$̑�ք �� 0��<������07shJ�H �v�À�sF��S*� ����̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(UL� &�(�,���0�\�?����̑�a�� ,e�����a�e�w�2ȫ�(�	�2�C��A/����\�+p�����2�1 (ܱ�CL S ����B̺��7F��h�?�<�lơ1L� ���c� ���u9�0����e/q��O���98�K��r9 (��,��Rs�ז�5�G�m20c��i��w�A2��:�0`�$��2�2 l�0�k�X�S� ,�ι�2��O���1!4�1w���2T@� _std��G�y� �ң�<H� jdgm���� w0\� �1L���	�P��~�W*�b��t 5P������3�,����E{������LL��5\L��3��L�|#~���~!���4��#��O����h�L6 A�������2璥���44�����[6\j4s��·��@�#��ol�E"w�8P k�����?0xj�H1�1`Rr�>��]�2a�#2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l��0`�&�"��|�`Am1�2@��ػ��3�HqB ��K�R��ˑb�W� ��Fs���)�ѐ�!����a�1����5��16�16C��C<����0\imBQ���d����b��\B5�-���DiL���O�_�<ѠPEtL�E�RH��ZǠPgω�am1l ��u���̑�b�<����<�$�T�̑�F�����Ȋ�Dpb��X"x��hr��p� ���Dp���9�0\� �j971\kckrcfJ�F�s������c��e "CTM�E�r���ɛ��a�`main.[��g�`Grun}�_vc�# 0�w�1Oܕ_u����bctme��Ӧ�`�ܑ�j735�-� KAREL U�se {�U���J���1���p� U ̑�9�B@��L�9����7j[�atk208 "K��Kя��\��9��a��̹�����cKRC�a�o ��kc�qJ�&s��� ��Grſ�fsD��:y�0�s��A1X\j|хr�dtB�, ��`.	v�q�� �sǑIf��Wfj52�TKQu�to Set��J�� H5K536�(�932���91�5�8(�9�BA�1(�7�4O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v���! conre;a�#�Controlw Re�ble��CNRE(�T�<�4��2���D�)���S�55i2��q(g�� (����4X�cOux�\s�futs�UTS `�i�栜���t�棈���? 6�T�!�S#A OO+D6����������,!��6�c+� igt�t6iB��I0�TW8 �0��la��vo58�o�b@Få򬡯i�Xh���!Xk�0Y!8\m6e�!6EC���v��6���������<1!6�A���A�6s��ƀ�U�g�T|ώ���rE1�qR��˔Z4�T������,#�eZp)g ����<ONO0���uJ���tCR;��F�a� �,e��f��prdsuchk �1���2&&?���t��*D %$�r(�✑�娟:r���'�s�qO��<s�crc�C�\At�trldJ"o�\�V�|���Paylo�nfirm�l�!�87��7��A�3ad�! �?ވI�?hplQ��3��3"�q��x pl�`���d87��l�calC�u�Du���;��movx�����initX�:s8O��a�r4 ���r67A4|�e GeneratiڲĐ��7g2q$��g =R� (Sh��c ,|�bE��$ԒA\�:�"��4���4�4�. sg��5��F$d6"e;Qp? "SHAP�T�Q ngcr pGC��a(�&"� ��"G3DA¶��r6�"�aW�/�$dataxX:s�"tpad��<[q�%tput;a__�O7;a�o8�1�yl+s��r�?�:�#�?�5x$�?�:c O�:y O�:H�IO�s`O%g�q�ǒ�?�@0\��"o�j�92;!�Ppl.C�ollis�QSkip#��@5��@J��D ��@\ވ�C@X��7��7�|s2��potcls�LS��DU�k?�\_ et1s�`�< \�Q䜐�@���`dcKqQ�F�C;��J,�n��` (��4eN����T�{���'j(�c������/IӸaȁ��̠GH�����зa��e\mcclmt "CLM�/��� �mate\��lmpALM�?>p7qCmc?����2vm�qp��%�3s��_sv90<�_x_msu�2L�^v_� K�o�{in��8(3r<�c_lo�gr��rtrcW� �v_3�~yac��d�<�ten��der$cCe�' Fiρ�R��Q��?�l�enteAr߄|��(Sd��V1�TX�+fK�r�a�99sQ9+�5�r�\tq\� "FN�DR���S�TDn$LAN]G�Pgui��D�`���S������sp�!ğ֙uf�ҝ�s����$�����e+�=�� �������������w�H�r\fn_�ϣ��|$`x�tcpma��- TCP�����?R638 R�Ҭ���38��M7p, ���Ӡ�$Ӡ�8p0Р��VS,�>�tk��99 �a��B3���PզԠ��0D�2�����UI��t� ��hqB���8��������p���re�ȿ��exe@4φ�B���pe38�ԡG�rmpWXφ�var@�φ�@3N�����vx�!ҡ���q�RBT �$cOPTN ask E0��1��R MAS0�H5�93/�96 H5�0�i�480�5�H0��m�Q�K��7�0�g�Pl�h0ԧ�2���DP��@"��_t\mas��0�a@��"�ԧ�����k�� �R����ӹ`m��bL��7�.f��u�d���r��splay�D�E���1w�UPD�T Ub��887 M(��Di{���v�� ��Ԛ⧔��#�B���|����o  ��� �a�䣣��60q��B�����qscan0��B���ad@�������q`�䗣��#��К�`2�� vl v��Ù�$�>�b����! S��Easyy/К�Util��|룙�511 J������R7 ��Nor|֠��inc),<6Q�� �`c��"4�[���986FVRx� So����q�nd 6����P��4�a\ (�@�
  �������d���K�bdZ���men�7���- Me`t!yFњ�Fb�0�T�Ua�577?i 3R��\�5�u?��!� n���f���<���l\mh�Ц�pűE|hmn�	���<\O���eD�1�� l!��y��Ù�\|p����B���Ћmh�@��:. aG!���/�t��55�6�!X�l�.u�s��Y/k)ensu)bL���eK�h��  �B\1;5g?y?�?�?D��?*rm�p�?Ktbox O2K|?0�G��C?A%ds���?�P"�!� �TR�� /��P�T6@�`�U�P�V�P�Ue�P0�U�PO��\3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ăd�Q3t.�P׀al��P+OP517F��IN0a��Q(}g���PESTf3ua@�PB�l�ig�h�6�a�q��P � ,9e��`  n�0m�bumpP�Q969g�69�Qq��P0��baAp�@Q� B�OX��,>vche8�s�>vetu㒣^=wffse�3�Ā�]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q8<twaǂ tp�Q҄�Taror Re'cov�b�O�P�642����a�q���a⁠QErǃ�Qr!y��`�P'�T�`�a�ar������	{'�paok971��71��`m���>��`jot���PXc��C�1�adb �-�ail��nagx���b�QR629�a�Q��b�P  ��
  �P���$$CL[q �����������$�PS_DIGsIT���"�!�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*���1:PRODU�CT�Q0\PGS�TK�bV,n��99�����$FEAT_IN�DEX��~������IL�ECOMP ;���)��"��S�ETUP2 <����  �N !�_AP2�BCK 1=�  �)}6/E+%,/i/��W/�/ ~+/�/O/�/s/�/? �/>?�/b?t??�?'? �?�?]?�?�?O(O�? LO�?pO�?}O�O5O�O YO�O _�O$_�OH_Z_ �O~__�_�_C_�_g_ �_�_	o2o�_Vo�_zo �oo�o?o�o�ouo
 �o.@�od�o� ��M�q��� <��`�r����%��� ̏[�������!�J� ُn�������3�ȟW� �����"���F�X�� |����/���֯e��� ���0���T��x��� ���=�ҿ�s�ϗ�@,ϻ�9�b�� P/� 2) *.V1Riϳ�!�*����`������PC�|7�!�FR6:"�"c��χ��T��� ��Lը��ܮx��ﶏ*.F��>� �	�N�,�k��ߏ��STM �����Qа����!�iPen�dant Panel���H��F����4������GIF �������u����JPG&P��<�����	PANE�L1.DT��@������2��Y�G��
3 w�����//�
4�a/�O///�/��
TPEINSO.XML�/����\�/�/�!Cust�om Toolb�ar?�PAS�SWORD/��FRS:\R?? �%Passwo�rd Config�?��?k?�?OH� 6O�?ZOlO�?�OO�O �OUO�OyO_�O�OD_ �Oh_�Oa_�_-_�_Q_ �_�_�_o�_@oRo�_ voo�o)o;o�o_o�o �o�o*�oN�or� �7��m�� &���\�����y� ��E�ڏi������4� ÏX�j��������A� S��w�����B�џ f�������+���O�� �������>�ͯ߯t� ���'���ο]�򿁿 �(Ϸ�L�ۿpς�� ��5���Y�k� ߏ�$� ���Z���~�ߢߴ� C���g�����2��� V����ߌ���?�� ��u�
���.�@���d� �����)���M���q� ����<��5r �%��[� &�J�n�� 3�W���"/� F/X/�|//�/�/A/ �/e/�/�/�/0?�/T? �/M?�??�?=?�?�? s?O�?,O>O�?bO�? �OO'O�OKO�OoO�O _�O:_�O^_p_�O�_ #_�_�_Y_�_}_o�_��_Ho)f�$FIL�E_DGBCK �1=��5`��� ( ��)
SUMMA�RY.DGRo�\�MD:�o�o
`�Diag Sum�mary�o�Z
C?ONSLOG�o�o�a
J�aCon�sole log�K�[�`MEMCHECK@'�o��^qMemory� Data��W��)�qHAD�OW���P��s�Shadow C?hangesS�-c�-��)	FTAP=��9����w`q�mment TB�D׏�W0<�)�ETHERNET�̏�^�q�Z��aE�thernet �bpfigurat�ion[��P��DCSVRFˏ��Ïܟ��q%�� ve�rify all�ߟ-c1PY���DIFFԟ��̟a��p�%��diffc���q��1X�?�Q��� ����X=��CHGD��¯ԯi��px��� ����2`�G�Y�� ��� �GD��ʿܿ�q��p���Ϥ�FY�3h�O�a��� ��(�GD�������y��p�ϡ�0�UPDATES.������[FRS:\������aUpda�tes List����kPSRBWLOD.CM.��\���B��_pPS_ROBOWEL���_�� ��o��,o!�3���W� ��{�
�t���@���d� ����/��Se�� ���N�r � =�a�r� &�J���/� 9/K/�o/��/"/�/ �/X/�/|/�/#?�/G? �/k?}??�?0?�?�? f?�?�?O�?OUO�? yOO�O�O>O�ObO�O 	_�O-_�OQ_c_�O�_ _�_:_�_�_p_o�_ o;o�__o�_�o�o$o �oHo�o�o~o�o7 �o0m�o� �� V�z�!��E�� i�{�
���.�ÏR��� �������.�S��w� �����<�џ`���� ��+���O�ޟH�������8���߯n�����$FILE_��P�R���������� �M�DONLY 1=�4�� 
 � ��w�į��诨�ѿ�� �����+Ϻ�O�޿s� ��ϩ�8�����n�� ��'߶�4�]��ρ�� �߷�F���j����� 5���Y�k��ߏ��� B�����x����1�C� ��g������,���P� ��������?��L�u�VISBCK�R�<�a�*.VD�|�4 FR:\���4 Vis�ion VD file� :Lb pZ�#��Y� }/$/�H/�l/� /�/1/�/�/�/�/�/  ?�/1?V?�/z?	?�? �???�?c?�?�?�?.O �?ROdOO�OO�O;O �O�OqO_�O*_<_�O�`_�O�__%_�_�M�R_GRP 1>�4�L�UC4 w B�P	 ]��ol`�*u����RHB ���2 ��� ��� ���He �Y�Q`orkbIh�oJd�o�Sc�o�oK��~�I�H�I޿�WF�5U�aR�!�`�o�o^`��4�EŰC ��ףQ7�Z/<��w!}>j!��>��lq�Q>|��U>���}E�� F@ �r��d�a}J��NJ�k�H9�H�u��F!��IP�s}?�`�.�9�<9��896C'�6<,6\b��  Au�_B�W��Ay;A?��@B{-��5�BlA1xA�7h��H���, A1�� ����|�ݏx���%���  @Ì�A�E�5@U�U@���4���j��� ��ǟ���֟��!���E�`r�UBH�P� �a`�Q�l�(v�K���ï�T
6�PQ��PQ��˯`�o�e�Q cB��P<5���@�33@����4�m�,�@UUU�U�~w�>u.�?!��]��տ����2��=[z�=��̽=V6<��=�=�=�$q��~��@8��i7G��8��D�8@9!�o��϶ϡ������D�@ D�� SCϫo4z��P��P'�6��_V� m�o�� To��xo�ߜo����� �A�,�e�P�b��� �����������=� (�a�L���p������� ����������*��N 9r]����� ���8#\n Y�}������ �/ԭ//A/�e/P/ �/p/�/�/�/�/�/? �/+??;?a?L?�?p? �?�?�?�?�?�?�?'O OKO6OoO�OHߢOl� �ߐߢ��O�� _��G_ bOk_V_�_z_�_�_�_ �_�_o�_1ooUo@o yodovo�o�o�o�o�o �oNu �������� �;�&�_�J���n��� ����ݏȏ��%�7� I�[�"/�描����� ٟ�������3��W� B�{�f�������կ�� �����A�,�e�P� b��������O�O�O ��O�OL�_p�:_�� ���Ϧ��������'� �7�]�H߁�lߥߐ� �ߴ�������#��G� 2�k�2��Vw���� �������1��U�@� R���v����������� ��-Q�u� ��r��6�� )M4q\n� �����/�#/ I/4/m/X/�/|/�/�/ �/�/�/?ֿ�B?� f?0�BϜ?f��?���/ �?�?�?/OOSO>OwO bO�O�O�O�O�O�O�O __=_(_a_L_^_�_ �_�_���_��o�_o 9o$o]oHo�olo�o�o �o�o�o�o�o#G 2kV{�h�� �����C�.�g� y�`����������Џ ���?�*�c�N��� r��������̟�� )��M�_�&?H?���? ���?�?�?����?@� I�4�m�X�j�����ǿ ���ֿ����E�0� i�Tύ�xϱϜ����� ����_,��_S���w� b߇߭ߘ��߼����� ��=�(�:�s�^�� ���������'� 9� �]�o����~��� ����������5  YDV�z��� ���1U@ yd��v����� /Я*/��
/�u/� �/�/�/�/�/�/�/? ?;?&?_?J?�?n?�? �?�?�?�?O�?%OO IO4O"�|OBO�O>O�O �O�O�O�O!__E_0_ i_T_�_x_�_�_�_�_ �_o�_/o��?oeowo �oP��oo�o�o�o �o+=$aL�p �������'� �K�6�o�Z������ ɏ��폴� ��D� / /z�D/��h/ş�� �ԟ���1��U�@� R���v�����ӯ���� ��-��Q�<�u�`� ��`O�O�O���޿� �;�&�_�J�oϕπ� �Ϥ��������%�� "�[�F��Fo�ߵ��� �ߠo��d�!���W� >�{�b�������� ������A�,�>�w� b����������������=��$FN�O ����\�
�F0l q  FL�AG>�(RRM�_CHKTYP � ] ��d ��] ��OM� _�MIN� 	����� �  XT S�SB_CFG �?\ ����O�TP_DEF_O/W  	��,�IRCOM� >��$GENOVRD7_DO��<�l�THR� d�d�q_ENB] �qRAVC_GR�P 1@�I X(/ %/7//[/ B//�/x/�/�/�/�/ �/?�/3??C?i?P? �?t?�?�?�?�?�?O OOAO(OeOLO^O�O.oROU�F\� �,�B,�8�?���O�O��O	__���  DaE_�Hy_�\@@m_B�=�vR/��I�O�WSMT�G�SU�oo&oRHOST�C�1H�I� Ĺ�zMSM��l[bo�	1�27.0�`1�o  e�o�o�o #z�oFXj|�l6�0s	anonymous�����F�Jao�&�&��o�x��o������ ҏ�3��,�>�a� O����������Ο�U %�7�I��]����f� x��������ү��� �+�i�{�P�b�t��� ���������S� (�:�L�^ϭ�oϔϦ� �������=��$�6� H�Zߩ���Ϳs����� ������ �2���V� h�z��߰������� ��
��k�}ߏߡߣ� ���߬���������C� *<Nq�_�� ����-�?�Q�c� eJ��n���� ���/"/E� X/j/|/�/�/� %'/?[0?B?T?f? x?��?�?�?�?�?? E/W/,O>OPObO�KDa�ENT 1I�K� P!�?�O  �P�O�O�O�O�O#_ �OG_
_S_._|_�_d_ �_�_�_�_o�_1o�_ ogo*o�oNo�oro�o �o�o	�o-�oQ u8n����� ���#��L�q�4� ��X���|�ݏ���ď�֏7���[���B�?QUICC0��h�z�۟��1ܟ��ʟ+��2,���{�!?ROUTER|�X��j�˯!PCJO�G̯��!19�2.168.0.�10��}GNAME� !�J!RO�BOT�vNS_C�FG 1H�I ��Aut�o-starte�d�$FTP�/ ���/�?޿#?��&� 8�JϏ?nπϒϤ�ǿ ��[������"�4ߵ& ����������濜��� �������'�9�K�]� o����������� ��/�/�/G���k��� �������������� 1T���Py�� ���"�4�	H- |�Qcu�VD� ���/�;/M/ _/q/�/����/
/ �/>?%?7?I?[?*/ ?�?�?�?�/�?l?�? O!O3OEO�/�/�/�/ �?�O ?�O�O�O__ �?A_S_e_w_�O4_._ �_�_�_�_oVOhOzO �O�_so�O�o�o�o�o �o�_'9Kno �o�����o*o <oNoP5��oY�k�}� ����pŏ׏���� 0���C�U�g�y���_��T_ERR J�;�����PDUSI�Z  ��^P�����>ٕWRD �?z���  �guest ���+�=�O�a�s�*��SCDMNGRPw 2Kz�Ð���۠\��K��� 	P01.�14 8�q  � y��B    ;�����{ �����������������������~ �ǟI�4�m�X��|��  i�  �  
����� ����+��������
����l�.x��
��"�l�ڲ۰s��d�������_G�ROU��L�� e��	��۠07K�QUPD  ����PČ�TYg������TTP_A�UTH 1M��� <!iPen'dan���<�_��!KAREL�:*�����KC�%�5�G��VISION SETZ���|��Ҽߪ��� ������
�W�.�@����d�v���CTRL� N�������
��FFF9E�3���FRS:DEFAULT��FANUC �Web Server�
������q�������������W�R_CONFIGw O�� ����IDL_CPU�_PC"��B���= �BH#MI�N.�BGNR_�IO��� ���% N�PT_SIM_D�Os}TPMO_DNTOLs �_PRTY�=!OLNK 1P���'9K]|o�MASTEr ������O_CFG���UO����C�YCLE���_?ASG 1Q���
 q2/D/V/h/ z/�/�/�/�/�/�/�/p
??y"NUM����Q�IPCH���£RTRY_�CN"�u���SC�RN������ ���R����?���$J23_D_SP_EN������0OBPROC��3��JOGV�1�S_�@��8��?�';ZO'??0CP�OSREO�KANJI_�Ϡu�A$#��3T ���E�O�ECL_LM B2e?��@EYLOGGI�N�������L�ANGUAGE Y_�=� }Q���LG�2U������ �x�����PZC � �'0������MC:\RSCH\00\˝�LN_DISP V�������T�OC�4Dz\A��SOGBOOK W+��o���o�o���Xi�o�o�o�o��o~}	x(y��	�ne�i�ekElG�_BUFF 1X���}2���� Ӣ������'� T�K�]����������� ɏۏ���#�P���~�qDCS Zxm =���%|d1h�`���ʟܟ�g�IOw 1[+ �?'����'�7�I�[�o� �������ǯٯ��� �!�3�G�W�i�{��������ÿ׿�El TM  ��d��#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U��g�yߋߝ߈t�SE�V�0m�TYP�� ��$�}�A�RS"�(_�s�2FLg 1\��0��� �����������5�STP<P���DmNGNAM�4�U�nf�UPS`GI�5��A�5s�_LOA�D@G %j%=@_MOV�u�����MAXUALRMB7�P8��y���3��0]&q��Ca]�s�3�~�� 8@=@^�+ طv	��V0+�P�A5d�cr���U� �����E( iTy����� ��/ /A/,/Q/w/ b/�/~/�/�/�/�/�/ ??)?O?:?s?V?�? �?�?�?�?�?�?O'O OKO.OoOZOlO�O�O �O�O�O�O�O#__G_ 2_D_}_`_�_�_�_�_ �_�_�_o
ooUo8o yodo�o�o�o�o�o�o��o�o-��D_LDXDISA^�� �MEMO_APX��E ?��
 �0y�����������ISC ;1_�� �O� ���W�i�����Ə �����}��ߏD�/� h�z�a��������� �����@���O�a� 5������������u� �ׯ<�'�`�r�Y��� ���y�޿�ۿ��� 8Ϲ�G�Y�-ϒ�}϶� ������m�����4���X�j�#�_MSTR� `��}�SCD 1as}�R���N� �������8�#�5�n� Y��}��������� ���4��X�C�|�g� �������������� 	B-Rxc�� �����> )bM�q��� ��/�(//L/7/ p/[/m/�/�/�/�/�/ �/?�/"?H?3?l?W?��?{?�?�?�?n�MK�CFG b����?��LTARM_��2cRuB� �3WpTNBpME�TPUOp�2�����NDSP_CM�NTnE@F�E�� d���N�2A�O|�D�EPOSCF�G��NPSTOL �1e-�4@�<#�
;Q�1;UK_YW7_ Y_[_m_�_�_�_�_�_ �_o�_oQo3oEo�o�io{o�o�a�ASIN�G_CHK  ��MAqODAQ2Cf�O�7J�eDEV �	Rz	MC:>'|HSIZEn@�����eTASK �%<z%$1234?56789 ��u��gTRIG 1g.�� l<u%����3���>svvYP�aq��kEM_IN�F 1h9G� `)AT?&FV0E0(����)��E0V1&�A3&B1&D2�&S0&C1S0}=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏ P��t�������]�ί �����(�۟�^� �#�5�����k�ܿ�  ϻ�ů6��Z�A�~� ��C���g�y������ ��2�i�C�h�ό�G� ���ߩ��ߙϫ���� ����d�v�)ߚ��߾� y��������<�N� �r�%�7�I�[���� ��9�&��J[��g��>ONIT�OR�@G ?;{ �  	EXESC1�3�2�3�E4�5��p�7�8�9�3�n�R �R�RRR R(R4R@RTLR2Y2e2qU2}2�2�2�U2�2�2�3Y�3e3��aR_G�RP_SV 1i�t��q(�?�/�e~q_�DCd~�1PL_N�AME !<u�� �!Defa�ult Pers�onality �(from FD�) �4RR2k! �1j)TEX)TsH��!�AX d�/ >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO@^OpO�O�O�Ox2-? �O�O�O__0_B_T_f_x_�b<�O�_�_�_ �_�_�_o o2oDoVotho&xRj" 1o�)�&0\�b, ��9��b�a @D��  �a?��c�a?x�`�a�aA'�6�e�w;�	l�b	� �xJp��`�`	p� �< ��(p� �.r� K��K ��K=�*�J���J���JV��kq`�q�P�x�|� @j�@T;f�r��f�q�acrs�I�����p����p�r�ph}�3��´  ���>��ph�`z���Ꜭa��3Jm�q� H�N���ac��'�aw�� ~ �  P� �Q� �� |  �а��/Ώqu	'�� � �I�� �  ��ވ�:�È�È�=���(����a	����I  �n @H�i~�ab�ӋB�b��w����N0��  'Ж�q�p�@2��@���X�r�q5�C�pC0C�@ C���=�`
�A1q "  @B�UV~X�
nwB0"h�A��p�ӊ�p�`���aDz���֏����Я	�pv�( �� -���I��-�=��A�a��we_q�`�p �?�ff ��m��>� ����Ƽ���@ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`���<
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC��������#/*/c/N/�wi�����v/C�`� CHs/`
=$�p��<!�!��ܼ�'��3A�A�AR�1AO�^?�$��?��] ±�
=ç>�����3�W
=�#��]�;e�׬a@�����{�����<�>(��B�u���=B0�������	R��zH�F��G���G���H�U`E����C�+��}I�#�I��H�D�F��E���RC�j=�>
�I��@H��!H�( E<YD0w/O*O ONO9OrO]O�O�O�O �O�O�O�O_�O8_#_ \_G_�_�_}_�_�_�_ �_�_�_"oooXoCo |ogo�o�o�o�o�o�o �o	B-fQ� u������� ,��P�b�M���q��� ��Ώ���ݏ�(�� L�7�p�[������ʟ ���ٟ���6�!�Z��E�W���#1(|��ٙ9�K���ĥ|������Ư!3��8���!4Mgqs��,�IB+8��J��a���{�d�d�����ȿ��쿔ڼ%P��P�= :GϚ�S�6�h�z���R�Ϯ����������  %�� ��h� Vߌ�z߰�&�g�/9�$�������7�����A�S�e�w�   ������������̿2 F�$�&Gb��������!C���@��������8�F� Dz�N�� F�P �D�������)#�B�'9K]o#?_���@@v
0ԥ8�8��8�.
 v��� !3EWi{�����:� ���ۨ�1��$M�SKCFMAP � ���� ���(.�ONREL  ��!9��EXC/FENBE'
#7%�^!FNCe/W$JO�GOVLIME'dtO S"d�KEYE'u�%�RUN�,��%�SFSP�DTY0g&P%9#S�IGNE/W$T1M�OT�/T!�_C�E_GRP 1p��#\x��?p� �?�?�?�?�?O�? OBO�?fOO[O�OSO �O�O�O�O�O_,_�O P__I_�_=_�_�_�_ �_�_oo�_:o��TCOM_CFG 1q	-�vo�o��o
Va_ARC_�b"�p)UAP_�CPL�ot$NOCHECK ?	+ �x�% 7I[m���������!�.+N�O_WAIT_L� 7%S2NT^ar�	+�s�_ERR�_12s	)9��  ,ȍޏ��x����&��dT_MO��t>��, W�*oq��9�PARAM��u	+��a�ß'g�{�� =?�345?678901�� ,��K�]�9�i�����`��ɯۯ��&g������C��cUM_RSPACE/�|�����$ODRDS�P�c#6p(OFFSET_CART�oη�DISƿ��PE?N_FILE尨!��ai��`OPTIO�N_IO�/��PW�ORK ve7s# ��V�ؤ�p�p�4�p�	 ���p��<���RG_DSBL  ���P#��ϸ�RIE�NTTOD ?�Cᴭ !l�UT__SIM_D$�"����V��LCT w}�h�iĜa[�1ԟ_PEXE�j�R�ATvШ&p%� ��2�^3j)TEX)T�H�)�X d 3�������%�7�I� [�m��������������!�3�E��2 ��u���������������c�<d�AS ew������`��Ǎ�^0OUa0�o(��(�����u2, ����O H @D��  [?�aG?��cc�D][�Z��;�	ls��xJ��������<� ��� ���2�H(��H3�k7HSM5G��22G���Gpc
͜�'f�/,-,2�CR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t3�!�/ �/�"�t32����/6 W ��P%�Q%��%�|T��S62�q?�'e	'� � ��2I� � � ��+==�̡ͳ?�;	�h	�0��I  �n �@�2�.��Ov;���ٟ?&gN�]O  �''�uD@!� C�C��@F#H!�/�O�O Nsb
���@�@E��@�e`0B��QA�0Yv: �13Uwz$oV_�/z_�e_�_�_	��( �� -�2@�1�1ta�Ua�c����:A-���.  �?�ff���[o"o�_!U�`oXÜQ8���o:�j>�1  Po�V(���eF0�f�Y����e�?����x�b�P<
6b<�߈;܍�<��ê<� <�#&�,/aA�;r��@Ov0P?fff?��0?&ip�T@�.�{r�J<?�`�u#	�Bdqt�Yc �a�Mw�Bo�� 7�"�[�F��j����� ��ُ����3�����,���(�E��� E��3G+� F��a��ҟ������,��P�;���B�pAZ�>��B��6�<O ίD���P��t�=����a�s�����6j�h�y�7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�<%?��?������(���#	Ę��P �N�||CH���Ŀx������@I�_��'�3A�A�A�R1AO�^??�$�?��� ��±
=ç>�����3�W
=�#� U��e����B��@��{�����<����(�B�u���=B0�������	�b�H��F�G���G���H�U`E����C�+��I�#�I��H�D�F��E��RC�j=[��
I��@H��!H�( E?<YD0߻� �������� �9�$� ]�H�Z���~������� ������#5 YD }h������ �
C.gR� ������	/� -//*/c/N/�/r/�/ �/�/�/�/?�/)?? M?8?q?\?�?�?�?�? �?�?�?O�?7O"O[O mOXO�O|O�O�O�O�O��O�O�O3_Q(���3���b��gUU���W_i_2�3ǭ8��_�_2�4M�gs�_�_�RIB+��_�_�a���{�miGo5okoYo(�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�u�,��  �p���o ��/��S��z
uү ܠ�������ڱ������������  /�M�w�e�������~�l2 F�$��'Gb��t��a�`�,p�S�C�y�@p�5��G�Y�۠F� D�z�� F�P D��]����پ��ʯܯ� ��~ÿ?���@@�J?�K�K���K���
 �|��� ����Ŀֿ������0�B�T�fϽ�V� ����{��1��$�PARAM_ME�NU ?3���  �DEFPULS�Er�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L��	�OPT���PTB4�.�C��R_DECSN ���e��ߑߣ����� ������!�3�\�W��i�{���USE_PROG %��q%�����CCR����e����_HOSoT !��!��:���T�`�V��/��X����_TIMqE��^��  ��?GDEBUG\�����GINP_FL'MSK����Tfp�����PGA  ��̹�)CH����TY+PE������� ����� - ?hcu���� ���//@/;/M/ _/�/�/�/�/�/�/�/��/??%?7?`?��W�ORD ?	=�	RSfu	P�NSUԜ2JO�K�DRTEy�]T�RACECTL �1x3��� }�`) &�`��`�>�6DT Q�y3�%@�0D �� �c��a:@V�@BR��2ODOVOhOzO�B �O�O�O�O�O�O�O_"_4_F_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����� ����0�B�T�f� x���������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�.Iv����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p��j��� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o��o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*���$PGTRACELEN  )��  ���(��>�_UP �z���m��u�Y�n�>�_C�FG {m�W�(�~���PКӂ��DEFSPD e|��'�P��>��IN��TRL �}��(�8����PE_CONFI��}~m��m�r���ղ�LID�����=�GRP s1��W��)��A ���&ff�(�A+33D��� D]� CÀ� A@1��Ѭ(�d�Ԭ��0�0�� 	 1�ح֚���G ´�����B� 9����O�9�s�(��>�T?�
5�������� =��=#�
���� P;t_��������  Dz (�
H�X ~i������ /�/D///h/S/�/���
V7.10�beta1��  A�E�"�ӻ�A (�� ?�!G��!>��r�"����!���!oBQ��!A\� P�!���!2p����Ț/8?J?\?n?};� ���/��/�?}/ �?�?OO:O%O7OpO [O�OO�O�O�O�O�O _�O6_!_Z_E_~_i_ �_�_�_�_�_�_'o 2o�_VoAoSo�owo�o �o�o�o�o�o.�R=v1�/�#F@ �y�}��{m��y =��1�'�O�a��? �?�?������ߏʏ� �'��K�6�H���l� ����ɟ���؟�#� �G�2�k�V���z��� �����o��ίC� .�g�R�d��������� �п	���-�?�*�c� ����Ϯ���� ��B�;�f�x����� ��DϹ��߶������ ��7�"�[�F�X��|� �����������!�3� �W�B�{�f������� �� �����/S >wbt���� ��=Ozό� �ψ����ϼ� / .�'/R�d�v߈߁/0 �/�/�/�/�/�/�/#? ?G?2?k?V?h?�?�? �?�?�?�?O�?1OCO .OgORO�OvO�O�O�� �O�O�O__?_*_c_ N_�_r_�_�_�_�_�_ o�_)oTfx�to ���/�o/ >/P/b/t/mo�| �������3� �W�B�{�f�x����� Տ�������A�S� >�w�b����O��џ�� ����+��O�:�s� ^�������ͯ���ܯ �@oRodo�o`��o�o �o��ƿ�o���*< N�Y��}�hϡό� �ϰ��������
�C� .�g�Rߋ�v߈��߬� ����	���-��Q�c� N�ﲟ���l����� ���;�&�_�J��� n�����������,� >�P�:L������� �����(�:�3 ��0iT�x�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?a?s? ��?�?X?�?�?�?�? O'OOKO6OoOZO�O ~O�O�O�O�O*\ &_8_r���_�_���$PLID_K�NOW_M  ~�� Q��TSV ��]�P��? o"o4o�OXoCoUo�o� R�SM_GRP� 1��Z'0{`J�@�`uf�e�`
�5� �gpk 'Pe]o�� ��������S+MR�c��mT�EyQ}? yR�������� ��폯���ӏ�G�!� �-������������ ����ϟ�C���)� ����������寧����QST�a1 1�j�)���P0� A 4��E2�D�V� h�������߿¿Կ� ��9��.�o�R�d�v�@���ϬϾ����2�90� Q�<3��A3�/�A�S��4l�~ߐߢ��5���������6
��.�@��A7Y�k�}���8���������MAD � )��P�ARNUM  �!�}o+��SCH
E� S�
��f���S��UPDf�x�|�_CMP_�`�H�� �'�UE�R_CHK-�a��ZE*<RSr��_�Q_MOG����_�X�_RES_G��!���D� >1bU�y�� ���/�	/����+/�k�H/g/ l/��Ї/�/�/�	� �/�/�/�X�?$?)? ���D?c?h?����?x�?�?�V 1��U��ax�@c]�@t�@(@c\�@��@D@c[�*@���THR_INR�r�J�b�Ud2FMA�SS?O ZSGMN�>OqCMON_QU?EUE ��U�V� P~P X�N$ U�hN�FV�@END8�A��IEXE�O�E���BE�@�O�COP�TIO�G��@PR�OGRAM %��J%�@�?���BT�ASK_IG�6^O?CFG ��Oz���_�PDATA�c�.�[@Ц2=�Do Vohozo�j2o�o�o�o �o�o);M j�INFO[��m� �D������ ��1�C�U�g�y��� ������ӏ���	�dwpt�l )�QE ?DIT ��_i�>�^WERFLX	C��RGADJ M�tZA�����?נ�ʕFA��IORIT�Y�GW���MPD�SPNQ����U�G�D��OTOE@1��X� (!A�F:@E� c�Ч!�tcpn���!�ud����!i�cm���?<�XY_��Q�X���Q)�� *�1�5��P��]�@�L���p��� �����ʿ��+�=Ϡ$�a�Hυϗ�*��P�ORT)QH��P��E��_CART�REPPX��SK�STA�H�
SSA�V�@�tZ	25?00H863���_�x�
�'��X�@�swPtS�ߕߧ���/URGE�@B��x	WF��DO�F"[�W\�������WRU�P_DELAY ��X���R_HO�TqX	B%�c���R_NORMALq^xR��v�SEMI�������9�QSKIP�'��tUr�x 	7�1�1��X�j�|� ?�tU������������ ��$J\n4 ������� �4FX|j� ������/0/ B//R/x/f/�/�/�/�tU�$RCVTM�$��D�� DCR�'���Ў!7���.1�Cc>��)�>�z�;��Z:��O8���j������:�o?�� <
�6b<߈;����>u.�??!<�&�?h? �?�?�@>��?O O2O DOVOhOzO�O�O�O�O �O�?�O�O__@_+_ =_v_Y_�_�_�?�_�_ �_oo*o<oNo`oro �o�o�o�_�o�o�o�o �o8J-n��_ �������"� 4�F�X�j�U������ ď���ӏ���B� T��x���������ҟ �����,�>�)�b� M������������ï կ�Y�:�L�^�p��� ������ʿܿ� �� ��6�!�Z�E�~ϐ�{� �ϗ�����-�� �2� D�V�h�zߌߞ߰��� ������
���.��R� =�v��k������ ����*�<�N�`�r� ������������� ��&J\?�� ������"�4FXj|��!G�N_ATC 1��	; AT�&FV0E0��ATDP/6/�9/2/9�A�TA�,A�T%G1%B96}0�+++��,�H/,�!IO�_TYPE  �%�#t�REFPOS1 1�V+� x�u/� n�/j�/
=�/�/�/ Q?<?u??�?4?�?X?x�?�?�+2 1�V+�/�?�?\O�?�O�?�!3 1�O*O<O�vO�O�O_�OS4 1��O�O�O_�_t_|�_+_S5 1�B_�T_f_�_o	oBo�_S6 1��_�_�_5o�o�o�oUoS7 1�lo~o�o�oH3l>�oS8 1��%_���SM�ASK 1�V/ � 
?�M��XNO�S/�r������!MOTE  n��$��_CFG �����q���"PL_RA�NG�����POW_ER ������SM_DRYP_RG %o�%��P��TART ���^�UME_P�RO-�?����$_E�XEC_ENB � ���GSPD���Րݘ��TDB���
�RM�
�MT�_'�T����O�BOT_NAME� o����O�B_ORD_NU�M ?�b!�H863  a�կ����PC_TIMEO�UT�� x�S2�32Ă1�� �LTEACH PENDAN���w��-���Maintena�nce Consȡ��s�"���KCL/Cm��

����t�ҿ No Use-��Ϝ��0�NPO�򁋁���.�CH_�L������q	���s�MAVAILȶ����糅��SPACE1 2��, j�߂�D��s��߂� �{S�8�?�k�v�k�Z� ���ߤ��ߚ� �2� D���hߊ�|��`��� ������� �2� D��h��|���`���������y���2�� ��0�B���f������{���3 );M_�� ����/� /44FXj|*/� ��/�/�/?(??=?5Q/c/u/�/�/G? �/�/�?O�?$OEO,OZO6n?�?�?�?�? dO�?�?_,_�OA_b_I_w_7�O�O�O�O �O�_�O_(oIoo^oofo�o8�_�_�_ �_�_�oo6oEf)�{���G ��o� ���
M� ���*�<� N�`�r�������w��@�o�収���d.� �%�S�e�w������� ����Ǐَ���Θ8� +�=�k�}�������ů ׯ͟����%�'�X� K�]���������ӿ忀�����#�E�W�; `� @���@����x�����\�e� ����������R�d� ��8�j߬߾߈ߒߤ� ���������0�r�� ��X������������8����
�ύ��_MODE  ��{��S ��{|�2�0�����3��	S|)CWO�RK_AD��D{+R  �{��`� �� _INOTVAL���d����R_OPTION�� ��H VA�T_GRP 2���up(N�k|�� _�����/0/ B/��h�u/T� }/�/ �/�/�/�/�/?!?�/ E?W?i?{?�?�?5?�? �?�?�?�?O/OAOO eOwO�O�O�O�OUO�O �O__�O=_O_a_s_ 5_�_�_�_�_�_�_�_ o'o9o�_Iooo�o�o Uo�o�o�o�o�o�o 5GYk-��� u�����1�C� �g�y���M�����ӏ 叧�	��-�?�Q�c� ��������������ǟ�;�M�_�����$SCAN_TI�M��_%}�R ��(�#((��<04Jd d 
!D�ʣ��u�/���V��U��25�$��@�d5�P�g��]	���������d�d�x�  P���� ��  8�� ҿ�!���D��$�M�_�qσϕϧ� ���������ƿv��F�X��/� ;�ob���pm��t�_�DiQ̡  � l�|�̡ĥ���� ���!�3�E�W�i�{� ������������� �/�A�S�e�]�Ӈ� ������������ );M_q��� ����r��� j�Tfx���� ���//,/>/P/ b/t/�/�/�/�/�/�%�/  0��6��!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O*�O�O �O�O__+_=_O_a_ s_�_�_�_�_�_�_�_ oo'o9oKo�O�OJ �o�o�o�o�o�o�o  2DVhz�� �����
�7?  ;�>�P�b�t��� ������Ǐُ���� !�3�E�W�i�{�������ß �ş3�ܟ ��&�8�J�\�n������������ɯ��v��,� ��+�	12345�678�� 	�
 =5���f�x�������������
� �.�@�R�d�vψϚ� ៾���������*� <�N�`�r߄߳Ϩߺ� ��������&�8�J� \�n�ߒ������� �����"�4�F�u�j� |��������������� 0_�Tfx� ������ I>Pbt��� ����!/(/:/ L/^/p/�/�/�/�/�/�/�2�/?�#/�9?K?]?�iCz � Bp˚   刅h2��*�$S�CR_GRP 1��(�U8(�\�xd�@� � ��'�	 �3�1�2�4(1 *�&�I3�F1OOXOn}m��D�@��0ʛ)���HUK�L�M-10iA 7890?�90;��F~;�M61C D�P:�CP��1
\&V�1	�6F��CW�9)A7Y	(R�_�_�_�_4�_�\���0i^ �oOUO>oPo#G�/ ���o'o�o�o�o�oB�0�rtrAA�0*  @蠈Bu&Xw?��ju�bH�0{UzAF@ F�`�r��o�� ���+��O�:�s� �mBqrr����������B�͏b����7�"� [�F�X���|�����ٟ ğ���N���AO�0�B�CU
L���E�jqBq�>7����$G@��@pϯ B����G�I
E�0EL_D�EFAULT  ��T���E��MIPOWERFL  
Ex*��7�WFDO�� *��1ERVE�NT 1����`(�� L!D?UM_EIP��>���j!AF_I�NE�¿C�!FIT������!o�:� ��a�!�RPC_MAIN�b�DȺPϭ�t�VI�S}�Cɻ����!�TP��PU�ϫ�d���E�!
PMON?_PROXYF߮�Ae4ߑ��_ߧ�f�����!RDM_S�RV�߫�g��)�!#R�Iﰴh�u�K!
v�M�ߨ�id����!RLSYN�C��>�8���!�ROS��4��4 ��Y�(�}���J�\��� ����������7�� ["4F�j|� ���!�Ei�o�ICE_KL �?%� (%SVCPRG1n >���3��3��"�4//�5./3/"�6V/[/�7~/�/���D�/�9�/�+ �@��/��#?�� K?��s?� /�?� H/�?�p/�?��/O ��/;O��/cO�? �O�9?�O�a?�O� �?_��?+_��?S_ �O{_�)O�_�QO �_�yO�_��Os� ���>o�o}1�o�o �o�o�o�o�o; M8q\���� �����7�"�[� F��j�������ُď ���!��E�0�W�{� f�����ß���ҟ� ��A�,�e�P���t���������ί�y_�DEV ���MC:���_!�OUT���2��REC 1q�`e�j� �	 �����˿��p�ڿ��
 �`e ���6�N�<�r�`ϖ� �Ϧ��Ϯ�������&� �J�8�n߀�bߤߒ� �߶�������"��2� X�F�|�j������� ��������.�T�B� x�Z�l����������� ��,P>`b t������ (L:\�d� ���� /�$/6/ /Z/H/~/l/�/�/�/ �/.��/?�/2? ?V? D?f?�?n?�?�?�?�? �?
O�?.O@O"OdORO �OvO�O�O�O�O�O�O __<_*_`_N_�_�_ x_�_�_�_�_�_oo 8oo,ono\o�o�o�o �o�o�o�o�o " 4jX����� �����B�$�f� T�v������������ ؏��>�,�b�P�r����p�V 1�}� �P
�ܟ�^�[J � 
��TYP�E\��HELL_?CFG �.��=͟  	�����RSR������ ӯ�������?�*� <�u�`���������Ῥ������%@�3�E��Q�\�Ұ1M�o�p��Ϸ��2Ұd]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&��1�OW_REG�_UI���IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he�#�� ��������Ҵ��) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������n���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( �}��>Pbt�� ,���� �;M_q��( ����//�7/ I/[/m//�/$/�/�/ �/�/�/?�/3?E?W? i?{?�? ?�?�?�?�? �?O�?/OAOSOeOwO �OO�O�O�O�O�O_ _�O=_O_a_s_�_�_ *_�_�_�_�_oo�_ 9oKo]ooo�o�o&o�o �o�o�o�o�o5G Yk}�"��� ����1�C�U�g� y��������ӏ��� 	���-�?�Q�c�u��� ��,���ϟ���� ��;�M�_�q�����(� ��˯ݯ�����7� I�[�m����$���ǿ ٿ���Ϣ�3�E�W��i�{ύ� �&cop�y mc:dio�cfgsv.io� md:=>in�spiron:3648������	���0��frs:or�derfil.d�at virt:?\temp\��`��r߄ߖ�)�(.�*.dB�T�W��������
xyzrate 61 ������n����%�.�O�H�Z������"�3.�@�mpbackN�b�t�܆��� }*��db��*C�U�Y�����6!�.x.�:\��8 @R���n��%�/.a6H_ ^� &�8�����m��� ����Z��/"4 �Xi/{/�/��C/ ��/�/?0BT e?w?�?��I?��?��?OO�$SNP�X_ASG 1�����9A�� P 0 �'%R[1]�@1.1O 9?�#3%dO�OsO�O�O�O �O�O�O __D_'_9_ z_]_�_�_�_�_�_�_ 
o�_o@o#odoGoYo �o}o�o�o�o�o�o�o *4`C�gy �������	� J�-�T���c������� ڏ�����4��)� j�M�t�����ğ���� ��ݟ�0��T�7�I� ��m��������ǯٯ ���$�P�3�t�W�i� �������ÿ���� :��D�p�Sϔ�wω� �ϭ��� ���$��� Z�=�dߐ�sߴߗߩ� ������ ��D�'�9� z�]��������� 
����@�#�d�G�Y� ��}������������� *4`C�gy ������	 J-T�c��� ���/�4//)/ j/M/t/�/�/�/�/�/��/�/?0?4,DPA�RAM �9E}CA �	��:�P�4�0$HOF�T_KB_CFG�  p3?E�4PI�N_SIM  9K�6�?�?�?�0,@�RVQSTP_DSB�>�21On8J0�SR ��;� G& =O{Op0�6�TOP_ON_E_RR  p4�9~�APTN �5��@A�BRING_PRM�O� J0VDT_G�RP 1�Y9�@  	�7n8_(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2Dkhz �������
� 1�.�@�R�d�v����� ����Џ�����*� <�N�`�r��������� ̟ޟ���&�8�J� \�����������ȯگ ����"�I�F�X�j� |�������Ŀֿ�� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�tߛߘߪ� ����������(�:� a�^�p������� ���� �'�$�6�H�Z� l�~���������������3VPRG_CO7UNT�6��A�5NENB�OM=��4J_UPD 1}��;8  
 p2������  )$6Hql~� ����/�/ / I/D/V/h/�/�/�/�/ �/�/�/�/!??.?@? i?d?v?�?�?�?�?�? �?�?OOAO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_��_�_YSDEBSUG" � �Pdk	��PSP_PASS�"B?�[LOG� ��mr�P�X�_  �g~�Q
MC:\d<�_b_MPCm�H�o�o�Qa�o �~vfSAV �m�:dUb�U\gS�V�\TEM_TI�ME 1�� �(�P�TNu]qT1SVGUNS} �#'k�spAS�K_OPTION�" �gospBC?CFG ��|� �b�{�}` ����a&��#�\�G� ��k�����ȏ����� �"��F�1�j�U��� y���ğ���ӟ��� 0��T�f��UR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz��rBr�|�|� ���z� �%��I� 4�m�X���|������� �֏���3��W�B� g���x�����՟���� ����S�>�w�b� ����'2A ��ʯܯ�� ����E�0�i�T��� x���ÿտ翢���� /��?�e�1�/���/ �ϜϮ��������,� �P�>�`߆�tߪߘ� �߼��������L� :�p�^������� ����� �6�H�>/`� r�������������� �� 0Vhz8 ������
 .�R@vd�� �����//</ */L/r/`/�/�/�/�/ �/�/�/�/?8?&?\? J?�?n?�?�?�?�?�� �?OO�?FO4OVOXO jO�O�O�O�O�O�O_ _�OB_0_f_T_v_�_ �_�_z_�_�_�_oo >o,oboPoroto�o�o �o�o�o�o(8 ^L�p���� ���$��H�6�l� ~�(O����f�d��؏ ���2� �B�D�V��� ����n����ԟ
��� .�@�R�d����v��� �����Я���*�� N�<�^�`�r�����̿ ���޿��$�J�8� n�\ϒπ϶Ϥ����� ��ߊ�(�:�L���|� jߌ߲ߠ��������� �0�B�T��x�f�� ������������,� �P�>�t�b������� ��������:( JL^����� � �6$ZH ~l��^���d� � //D/2/h/V/x/ �/�/�/�/�/�/�/? 
?@?.?d?v?�?�?T? �?�?�?�?�?OO<O *O`ONO�OrO�O�O�O �O�O_�O&__6_8_ J_�_n_�_�_�_�_�_ �_�_"ooFo��po �o,oZo�o�o�o�o �o0Tfx�H �������,� >��b�P���t����� ����Ώ��(��L� :�p�^�������ʟ�� �ܟ� �"�$�6�l� Z���~�����دꯔo ��&�ЯV�D�z�h� ������Կ¿��
�� .��R�@�v�dϚτ��  ���� ��������$TBJ�OP_GRP 2�ǌ�� � ?������������_xJBЌ���9� �< ��X���� @����	 �C��} t�b  C��<��>��͘Ր���>̚йѳ33�=�CLj�f�ff?��?�ff�BG��ь�����t��ކ�>�(�\�)�ߖ�E噙�;���hCYj�� � @h��B�  �A����f��C�  Dhъ�1���O�4�N����
:���Bl^���j�i�l�l����A�ə�A�"��D9��֊=qH����нp�h�Q�;�A�j��o��@L��D	2��������$�6�>B��\��T���Q�ts>x�@33@���C���y�1�����>��Dh�����x�����<{�h�@i� ��t ��	���K& �j�n|��� p�/�/:/k/������!��	V�3.00J�m61cI�*� IԿ���/�' Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I�!CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;��;Q�T,8�4`� *�ϴ?�2����3\�X/O��ESTPARS  ���	���HR@ABL/E 1����0�É
H�7 8��9
GB
H
H����
G	
HE

H
HYE��
H�
H
H6FRD	IAO�XOjO|O�O�O�ETO"_4[>_P_�b_t_�^:BS _�  �JGoYoko}o�o�o�o �o�o�o�o1C Ugy����`#o RL�y�_�_�_�_�O�O��O�O�OX:B�rNUoM  ���P��� V@P:B_CFG ˭��Z�h�@��IMEBF_TT%AU��2@��VERS�q���R 1���
 �(�/����b�  ����J�\���j�|��� ǟ��ȟ֟����� 0�B�T���x�������R2�_���@�
��MI_CHAN��� � ��DBGL�V���������E�THERAD ?U��O������h�����ROUT6�!��!����~��SNMASKD�|�U�255.���#�����OOLO_FS_DI%@�u�.�ORQCTRL �����}ϛ3r� �Ϲ���������%� 7�I�[�:���h�z߯��APE_DETA�I"�G�PON_S�VOFF=���P_?MON �֍��2��STRTCH/K �^������VTCOMPAT���O�����FPRO�G %^�%  BCKEDT-Q�<��9�PLAY&H��_INST_Mްe ������US��q��LCK���Q?UICKME�=�ރ�SCREZ�>G�tps� �� �u�z����_��@@�n�.�SR_GRP� 1�^� �O����
��+ O=sa�쀚 �
m������L/ C1gU�y �����	/�-/�/Q/?/a/�/	1?234567�0�/��/@Xt�1���
� �}ipnl�/� gen.htm�? ?2?D?V?`�Panel _setupZ<}P���?�?�?�?�?�?  �??,O>OPObOtO�O �?�O!O�O�O�O__ (_�O�O^_p_�_�_�_ �_/_]_S_ oo$o6o HoZo�_~o�_�o�o�o �o�o�oso�o2DV hz�1'�� �
��.��R��v����������ЏG���U�ALRM��G ?9� �1�#�5� f�Y���}�������џ�ן���,��P��S�EV  �����ECFG ���롽�A�� :��Ƚ�
 Q��� ^����	��-�?�Q��c�u�����������Ԇ� �����I2��?���(%D�6�  �$�]�Hρ�lϥϐ� �ϴ�������#��Gߌ��� �߿U�I�_Y�HIST 1}��  (��� ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1����(�:�� ����936�߆����K� ������	��-�?��� c�u���������L��� ��);��_q �����Z� %7I�m������f��f //'/9/K/]/`�/ �/�/�/�/�/j/�/? #?5?G?Y?�/�/�?�? �?�?�?�?x?OO1O COUOgO�?�O�O�O�O �O�OtO�O_-_?_Q_ c_u__�_�_�_�_�_ �_��)o;oMo_oqo �o�_�o�o�o�o�o �o%7I[m�  ������� 3�E�W�i�{������ ÏՏ�������A� S�e�w�����*���џ �����ooO�a� s���������ͯ߯� ��'���K�]�o��� ������F�ۿ���� #�5�ĿY�k�}Ϗϡ� ��B���������1� C���g�yߋߝ߯��� P�����	��-�?�*� <�u��������� ����)�;�M����� ������������l� %7I[��� ����hz! 3EWi���� ���v////A/�S/e/P���$UI�_PANEDAT�A 1������!  	�}w/�/�/�/�/?? )?>?��/ i?{?�?�?�?�?*?�? �?OOOAO(OeOLO �O�O�O�O�O�O�O�O\_&Y� b�>R Q?V_h_z_�_�_�__ �_G?�_
oo.o@oRo do�_�ooo�o�o�o�o �o�o*<#`G ��}�-\�v�# �_��!�3�E�W�� {��_����ÏՏ��� `��/��S�:�w��� p�����џ������ +��O�a������� ��ͯ߯�D����9� K�]�o��������ɿ ���Կ�#�
�G�.� k�}�dϡψ����Ͼ� ��n���1�C�U�g�y� ���ϯ���4�����	� �-�?��c�J��� ������������� ;�M�4�q�X����� ������%7�� [������� @��3Wi P�t����� /�//A/����w/�/ �/�/�/�/$/�/h? +?=?O?a?s?�?�/�? �?�?�?�?O�?'OO KO]ODO�OhO�O�O�O �ON/`/_#_5_G_Y_ k_�O�_�_?�_�_�_ �_oo�_Co*ogoyo `o�o�o�o�o�o�o�o -Q8u�O�O}��������)�>��U-�j�|� ������ď+��Ϗ� ��B�)�f�M����� ���������ݟ�&��S�K�$UI_P�ANELINK �1�U � �  ���}1234567890s������� ��ͯդ�Rq����!� 3�E�W��{�������ÿտm�m�&����Qo�  �0�B�T� f�x��v�&ϲ����� ����ߤ�0�B�T�f� xߊ�"ߘ��������� �߲�>�P�b�t�� ��0���������� ��$�L�^�p�����,� >������� $�0,&�[gI�m ������� >P3t�i�� Ϻ� -n��'/9/ K/]/o/�/t�/�/�/ �/�/�/?�/)?;?M? _?q?�?�UQ�=�2 "��?�?�?OO%O7O ��OOaOsO�O�O�O�O JO�O�O__'_9_�O ]_o_�_�_�_�_F_�_ �_�_o#o5oGo�_ko }o�o�o�o�oTo�o�o 1C�ogy� ����B�	�� -��Q�c�F�����|� ������֏�)�� M���=�?��?/ȟ ڟ����"�?F�X� j�|�����/�į֯� ����0��?�?�?x� ��������ҿY��� �,�>�P�b��Ϙ� �ϼ�����o���(� :�L�^��ςߔߦ߸� ������}��$�6�H� Z�l��ߐ������� ��y�� �2�D�V�h� z����-��������� 
��.RdG� �}����c� ��<��`r��� �����//&/8/ J/�n/�/�/�/�/�/ 7�I�[�	�"?4?F?X? j?|?��?�?�?�?�? �?�?O0OBOTOfOxO �OO�O�O�O�O�O_ �O,_>_P_b_t_�__ �_�_�_�_�_oo�_ :oLo^opo�o�o#o�o �o�o�o ��6H �l~a���� ����2��V�h� K�������1�U 
��.�@�R�d�W/�� ������П������ *�<�N�`�r��/�/? ��̯ޯ���&��� J�\�n�������3�ȿ ڿ����"ϱ�F�X� j�|ώϠϲ�A����� ����0߿�T�f�x� �ߜ߮�=�������� �,�>���b�t��� ���+������ :�L�/�p���e����� ������ ��6��🯡�ۏ��$UI�_QUICKME�N  ����}��RESTORE 1٩��  ��
�8m 3\n���G� ���/�4/F/X/ j/|/'�/�/�//�/ �/??0?�/T?f?x? �?�?�?Q?�?�?�?O O�/'O9OKO�?�O�O �O�O�OqO�O__(_ :_�O^_p_�_�_�_QO [_�_�_I_�_$o6oHo Zoloo�o�o�o�o�o {o�o 2D�_Q cu�o����� ��.�@�R�d�v���������Џ⏜SC�RE� ?��u1sc� uU2�3�4�5��6�7�8��UGSER����T����ks'���4��5*��6��7��8��� �NDO_CFG �ڱ  �  �� PDATE �h��Non�e�SEUFRA_ME  ϖ���RTOL_AB�RT����ENB�(��GRP 1���	�Cz  A�~�|�%|��������į֦��X�� U�H�X�7�MSK  �K�S�7�N�%�uT�%�����VI�SCAND_MA�XI�I�3���FAIL_IMGI��z �% #S���IM�REGNUMI�
����SIZI�� ��ϔ,�ONT�MOU'�K�Ε��&����a���a��s�F�R:\�� � �MC:\(�\wLOGh�B@Ԕ !{��Ϡ������z MCV�����UD1 �E�X	�z ��PO�64_�Q���n6��PO!�LI��Oڞ�e�V�N��f@`�I�� =	�_�SZVmޘ���`�WAImߠ�ST�AT �k�% @��4�F�T�$#�x� �2DWP  ���P G��=���͎���_�JMPERR 1�ޱ
  �p23�45678901 ���	�:�-�?�]� c���������������x��$�MLOW��8������_TI/�˘�'��MPHASOE  k�ԓ� ���SHIFT%�15 Ǚ��<z� �_����F /|Se��� ����0///?/ x/O/a/�/�/�/�/�/�����k�	VSwFT1\�	V���M+3 �5�Ք �p����A�  BU8[0[0�Πpg3�a1Y2�_3Y�7ME���K�͗	6e���&+%��M���b���	��$��TDI�NEND3�4��4O H�+�G1�OS2OI�V I���]LRELEvI��4.�@��1?_ACTIV�IT�<�B��A �m��/_��BRDBГOZ�YBOX �ǝ�f_\��b�2�T�I190.0m.�P83p\�V�254p^�Ԓ	� �S�_�[b��robot84�q_   px�9o\�pc�P ZoMh�]Hm�_Jk@1�o^�ZABCd��k�,���P\�Xo}�o0 );M�q�� ������>��a	Z�b��_V