��   I�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��ETH_FLT�R.� $� �  �FT�P_CTRL.� @ $LOG�_8	�CMO>�$DNLD_FI�LTE� � SUB�DIRCAP�!�(�HO��NT�. 4� H_NAME !ADDRTYP�A H_LENGT1H' �z +�LS D $ROBOTIG �PEER^� MwASKMRU~�OMGDEV#�� RDM*�D_ISABL&�OTCPIG/ 3 �$ARPSIZ�&_IPF'W�_MC��F_I�N� FA~LAS�Ss�HO_� I�NFO��TEL�K PV��b	 WORD  �$ACCES�S_LVL?TI�MEOUTuOR�T � �ICEU�S=   ��$#  �����!�� � � VIRTUAL�/�!'|0 �%
���F�����$�%����+ ������$�� �-2�%;�SHARED� 1�)  CP!�!�?���!|? �?�?�?�?O�?%O�? 1OOZOOBO�OfO�O �O�O�O_�O�OE__ i_,_�_P_�_t_�_�_ �_o�_/o�_SooLo �oxo�opo�o�o�o�o �o*Os6� Z�~����� 9��]� ���D�V��� z�ۏ����#����Y�H�}�@���)7z _LIST 1=_x!1.ܒ0���d�ە1�d�25c5.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I���� o�������O�6����8������ �$ ���-� ���-� ��&�%��&!Ò�)��0H!� ����rj3_tpd����! � �!!KC� e�0ٙ��&W�!Cm ��w߉�~S�!CON� ���1�=�smon��W�