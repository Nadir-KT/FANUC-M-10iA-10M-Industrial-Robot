��   I�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETGRO��ETH_FLT�R.  $��   ��FTP_CTRL�. @ $L�OG_8	�CMO�>$DNLD_�FILTE� � S�UBDIRCAP�����HO��NT�. 4� H_NAME !ADDRTYP�A H_LENGT1H'�z +�LS D $ROBOTIG �PEER^� MwASKMRU~;OMGDEV#��RDM*�DI�SABL&.S?V�TCPIG/ �3 $ARPS�IZ&_IPF�'W_MC��F�_IN� FA~L�ASSs�HO_ބ INFO��T;ELK PV��b	 WORD�  $ACCESS_LVL?TIMEOUTu�ORT � �ICgEUS= ��$#  ����!��� � � VIRTUAL�/�!'0 �%_
���F��e���$�%��;�+ ����#�$�� �-2%;��SHARED 1��)  P!�!�?���!|?�?�? �?�?O�?%O�?1OO ZOOBO�OfO�O�O�O �O_�O�OE__i_,_ �_P_�_t_�_�_�_o �_/o�_SooLo�oxo �opo�o�o�o�o�o *Os6�Z� ~�����9�� ]� ���D�V���z�ۏ ����#���Y�H��}�@���)7z _LI�ST 1=x!1.ܒ0��d�ە�1�d�255.�$������%ړ2 ��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I����o�������O�6���8��0���� �$�� �-� ���-��%�%���&!Ò�)�0H�!� ���r?j3_tpd���!� � �!!KC�� e�0ٙ��&W�!�Cm ��w߉�S�!CON� ��1�==�smon��W�