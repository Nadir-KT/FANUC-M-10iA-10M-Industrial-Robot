��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �ET�H_FLTR.�� $�  � �FTP_C�TRL. @ ?$LOG_8	��CMO>$DN�LD_FILTE�� � SUBDIR�CAP�� HOv��NT. 4� �H_NAME �!ADDRT�YPA H_LE�NGTH' ��z +LS �D $ROBO�TIG PEER�^� MASKM�RU~OMGDEuV#� RDM*��DISABL�&1� TCPI�G/ 3 $AR�PSIZ&_I{PF'W_MC�ދF_IN� FA�~LASSs�H{O_� INFO���TELK P�V�b	 WO�RD  $A�CCESS_LV�L?TIMEOU=TuORT � ��ICEUS=  �1 �$#  ����!�� � � VIRTUAL�/�!'0 �%
U���F�����$��%���+3 �����$�� ��-2%;�SHAR�ED 1�)  P!�!�?���!|?�?�?�?�?O�? %O�?1OOZOOBO�O fO�O�O�O�O_�O�O E__i_,_�_P_�_t_ �_�_�_o�_/o�_So oLo�oxo�opo�o�o �o�o�o*Os 6�Z�~��� ��9��]� ���D� V���z�ۏ����#� ��Y�H�}�@���)7�z _LIST 1}=x!1.ܒ�0��d�ە�	�f��255.$����	��%ړ2��X���+�=�O�3Y��Р �������O�4ѯ�@H���	��-�O�5I�����o�������O�6 ���8������ �$���-� ����-� �&�%��&!Ò:�)�0H!� ����rj3_t�pd���! � �!!KC� e�0ٙ�<�&W�!Cm ���w߉�S�!CO�N� ��1�=�smon��W�