��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ��'�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"�SBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�� W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2F�G1_�3�B�2��XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�0@� �zsa�!ip;G0� � 
$WARNM�0f�!,P� ܁s�pNST� CO�RN�"a1FLTR^�uTRAT� T�p; H0ACCa1�p��{�ORI
`l"S={RT0_S�BְqHG,I1 E[ Tp�"3I9�CTY�D,P*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7���8��94�G CO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0����p� �v�p��PzPb26����"J��_R��BC�J��3�JVP��tB�S��}Aw��"�tP_�*0OFSzR @�� RO_K8���aIyT�3��NOM_�0��1ĥ3W ��TC �� $���AxP��K}EX�� �0g0I0x1��p�
$TFa�ކC$MD3��TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF�vF���Pp@�a2 6
P$A`PU�3N�)#�dR*�AqX�!sDETAI�3�BUFV��p@1c |�p۶�pPIdT�� PP[�MZ�M�g�Ͱj�F[�SIMQSI�"0��A.�����kx Tp|zM��P�B�FACTrbHPEW7�P1Ӡؖ�v��MCd�5 �$*1JB�p<�*1DECHښ�H��ľb� � +PN�S_EMP��$GP���,P_��3�p2�@Pܤ��TC��|r ��0�s��b�0�� �B0���!
���JR� ��_SEGFR��Iv *�aR�TkpN&S,��PVF4��� &k�Bv�u�cu� �aE�� !2��+�MQ��E�SIZ�3�����T��P�����aRSINF�����kq�� ������LX������F�CRCMu�3CClpG��p���O}�� �b�1�������2�V�DxIC��C���r��`��P��{� EV ��zF_��F�pNB0�?������A�! �r�Rx�� ��V�lp�2��aR�t��,�g�RTx #�5�5"2��uA�R���`CX�$LG�p��B�1 `s�P�tB�aA�0{�У+0R���tME�`!BupCfrRA 3tAZ��h��pc�OT�FC�b�`�`FNp���1��ADI+�a%��b �{��p$�pSp�c�`aS�P��a,QMP6䒁`Y�3��M'�pUt��aU  $>�TITO1�S�S�!���$�"0�DBPX�WO��!��$3SK��FDB��"�"@�PR8� �
� ���# l>�q1$��$��
+�L9$?(�V�)%@?R4C&_?R4gENE��'~?�(�� RE�pY2(�H �OS��#$L�3$$3R�h�;3�MVOk_D@!V�ROScrr�w�S����CRIGGER�2FPA�S��7�ET�URN0B�cMR_���TUː[��0EkWM%���GN>`���RLA���Eݡ<�P�&$P�t�'�@4a��C�DϣV��DXQ��4�1��MVG�O_AWAYRM�O#�aw!�D�CS_)  `IS#� �� �s 3S�AQ汯 4Rx�@ZSW�AQ�p�@1UW��NcTNTV)�5RV
a����|c�éWƃ��J�B��x0��SAFE�ۥ�V_SV�bEX�CLUU�;��ONL��cYg�~az��OT�a{�HI_V�? ��R, M�_ �*�0� ��_z�2�� CdSGO  +�rƐm@�A�c~b���w@��V�i�b�fANNUNx0�$�dKIDY�UABc�@@Sp�i�a+ �j�f��!��pOGIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�� 6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6CqibMSW�U. 8��KEYI��5�TM�1�s�qoA�vINޱw��", �/ D��HOST�P!4���<���`<�°<��p<�EM'����Z�� SBL� U}L��0  �	���E�� T�01� � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0QSp�����#��SAV� ����c�S< 9�`�f�P$�0E!� YN�_B�#2 0��D�I�d�pO|�m��#�$F�R_IC� �ENC2_Sd3  ��< 3�9���� cgp����!4�"��2�A��ޖ5���`ǻ�@�Q@K&D-!�a�AV�ER�q����DSP
���PC_�q��"��|�ܣ�VALU�3�HE�(�M�I�P)���OPPm ��TH�*��SH" T�/�Fb�;�d��`��d ��Ш�ET�6 H(rLL_DUǀ�a�@��k���֠OT�"U�/���q@@NOAUT5O70�$}�x�~�@s��|�C͠���C� 2��z�L��� 8H *��L� ���Բ@sv� �`� �� ÿ���Xq��@cq���q���q��7���8��9��0���1��1 �1-�1:�1�G�1T�1a�1n�2R|�2��2 �2-�U2:�2G�2T�2a�U2n�3|�3�3˪ �3-�3:�3G�3*T�3a�3n�4|��q8���9 <���z�ΓKI����H硵�BaFEq@{@: y,��&a? PF_P?��>�����E�@��QQ��;�fp$TP�$�VARI����,�U�P2Q`< W�߃TD��g���`�������͠��BAC�"= T2����$)�,+r³�p IFI��p�� q M�P"�0��Fl@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� Fa@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(�q�#5T�DG���� �%�'�FSS� )�? P(q1�1�E`_1"811��EC13D;5D6��GRA���@��4���PW�ON2EBUG�S�2�C`�gϐ_E A ��o� �TE�RM�5B�5�O�ORIw�0C�5���SM_-`����0D�5&���TA�9E�5DG��UP��F� -QϒA�P�3�@�B$SEGGJ� E�L�UUSEPNFI��pBx��1@��4�>DC$UF�P��C$���Q�@C��ĳG�0T�����SNSTj�PATۡg��AOPTHJ�A�E*� Z%qB\`F�{E��F�q��pARxPY�aSHF�T͢qA�AX_SH�OR$�>��6 @$�GqPE���OVRH���aZPI@P@$U?r= *aAYLO���j�I�"��Aؠ��ؠERV��Qi�[Y)� �G�@R��i�e��i��R�!P�uASYM���uqAWJ�G)��AE��Q7i�RD�U[d@�@i�U��C�%UP��X�P���WOR�@M��k0SMT��GƇ�GR��3�aPA�@��p5�'�H �� j�A�TOC�jA7pP]Pp$O�Pd�O��C�%�p��O!��RE.pRĈC�AO�?��Be�5pR�EruIx'QG�eo$PWR) IMdu��RR_$s��5��B �Iz2H8�=�_A�DDRH�H_LE�NG�B�q�q:�x�Rj��So�J.�SS��SK������ ��F-�SE*���rSN�[MN1K	�j�05�@r�֣OL��\��WpW�Q�>pACRO �p���@H ����Q�� ��OUPW3�b_">�I��!q�a1���� ����|���������-���:���iIO
X2S=�D�e��]���L $��p�!�_OFF[r_�PR�M_�̱HTT�P_�H��M (��pOBJ�"�pG�-$H�LE�C��ٰ�N � 9�*�AKB_�T��
�S�`l�S��LV��KRW"~duHITCOU?[BGi�LO�q�����d� Fpk�GpS9S� ���HWh�wA��O.��`INC�PUX2VISIO ��!��¢.�á<�á~-� �IOLN)�P 87�R'�[p�$SL�bd PU�T_��$dp�P�z �� F_AS:2Q/�$LD����D�aQT U�0]P�A0������PHYG灱�Z���5�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp��㱰x��ٶ��UJ��S����NE�WJOG��G �DIS��&�K�Ġ��3T |��AV8��`_�CTR!S^��FLAGf2&�LG�dU �n�:��3?LG_SIZ��`�ň��=���FD��I����Z �ǳ��0�� ��@s��-ֈ�-�=�-����-��0-�ISCH�_��Dq��N?���V
��EE!2�C��"n�U�����`L�Ӕ�7DAU��EA��Ġt����GHr��I��BOO)�WL ?`�� ITV���0�\�REC�SCR�f 0�a�D^�����MARG��`!P�)�T��/ty�?I�S�H�WpW�I���T�JGM���MNCH��I�FN�KEY��K��PR�G��UF��P��F�WD��HL�STP��V��@�����RSS�H�` �Q�C��T1�ZbT�R ���U �����|R��t�i���G��8PPO��6�F�z1�M��FOCU���RGEXP�TUI��IЈ�c��n ��n����ePf���!p�6�eP7�N���CAN�AI�jB��VAIL杆CLt!;eDCS�_HI�4�.��O��|!�S S�n瘱I�BUFF�1XY��PT�$�� �v��f���װA�rYY��P ���\��pOS1�2��3�K�0Z �  ��aiE�*���IDX�dP�RhrO��+��A&ST��R���Yz�<! Y$EK&CK+���Z&pm&�F�1[ L�� o�0��]PL�6pwq�t�^����w��7�_ \ �`��瀰�7�t�#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3�1DM�R7��LDR5<4R5ORG.���e2(` ���V�8.��T<�4�d^ �q�<4��-4R5�S�`T00m��0D>FRCLMC!D�?0�?3I@��MIC��dg_ d���RQm�=q�DSTB	� c �Fg�HAX;b� �H�LEXCE�SZr�oEMup�a`Z��B;d�rB`��`5a��F_A�J���$[�O�H0K�db q\��ӂS�$MB���LIБ}SREQU�IR�R>q�\Á�XD�EBU��oAL� MP�c�ba��P؃ӂ!B�oAND���`�`d0�҆�c�cDC1��IN�����`@�(h?�Nz�@q��o� ��SPST8� en�rLOC�RI�p�EX�fA�p��A�oAODAQP�f �X��ON��[rMF �����f)�"I��%�e؃�T��FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y��RFЭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?
�uD�)�b�	@Ð�i �@CU��V��T0�eRR2�j� Dɐ�Qނ�Bd$OCALI�@F�G�:s�2�RIN��v��<NV�INTE���kE���,��b����_Nl��ڂ���kDׄRm�DIVFiFDH�@ـn��$V��'c!$��$Z������~�[��oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS�@#2L  �Ė83ಀ����� ��PAT!H��������3̒Vp�A_�Q�.�4�B��Cᐈ�_MGh��$DDQ���G�$FWh��p��m������b�DE��PPAB�NԗROTSPE!ED����00J�Я�8��@��̐$US�E_��P��s�S�Y��c�A kqYNru@Ag��OFF�qn�MOUN�NGg��K�OL�H�INC *��a��q��Bj�L@�BENCS��q�BđX���D��IN#"I̒0��4�\BݠVEO�w�>Ͳ23_UPE�߳/LOWL���00����D���BwP���� �1RCʀƶMO3SIV�JRMO���@�GPERCH  �OV��^��i� <!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸUPp������TRKr�>"AYLOA'a��  Q-�̒<�1Ӣ`0 ���RTI$Qx�0 MO ���МB R�0J��D���s�H����b�DU�M2(�S_BCKLSH_C̒��>� =�q�#�U��ԑ���2�<t�]ACLALvŲp�1n�P�CHK00:'%SD�RTY4�k���y�1�q_6#2�_�UM$Pj�Cw�_�S�CL��ƠLMT_OJ1_LO��@���q��E�����๕�幘SPC��7���L���PCo���H� ȰPU�m�C/@�"XT\_�c�CN_��N��Le���SFu���V��&#����9�̒��=�C�u�SH6#��c��� �1�Ѩ�o�0�͑
��f_�PAt�h�_Ps�W�_10��4�R�01D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�sR0Hљ��_W��-ԁ_=��C��I��I*�I�II�F�`�aJLA.�1[�VC��0�D�BO1U�@i�B\JRKU��~	@DBL_SMd�:BM%`_DLC�BGRV��C��I���H_� �*CcOS+\�(LN� 7+X>$C�9)I�9)u*c,)�Z2 HƺcMY@!�( "TH&-��)THET0�N�K23I��"=�A C-B6CB=�C�A�B�(261C�616SB8C�T25GTS QơC��aS$" �4c#<�7r#$DUD�EX��1s�t��B�6���AQ�|r�f$NE�DpI B U�\B5��$!��!�A�%E(G%(!LCPH$U�2׵�2SX pCc%pCr%�2�&�C�J�&!�VAHV6H3�YLUVhJVuKV�KV�KUV�KV�KV�IHAH@ZF`RXM��wXuKH�KUH�KH�KH�KH�I�O2LOAHO�YWNO�hJOuKO�KO�KO*�KO�KO�&F�2#1�ic%�d4GSPBA?LANCE_�!�c�LEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%�Ċ1ky�UTO_<?�jT1T2Cy��2N&�v�ϰctw�gѠp�0Ӓ~���T��O����� INSEGv�!�REV�v!���gDIF��1l�w6�1m�0OB�q
����MIϰ1��L�CHWAR����A�B&u�$MEC�H,1� :�@�U�AX�:�P��Y�G$�8pn� 
Z��|���RO�BR�CR̒��N�'�MSK_�`�f�p P Np_���R����΄ݡ�1 ��ҰТ΀ϳ��΀"��IN�q�MTC�OM_C@j�q � L��p��$ONORE³5����$�r 8� GRl�E�SD�0ABF��$XYZ_DAx5A���DEBU�qXI��Q�s �`$�wCOD�� ���k�F�f�$BU�FINDXР��
��MOR��t $-�U��)��rРB��Ӱ��Gؒu� � $SIMULT ��~�� ����OBJE�` �AD�JUS>�1�AY_	Ik��D_����C��_FIF�=�T � ��Ұ��{��p� ��З��p�@��D�FRiI��ӥT��RO� �E��S�OPsWO�ŀv0���SYSBU�@ʐ$�SOP����#�U<"��pPRUN�I�PA�DH�D����_OU�=��qn�{$}�IMAG��iˀ�0P�qIM��Ơ�IN�q���RGOVRDȡ:���|�aP~���Р�0L_6p0���i��RB���0e��M���EDѐ*F� ��N`M*�������˱SL�`ŀw� x $OVS�L�vSDI��DEXm�g�e�9w�����	V� ~�N���w���ІÛǖȳ�M�����q<��� x �HˁE�F�ATUS
���C�0àǒ�çBTM����If�¿�4����(�ŀy �DˀEz�g���PE��r�����
���EXE��V��E�Y�$Ժ �ŀz @ˁ��UP�{�h�$�p��XN����9�H� ��PG"�{ h �$SUB��c��p_���01\�MPWAI2��P����LO��<��F�p�$RCV?FAIL_C�f��BWD"�F���DE�FSPup | Lˀ`�D�� U�UNI��S���RX`���_L�pP��%�P�ā}��� @B�~���|��`�N�`�KET��y���Pԙ $�~���0SI�ZE��ଠ{���S�<�OR��FORMAT/p � F���r�EMR��y�UX����LI7�ā�  $�P_�SWI�M��_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W ��U����� A$PI�6 ���	��)�4�l�}69��Q�����S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�aO�0\H��6@�R�� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�H�t��W�UpS���R�M��O㵐.'}q��C�g���@ʣ����S�M��AÂ� � $sPY��$WH`'�NGp���H`��Fb`��Fb��Fb��PLM�@��	� 0h�H�{�X��	O��z�Z�eT�M���G� pS��C���O__0_B_�a��_%�� |S����@	 �v��v �@���w�vr��EM��% ����dt�B�����ftPn��PM��QU� �U�Q��Af�wQTH=�HOL��oQHYS�ES�F,�UE��B��O#��  ��P0�|�gAPQ���ʠu���O��ŀ�ɂv�-�A;ӝGROG��a2D��E�Âv�_�ĀZ�INFO&��+����b�Ȝ�OI킍 ((@SLEQ/�#�����pO�o���DS`c0O�0�01�EZ0NUe�_�AUyT�Ab�COPY�P�Ѓ�{��@M��N������1�P�
� ��RiGI�����X_�P�l�$�����`�W��P��j@�G���EXT_CYCtb!���p����h�7_NA�!$�\��<�RO�`]�� � m��PORp�ㅣ���SRVt��)����DI �T_ l���Ѥ{�ۧ��ۧ Ъۧ5٩6٩7٩8�����S�B쐒���$�F6���PL8�A�A^�TAR��@ E `�Z�����<��d7� ,(@FLq`hѦ�@YNL���M�C���PWRЍ��=�e�DELAѰ�mY�pAD#q�w��QSKIP�� iĕ�x�O�`NT!���P_x���� �@�b�p1�1�1� ��?� �?��>��>��&�>�3�>�9�Js2R;쐖 4��EX� TQ����ށ +����[�KFд�w�wRDCIf� �U`
�X}�R�#%M!*��0�)��$RGEAR�_0IO�TJBFL1G�igpERa��T�C݃������2TH�2N��� 1��b��Gq T�0 I����M���`Ib�\�v�REF�1�� l�h��ENA9B��lcTPE?@�� ��!(ᭀ����Q�#��~�+2 H�W���2�Қ���"�4�F�X�
j�3�қ{����\���� ��4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:Lj�7�ҟo@�����j�8�����"4Fj�SMSK������a��E�A O���MOTE�������@ "1�+��I�O�5"%I��p��PsOWi@쐣  �@����X�gpi�쐤���Y"$DSB_SICGN4A�Qi�̰C��^>%S232%�Sb��iDEVICEU�S#�R*�PARI�T�!OPBIT��Q��OWCON�TR�+�ⱓ*�C�U� M�SUXTA�SK�3NB��0�$T�ATU�P�qRIS@@쐦F�6�_�P�C}�$FREEFROMS]p�ai��GETN@S�UPDrl�ARB��RSP%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG �G|�.2���F��1�!d�9Z�8+5K�+5�� �y�L0�4��X �0m�L
N�T�3Hz��89��%��4�3G��W�0�W�RdD�Z��Tܳ���K�a3d��$cV �2���1��I1TH�02K2sk3K3Jci�aI�i�a�0L��SL��R$Vؠ�B�V�EVk�]V*R��� �,6Lc���9V2�F{/P:B��PS_�E�t�$rr�C�ѳ3$A0��wPR���v�U�cSk�� {��8��G� 0���VX`�!�tX`��0P�Ё��
�5SK!� �"-qR��!0���z�MNJ AX�!h�A�@�LlA��A�THIC��1�������1TF�E���q>�IF_C	H�3A�I0�����G1�x������9��Ɇ_JF҇PR|(���RVAT�� �-p��7@�����DO�E��COU�(��AXIg��O�FFSE+�TRIG�SK��c���Ѽ�e��[�K�Hk���8�IG#MAo0�A-��ҙ��ORG_UNEV���� �S�쐮�d �$�������GROU��ݓTqO2��!ݓDSP���JOG'��#	�_P'�2OR���>P67KEPl�IR�0�2PM�RQ�AP�Q���E�0q�e���SYS�G��"��PG��BRAK*Rd�r�3�-���0����ߒ<pAD��ݓ�J�BSOC� N��DUMMY14��p\@SV�PDE_�OP3SFSPD�_OVR��ٰC�O��"�OR-��Nı0.�Fr�.��OV��SFc�2�f��F���!4�S��RA�"L�CHDL�REC�OV��0�W�@M�յ�RO3��9_�0� @�ҹ@�VERE�$OF�S�@CV� 0BWD�G�ѴC��2j�
�T�R�!��E_F�DOj�MB_CM4��U�B �BL=r0�w�=q�tVfQ��x0spd��_�Gxǋ�AM��`k�J0������_M���2{�#�8$CA��{Й���8$HB�K|1c��IO��8.�:!aPPA"�N��3�^�F���:"�DVC_DB�C��d�w"����!��1���ç�y3����ATIO� �q0�UC�&CAB�BS�PⳐ�P�Ȗ��_0c�S�UBCPUq��S �Pa aá�}0�Sb��c���r"ơ$HW_AC���:c��IcA�A~-�l$UNIT��l��ATN�f�����CYCLųNEC�A��[�FLTR_2_FI���(��}&Ɩ�LP&�����_S[CT@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb��r�: _T��PROX��O�� EM�_�r��8u�q u��q��DI�0e�RAOILAC��}RMƐCLOԠdC��:anq���wq����PR��S�LQ�pfC��30	���FUNCŢ�rRINkP+a�0 ��!3RA� >R 
Я8�ԯWAR�#BLFQ��A�����DA�����LDm0�aB9�2�nqBTIvrb8ؑ���PRIAQ1�"AFS�P�!���𰠓�`%b���M�I1U�DF_j@��y1�°LME�FA�@H�RDY�4��Pn@R�S@Q�0"�MUL�SEj@f�b�q ��X��ȑ���m$.A$�1$c1�Ó���� x~�EG� ݓ�q!cAR����09>B��%��AXE��RKOB��W�A4�_�-�֣SY���!6��&S&�'WR���-1����STR��5�9�E�� 	5B��=Q�B90�@6������O�T�0o 	$�A�RY8�w20���	�%�FI��;�$LGINK�H��1�aI_63�5�q�2XYZ"��;�q�3@�R�1�2�8{0B�{D��� CFI��6G��
�{��_J��6��3aO�P_O4Y;5�QT�BmA"�BC
�z�D�U"�66CTURN3�vr�E�1�9���GFL�`���~ �@��5<:7�� 1��?0K�Mc�68�Cb�vrb�4�ORQ ��X�>8�#op�������wq�Uf�����TOVE�Q��M;�E# �UK#�UQ"�VW�ZQ �W���Tυ� ;��� �QH�!`�ҽ��U�Q�W`keK#kecXER�
�	GE	0��S�dAWaǢ:D���7!�!AX�rB!{q ��1uy-!y�p z�@z�@z6Pz\P z� z1v�y� y�+y�;y�Ky� [y�ky�{y��y�qޜyDEBU��$ ����L�!º2WG` � AB!�,��SV���� 
w���m� ��w����1���1���A ���A��6Q��\Q���!��m@��2CLAB�3B�U�����S 7 ÐER����� � $�@� A6ؑ!p�PO���Z�q0w�^�_MRA�ȑ� d  T�-�ERR��ÏSTYz�B�I�V3@��cΑTOQ�d:`L�� �d2�]�X�C�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	�SFZN�_CFG_!� 4 ��?º�|�ų����@�ȲW �]���\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(����$�!s�Q�g�P{RV �HELLĥ�� 56�B_BAS�!�RSR��ԣo ��#S��[��1r�%���2ݺ3ݺ4ݺ5*ݺ6ݺ7ݺ8ݷ���ROOI䰝0�0NLK!�CAB� ���ACK��IN��T�:�1�@�@ z�m�_�PU!�CO� ��OU��P� Ҧ) ��޶���TPFWD_�KARӑ��RE�~��P��(��QU�E�����P
��CSTOPI_AL������0&���㰑�0S#EMl�b�|�M��dЛTY|�SOK�}�D�I�����(���_�TM\�MANRQ�ֿ0E+�|�$K�EYSWITCH�&	���HE
�B�EAT����E� LQEҒ���U��FO������O_HOM��O�REF�PPARz��!&0��C+�9OA�ECO��B<�rIOCM�D8׆��]���8�` �# D�1����U��&��MH�»P�CFOR�C��� ���O}M�  � @V�T�|�U,3P� 1-��`� 3-�4���N�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��C@�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fim7s�'��VP��UPD��  ���|�԰��YSL}OǢ� � z� �и���o�E��`>�^t��АALUץ�����CU���wFOqID�_L�ӿuHI�zI~�$FILE_����t��$`�JvSAΒ�� h���E_BLCK�#�C,�D_CPU<�{�<��o����tJr��Rw ��
PW �O� ��LA��Sp��������RUNF� Ɂ��Ɂ����F�ꁡ�|ꁬ� �TBCu��C� �X -$�LENi��v�������I��G�LO�W_AXI�F1��t2X�M����D�4
 ��I�� ��}�GTOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑTCV����T���&��ݡ����HJ�����J����Mo�"��J�Ǜ �������2��� v�����6F�JK��VKi�Ρ4v�Ρ3��J0�ң�JJڣJJ�AAALң�ڣ��4�5z�&�N1-�9����␅�L~�_Vj�{x+p���� ` ��GROU�pD��B>�NFLIC��REQUIREa�EBUA��p����2¯�����c��� \��APP�R��C���
�E�N�CLOe��SC_M v�,ɣ�
�ޣ�� ���MCp�&���g�_MG�q�C� �{�9���|�wBRKz�NOL��t|ĉ R��_LI|�H�Ǫ�k�J����P
� ��ڣ�����&���/�"��6��6��8���|���� ���8�%�W�2�e�PATHa�z�p�z�=�vӴ��ϰ�x�CN=�CaA�����p�IN��UC��bq��CO�U�M��YZ������qE�%���2������PA�YLOA��J2L�3pR_AN��<�L���F�B�6�R�{�R_?F2LSHR��|�LOG��р��ӎ���ACRL_u��������.���H�p�$yH{���FLEX
��s�J�� :�/����6�2���0��;�M�_�F16�� ��n���������ȟ��Eҟ�����,�>� P�b���d�{�����@�������5�T��X��v���Eť mFѯ��������&�/�A�S�e�D�J>x�� � ������j�4pAT����n��EL  �%øJڪ��ʰJE��CTYR�Ѭ�TN��F&���HAND_VB�[
�pK�� $�F2{�6� �rS�Wi�yr�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�(#�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������uN���2�H̟�����"CqENL� a�DI��>�Obt8C�Dpx�� ��2IxQA����q��-���s �� ����� ���OMME���rr/�TVpPT@�P ���qe�i�����P�x ��yT�Pj�� $DUMMY}9�$PS_��RFq�  ��:�� ���!~q� �X����K�STs��ʰSBR��M21�_Vt�8$SV_�ERt�O��z���C+LRx�A  O�r?p�? Oր � D $GLOB���#LO��Յ$�o���P�!SYSA�DR�!?p�pTCH>M0 � ,��ސ�W_NA���/�e�$%SR��l (:]8:m� K6�^2m�i7m�w9m� �9���ǳ��ǳ���ŕ ߝ�9ŕ���i�L� ��m��_�_�_�TDџXSCRE�ƀӚ� ��STF���1}�pТ6��D�] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��tC�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$��VSHIF��|s�P�p�6��s���R���OSU�RW�pRADIz��2�_�q�h�g!� �q)�LUza�$OUTPUT_3BM��IML�oRp6(`)�@TIL<'SCO�@Ce�; ��9��F��T��a ��o�>�3�����w�2u�sqV�zu✫�%�DJU��|#_�WAIT������%ONE���YBOư ��� $@p%�C�S�Bn)TPE��NE�C��x"�$t$���*B_T��R��%�qRH� ���sB�%�tM�+ ��t�.�F�R!݀���OPm�MAS�_�DOG�OaT	�D�����C3S�	�O2DE�LAY���e2JO ��n8E��Ss4'#J�aP`6%�����Y_��O2$��2���5��`?� n=pZAB�CS��  $��2��J�
sp�$$�CLAS������AB�sp'@@V�IRT��O.@AB�S�$�1 <E�� < *AtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v�����M@[�AXLրK�*B��dC  ���IN8��ā��PRE������LARM�RECOV �<I䂥�NG�� �\K	 =#�
�J�\�M@PPLIC��?<E�E��HandlingTool ��� 
V7.50�P/28 *A�(�m��
�_S�W�� UP*A�� ��F0ڑ����A�G@�� 20���*A���:�����xFB �7DA5�� ~'@)m@�𞝓None������� ��T���*A4lx��P_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ�:�i�n�����#BGB ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��e��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���oe�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� ��PB�Z?����5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`ϖ�S:�(����Yp0�_)o�S`�BBia�P�_mo8j�(�aKoo�o9i�(�E�og�o�o�m�o�f�oGq:I�ZDE�F f8��)��R6pbuf.txAtm�]n�@�����# 	`(Ж�A=L����zMC�21B�=��9���4�=��n׾�Cz  B�HBCCPUeB���CF�;.�<C���C�5rSZE@D�ny�DQ��D���>��D�;�D����F���>F�$G}�RB�Gz&ր��SY��!�vqG����Em�(�.*��(�(��<�qѦG�x2��Ң �L� a�D�j���E�e���EX�EQ��EJP F�E��F� G��ǎ^F E��� FB� H,-� Ge��H3Y����  >�3�3 ���xV � n2xQ@��5Y���8B� A�AST<#�
� �_'�%�~�wRSMOFS����~2�yT1�0DOE �O c
�v(�;�"�  <�6�z�R���?�j�KC4��SZm� W�Q�{�m�C��B-JG�C�`@$�q���T{�FPROG C%i����c�I���� �Ɯ�f�KEY_�TBL  �vM��u� �	
��� !"#$%&�'()*+,-.�/01c�:;<=�>?@ABC�pG�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������p���͓���������������������������������耇����������������������!j�LC�K��.�j���STA�T���_AUTO�_DO���W/�INDT_ENB�b�2R��9�+�T2wߞXSTOP\߿2T{RLl�LETE�����_SCREE�N ik�csc��U��MM�ENU 1 i  <g\��L� SU+�U��p3g���� ���������2�	�� A�z�Q�c��������� ������.d; M�q����� �N%7]� m���/�� /J/!/3/�/W/i/�/ �/�/�/�/�/�/4?? ?j?A?S?y?�?�?�? �?�?�?O�?O-OfO =OOO�OsO�O�O�O�O��O_�O_P_Sy�_?MANUAL��n��DBCOU�RIG|���DBNUM�p���<���
�QPXWORK 1!R�ү�_oO.o@oRk��Q_AWAY�S^��GCP ��=��df_AL�P�db�R�Y�������X_�p �1"�� , 
��^���o xvf`M�T�I^�rl@�:sOoNTIM�������Zv�i
õ�cM?OTNEND���d�RECORD 1�(R�a��ua�O��q��sb�.�@� R��xZ�������ɏ ۏ폄���#���G��� k�}�����<�ş4�� X���1�C���g�֟ ��������ӯ�T�	� x�-���Q�c�u����� �����>����)� ��Mϼ�F�࿕ϧϹ� ��:�������%�s`Pn &�]�o��ϓ�~ߌ��� 8�J�����5� �� k����ߡ��J����� X��|��C�U���� ������0�����	���dbTOLERE�NCqdBȺb`L��͐PCS_CF�G )�k)wd�MC:\O L%04d.CSV
��Pc�)sA �CH� z�P)~����hMRC_OU/T *�[�`+~P SGN +�e��r��#�10-�MAY-20 0�9:27*V27-�JANj21:4�8�k P;����)~�`p�a�m��PJ�PѬVERS�ION S?V2.0.�6t�EFLOGIC {1,�[ 	DX��P7)�PF."PR?OG_ENB�o�r.j ULSew �T��"_WRSTJN�Ep�V�r`dEMO_�OPT_SL ?�	�es
 	R575)s7)�/?�?*?<?'�$TO � �-��?&V_V@pEX�Wd�u�3PATH AS�A\�?�?O/{IkCT�aFo`-�g�dseg�M%&ASTBF_TTS�x�Y^C��Sq:qF�PMAU� t/.XrMSWR.�i6Q.|S/�Z!D_ N�O0__T_C_x_g_��_�tSBL_FA�UL"0�[3wTD�IAU 16M6p��A1234?567890gFP?BoTofoxo�o �o�o�o�o�o�o@,>Pb�S�pP�_ ���_s��  0`�����)�;� M�_�q���������ˏpݏ��|)UMP�!f� �^�TR�B8�#+�=�PMEfEI��Y_TEMP9 Ç��3@�3A v�U�NI�.(YN_B�RK 2Y)E�MGDI_STA��%WЕNC2_S_CR 3��1o "�4�F�X�fv�����`����#��ޑ14� ���)�;�����ݤ5�����x� f	u�ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/߭ P�b�t�� ��xߞ߰� ��������
��.�@� R�d�v������� ������*�<�N��� r��������������� &8J\n� ������� "`�FXj|�� �����//0/ B/T/f/x/�/�/�/�/ �/�/�/4?,?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO �O�O�O�O�O?�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�O �O�o�o�o
.@ Rdv����� ����*�<�N�`� r����o����̏ޏ�� ��&�8�J�\�n��� ������ȟڟ�����H�ETMODE �16��� ��ƨ
R�d�v��נRROR_PR�OG %A�%��:߽�  ��TAB_LE  A�������#�L�RRSE�V_NUM  <��Q��K�S����_AUTO_ENB  ��I�Ϥw_NOh� 7A��{�R�  *�*�����������^��+��Ŀֿ迄�HI�SO�͡I�}�_AL�M 18A� �2;�����+�e�@wωϛϭϿ��_H�.��  A���|���4�TCP_VE/R !A�!�����$EXTLOG_7REQ��{�V��SIZ_�Q�TOL�  ͡Dz���=#׍�XT_BWD����r���n�w_DI�� 9���}�z�͡m���S�TEP����4��O/P_DO���Ѡ�FACTORY_�TUN�dG�EATURE :�����l�Ha�ndlingTo�ol ��  - �CEngli�sh Dicti�onary��OR�DEAA V�is�� Mast�er���96 H���nalog I�/O���H551���uto Sof�tware Up�date  ��J���matic B�ackup��Pa�rt&�gro�und Edit���  8\apCamera��F��t\j6R�e�ll���LOADnR�omm��shq�ޝ�TI" ��co<��
! o����pane�� 
�!��tyle �select��H�59��nD���onoitor��48�����tr��Reli�ab���adin�Diagno�s"����2�2 ua�l Check �Safety UIF lg\a���hanced Rob Serv �q ct\��lU?ser FrU���DIF��Ext.� DIO ��fi�A d��end.r Err L@��KIF�r��  �����90��FCTN_ MenuZ v'���74� TP I�n��fac  SU (G=�}p��k Excn �g�3��High�-Sper Ski.+�  sO�H9 � �mmunic!�oknsg�teur� 4����V�����conn��2��E�N��Incrs�tru���5.f�dKAREL Cmd. L?�uaA� O�Ru�n-Ti� Env�����K� ��+%�sn#�S/W��74��LicenseT��  (Au* o�gBook(Sy���m)��"
�MACROs,~V/Offse��ap��MH� �����pfa5�Mech�Stop Pro�t��� d�b i��Shif���j545�!xr ��#�ޜ�,+{b od�e Switch.��m\e�!o4=.�& pro�4���g��Mult�i-T7G��net.Pos �Regi��z�P>��t Fun����3 Rz1��Numx �����9m�1� � Adjuj��1' J7�7�* ����6tatuq1EI�KRDMto}t��scove�� ��@By- }u'est1�$Go� � �U5\SNPX� b"���YA�"Libr����#��1 �$~@h�pd]0��Jts in V�CCM�����0� 8 �u!��2 R�0��/I�08��TM�ILIB�M J9u2�@P�Acc>��F�97�TPTXl�+�BRSQelZ0�M8 Rm��q%���692��Unex�ceptr mot}nT  CVV�P���KC����+-|��~K  II)�VSP CSXC�&�.c�� e�"�� t��@Wew�A3D Q�8bvr ngmen�@�iP� �a0y�0�pfGr�idAplay �!� nh�@*�3R�1M�-10iA(B2�01 �`2V"  �F���scii�l�oad��83 M��l����Guar��d J85�0�mP�'�L`���stuaPsat�&]$Cyc���|0ori_ x%D7ata'Pqu����ch�1��g`� j6� RLJam�5��|��IMI De-By(\A�cP" #^0�C  etkc>^0asswo%q�)650�ApU�Xsnt��Pven�C�TqH�5�0Y�ELLOW BO�?Y��� Arc�0v�is��Ch�We{ldQcial4Izt�Op� ��gs֛` 2@�a��pofG yRjT1 �NE�#HT� xy�Wb��! �p�`g�d`���p\� =P��JPN ARCP*�PR�A�� O�L�pSup̂fi�l�p��J�� ��cro�670�1C~E�d���SS�pe�teex�$ �P� So7 �t� ssagN5 D<Q�BP:� �9 "0F�QrtQC��P�l0dpn�笔�rpf��q�e�ppma�scbin4ps{yn�' ptx]0�8�HELNCL� VIS PKGsS �Z@MB �&��B J8@IP�E GET_VA�R FI?S (U�ni� LU�OOL�: ADD�@29�.FD�TCm���E�@DVp���`A�Т�NO WTWTE'ST �� 6�!���c�FOR ��EC�T �a!� ALS�E ALA`�CP?MO-130��� �b D: HANG FROMg��2���R709 DR�AM AVAIL�CHECKS 5�49��m�VPCS� SU֐LIMC�HK��P�0x�FF� POS� F�� �q8-12 oCHARS�ER6��OGRA ��Z@A�VEH�AME��.#SV��Вאn$���9�m "y�TRC�v� SHADP�U_PDAT k�0���STATI��� �MUCH ���T�IMQ MOTN�-003��@O�BOGUIDE DAUGH���b��@$tou� �@C�y �0��PATH�_�MOVET�� �R64��VMXP�ACK MAY ?ASSERTjS��oCYCL`�TA���BE COR 7�1�1-�AN��RC� OPTIONS�  �`��APSH;-1�`fix��2�SO��B��XO򝡞�C_T��	�i��0j���du�byz p w1a��y�٠HI�����U�pb XSPD� TB/�F� \h�chΤB0���EN�D�CE�06\Q�p�{ smay n�@�pk��L ��tOraff#�	� ���~1from s�ysvar sc�r�0R� ��d�DJ�U���H�!A��/���SET ERR��D�P7����ND�ANT SCRE�EN UNREAO VM �PD�D���PA���R�IO� JNN�0�FI���B��GROUNנD Y�Т٠��h�SVIP 53� QS��DIGIT VERS��ká��NEW�� P06z�@C�1IMAG�hͱ���8� DI`<���pSSUE�5���EPLAN JO�N� DEL���15�7QאD��CAL�LI���Q��m���I�PND}�IMG oN9 PZ�19���MNT/��ES ܏��`LocR Ho�l߀=��2�Pn� P�G:��=�M��ca�n����С: 3�D mE2view� d X��eat1 �0b�pof Ǡ�"HCɰ�ANN�OT ACCESS M cpie�$Et.Qs a� l�oMdFlex)a:z��w$qmo G�s�A9�-'p~0��h0p�a��eJ AUTcO-�0��!ipu@�Т<ᡠIABLE�+� 7�a FPLNs: L�pl m6� MD<�VI�и�WIT HOC�;Jo~1Qui��":��N��USB�@�P�t & remo�v���D�vAxisO FT_7�PGɰ�CP:�OS-1�44 � h s s268QՐOST�p�  CRASH �DU��$P��WO�RD.$�LOG3IN�P��P:	�0��046 issu�eE�H�: Sl�ow st�cB�`6����໰IF��IMPR��SPO�T:Wh4���N1S�TY��0VMGR��b�N�CAT��4�oRRE�� � �58�1��:%�RT�U!Pe -M a�SE�:�@pp���AGpL���m@allء�*0a�OCB W�A���"3 CNTw0 T9DWroO0alarm�ˀm0d t�M�"0�2|�s o�Z@OME<�x� ��E%  #1-�gSRE��M�st}0g     5�KANJI5no� MNS@�IN�ISITALIZf'� E�f�we���6@� dr�@ fp� "��SCII �L�afails �w��SYSTE0[�i��  � Mq��1QGro8�m n�@vA����&���n�0q��RWRI� OF Lk��� �\ref"�
�up�� de-rela��Qd 03.�0S�Schőbetw�e4�IND exm ɰTPa�DO� �l� �ɰGig�E�soperab�il`p l,��H0cB��@]�le�Q0cflxz�Ð���OS {����v4pf;igi GLA�$��c2�7H� lapn�0ASB� If��=g�2 l\c�0���/�E�� EXCE 㰁�P���i�� o0��Gd`]Ц�yfq�l lxt��EFal��#0�i�xO�Y�n�CLOS��SRNq1NT^�F��U��FqKP�ANIOO V7/ॠ1�{8����DB �0���ᴥ�ED��DET�|�'� �bF�NLwINEb�BUG�Tt���C"RLIB���A��ABC JA�RKY@��� rk�ey�`IL���PRr��N��ITGAR� D$�R �Er *�T��a�U�0��h��[�ZE V� T�ASK p.vr��P2" .�XfJ�s�rn�S谥dIBP�	c���B/��BU]S��UNN� j0�-�{��cR'���L�OE�DIVS�CU�Ls$cb����BW !��R~�W`P�����IT(঱tʠ�O=F��UNEXڠ+�Ҧ�p�FtE��SV�EMG3`NML �505� D*�CC_SAFE�P*� �8ꐺ� PET��'P��`�F  !���IQR����c i S>�� K��K�H G_UNCHG��S�/MECH��M���T*�%p6u��tPORY LEAK�9J���SPEgD���2V 74\GR�I��Q�g��CTLN��TRe @�_�p l���EN'�IN�������$���r��T3\)�i�STO�A�s�L��͐X	���qb��Y� ��TO2�J m��0F<�K����SDU�S��O��3 9�J F�&��~�SSVGN-1#�I���RSRwQDAU��Cޱ� �T6�g��� �3�]���BRKCTqR/"� �q\j5�p�_�Q�S�qINVJ0D ZO�Pݲ���s ��г�Ui ɰ̒�a��DUAL� J5�0e�x�RVO117 AW�TH!Hr�%�N�247%�528��|�&aol ���RP���at�Sd�cU���P,�LER��iԗQ<0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�c�豓�{�U��ROP� 2�b�pB��IT�P4M��b !A�Ut c0< � pleste�N@� z1�^qR635 (AccuCal2kA=���I) "�ǰ�1a\�Ps��ǐ� �bЧ0P򶲊���i�g\cbacul "A3p_ �1��ն|���etaca��AT���PC�`����v�_p�.pc!�x���:�circB���5�tl��Bɵ�:�Cfm+�Ί�V�b�����r�upfrm.0����ⴊ�xed��Μ��~�pedA�D �|}b�ptlibB�� �_�rt��	��_\׊ۊ�6�fm �݊�oޢ�e��̆Ϙ�"��c�Ӳ�5�j>���F��tcȐ��	�r�����mm 1��T�sl^0��T�mѡ�#�rm3��ub Y�q�gstd}��pl;��&�ckv�=�r�vf0�䊰��9�vi�����ul�`�0fp�q ��.f��� da�q; i Data Acquisi���n�
��T`��1�89��22 �DMCM RRS�2Z�75��9 3� R710�o5�9p5\?��T ="��1 (D�T� nk@��������E �Ƒȵ��Ӹ�etdmm ��ER�����gE��1�q\mo ?۳�=(G���`[(

�2�` ! �|@JMACRO���Skip/OffCse:�a��V�4oy9� &qR662�H��s�H�
 6Bq�8����9Z�43� J77� 6�J783�o ��n��"v�R5IKC~Bq2 PTLC�vZg R�3 (�s, ��������03�	зJԷ\s�fmnmc "M�NMC����ҹ�%m;nf�FMC"Ѻ|0ª etmcr� ��8���� �,+{D6{�   874\Oprdq>,jF0����axisHP�rocess A�xes e�rol�^PRA
�Dp� 5�6 J81j�59� 56o6� ���06w�690 98� [!GIDV�1��2(x2��2ont�0�
� ���m2���?C���etis "IS�D��9�� FpraxRAM�P� D�чdefB�,�G�i�sbasicHB��@޲{6�� 708*�6��(�Acw:� �����D
�/,��AMOX�� ��DvE��?;Td��>Pi� RAFM';�]�!PAM�V�W�E�e�U�Q'
bU�75��.�ceNe� nterface^4�1' 5&!54�K��b(Devam±�/@�#���/<�Tane`�"DNEWE���bt�pdnui �AI��_s2�d_rso!no���bAsfjN�>�bdv_arFvf�`xhpz�}w��hkH�9xstc��gApocnlGzv{�ff� �r���z�3{q�'Td>pcham�pr;e�p� ^59�77��	܀�4}0��m�Ɂ�/�����lf�!�p�cchmp]aMP�&B�� �mpevp�����pcs���YeS�� Macr%o�OD��16Q!)* �:$�2U"_,��Y�(PC ��$_;������o��J�gege=mQ@GEMSW�~Z>G�gesndy��OD�ndda��S��csyT�Kɓ�su^҈����n�m���L�� ' ���9:p'ѳ�޲��spotplusp���`-�W�l��J�s��t[�׷p�key�ɰ�$��s�-����m���\featu 0FEAWD�woolo�srn'!2 p���a�As3���tT.� (N. A.)��!e!�J# (j�,��oBLIB�oD -�.�n��k9�"K��u[-��_���p� "PS�EqW����wop "sEЅ�&�:�J� �����y�|��O8�� 5��Rɺ���ɰ[��X �������%�(
���q HL�0k�
�z�a!�B�Q�"( g�Q�����]�'�.� ����&���<�!ҝ_�#��tpJ�H�~Z��j� ����y������2�� e������Z����V�� !%���=�]�͂��^2n�@iRV� on�IQYq͋JF0� 8ހȖ`�	(^�dQueue���X\1�ʖ`��+F1tpvtsn���N&��ftpJ0v �RDV�	f��J1� Q���v�en���kvstk��m�p��btkclrqq���get�����r��`ka�ck�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�mc�N+v3�_� �����.v�/\=jF��� �`Q��΋ܒ�N50 (F�RA��+��͢fraparm��Ҁ�z} 6�J643p:~V�ELSE
#��VAR $SGSYSCFG.$�`�_UNITS 2��DG~°@�4Jgfr8��4A�@FRL-��0 ͅ�3ې���L�0NE �:�=�?@�8�v�9�~Qx304��;�BP�RSM~QA�5TX�.$VNUM_O�L��5��DJ507���l� Funct�ʂ"qwAP��琉�3# H�ƞ�kP9jQ�QA5ձ� ��@jLJzB J[�6N�kAP���|�S��"TPPR����QA�prnaS�V�ZS��AS8Dj5150U�-�`cr�`8 ���ʇ�DJR`jYȑH�  �Q ��PJ6�a21��4�8AAVM �5�Q�b0 lB�`T�UP xbJ5�45 `b�`616����0VCAM� 9�CLIOn b1�5 ����`MSC8�
rP �R`\sSTY�L MNIN�`J�628Q  �`N�REd�;@�`SCH� ��9pDCSU �Mete�`ORSsR Ԃ�a04 kREIOC �a]5�`542�b9vp�P<�nP�a�`�R�`7��`�MASKg Ho�.r7 �2��`OCO :��r3@��p�b�p���r0X�|�a�`13\mn�a39 HRM"�q��q��LCHK>�uOPLG B��a�03 �q.�pHC�R Ob�pCpPo�si�`fP6 is�[rJ554�òpDSW�bM�D�pqR�ag37 }Rjr0 �1��s4 �R6�7��5�2�r5 �2�r7 �1� P6���Reg�i�@T�uFRKDM�uSaq%�4�`�930�uSNBA��uSHLB̀\suf"pM�NPI��SPVC�J52�0��TC�`"MN�рTMIL�IF�V�PAC W�pT�PTXp6.%�T�ELN N Me��09m3UEsCK�b�`UFR�`ކ�VCOR��VI�PLpq89qSXC��S�`VVF�J�T�P �q��R626.l�u S�`Gސ�2?IGUI�C���PGSt�\ŀH8�63�S�q�����q3u4sŁ684��0�a�@b>�3 :B��s1 T��96 .��+E�51 y�q5�3�3�b1 ���b1� n�jr9 ���`V�AT ߲�q75 �s�F��`�sAWSM<��`TOP u�ŀ�R52p���a80 �
�ށXY q���0� ,b�`885�QXрOLp}�"pE࠱;tp�`LCMD���ETSS���6 |�V�CPE oZ1��VRCd3
�NL:H�h��001m2Epƌ�3 f��p��4 _/165C��6l�ꌰ7PR��008� tB��9 -20-0�`U0�pF�1޲1 ��޲2L"���p���޲4��5 \�hmp޲6 RBC�F�`ళ�fs�8 ��Ҋ��~�J�7 r'bcfA�L�8\PC����"�32m0u�n��K�Rٰn�5 5E7W
n�9 z��g40 kB��3 ���6ݲ�`00iB/���6�u��7�u��8` µ������sU0�`��t �1 05\rb��2 E���K�Ȇ�j���5˰��60 ��a�HУ`:�63�jA0F�_���F�7 ڱ݀�H�8�eHЋ��cU0$��7�p��1u��y8u��9 73��L����D7� ��5t󮊱97 ��8U�1(��2��1�1:���Eh��1np�"��8(�{U1��\pyl���,࿱v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6 B���цp��1�����1�`͵155�ض157 �2��6A2�S����1b�H�2����1Π"�2��&�B6`�1<c�34 7B�5 DR���8_�B/��187y uJ�8 06��90 rBn�1 (���202 0EWE,ѱ2^��2��90�cU2�p�2��2 b��4��2�a"RB4����9\�U2�`w�<l���4 60Mp��7������b�s
5� ��3����pB"9� 3 ����`ڰR,:7 �2��V�2��5���2^��a^	9���qr����n�A5����5᥁"�8a�$Ɂ}�5B���5���B�`UA���� ��86 V�6 S�0��5�px�2�#�529 �2P^�b1P�5~�A2`���&P5��E8��5��u�!�5���ٵ544��5��R��ąP nB^z�c �(�4�����U)5J�V�5��1�1^���%�����5 b�21��gA��58�W82� rb��5N�E�5890r� 1�95 �"���� ��c8"a��|�L ���!J"5|6��^!�6��B�"8�`#��j+�8%�6B�AME�޶"1 iC��62�2�Bu�6V��d� 4���84�`ANRS�P�e/S� C@�5� �6� ��� \� ��6� �V� 3t��� T20CA�R���8� Hf� 1DH�� �AOE� �� ;,+|�� �0\�,� �!64K��ԓrA|� �1 (M-7�!/50T�[PM��P�Th:1�C�#Pe�� �3�0� 5`M7�5T"� �D8p� ��0Gc� u�4��i1-O710i�1� Skd�7j�?6�:-HS,� �RN�@�UB�xf�X�=m75sA*A6an���!/CB�B2.6A �0;A�CIB@�A�2�QF1�UB2�21� /70�S� �4�����Aj1�3p�p��r#0 B2\m*A@C��;bi"i1K�u"�A~AAU� imm7c7��ZA@I�@�D�f�A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A �5*A�EA�5B�4>\77
B7=Q�D�2�Q�$B�E7�C�D/qAHEE�W7�_|`jz@�  2�0�Ejc7�`�E"l7�@7�A
1�EH�V~`�W2%Q�R9�.�@0L_�#����"�A���b��H3s=rA/2�R5nR4�74r�NUQ1ZU�A�s\m9
1M92L2�!F!^Y:�ps� 2ci��-?�qhimQ�t  w043 �C�p2�mQ�r�H_ �H20�Evr�QHsXBSt#62�q`s����� x��Pxq350_*AF3I)�2�d�u0�@�� '4TX�0�pa3i1A3sQ25�c&��st�r�VR1%e�q0
��j1��O2� ���A�UEiy�.�‐ ț0Ch20$CXB79�#A�ᓄM Q1]�~�� 9�Q��?PQ��qA !Pvs� 5	15aU����?PŅ���ဝQ9#A6�zS*�7�qb5��1����Q��00P(��V7]u�aitE1�� �ïp?7� !?�z��{rbUQRB1PM=��Qa9��H��QQ�25L�������Q��@�L��8ܰ��y00�\ry�"R2BL��tN  ���; �1D6{�2�qeR�5���_b�3��X]1m1lcqP1�a�E�Q� 5F����!y5���@M-16Q� � f���r��Q�e� p��� PN�LT_�10��i1��9453��@8�e�|�b1l>F1@u*AY2�
��R8�Q0����RJ�J3�D}T� 85
Qg�/0��*A�!P�*A�Ð𫿽�2,ǿپ6t�6=Q��`�Pȓ��� AQ� g�*ASt]1^u�ajr I�B����~�|I�b�L�yI�\m�Qb�I�u�z�A�c3Apa9q� B6S��S��m���}��85`N�N�  �(M���f1��@�6����161��5�s`�SC��U��A�����5\set06�c����10�y�h8��a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��@���5�B��B��h`� F���X0���A:���C�M��AZ��@��4�6@i����� e�O�-	 ���f1��F �ᱦ��1F�Y	���T6HL3��U66~`���U�9dU�9D20Lf0�� Qv� ��fjq��N�� ����0v
� ��i	�\	��72lqQ2������� \chn?gmove.V���d���@2l_arf	�f~��6� �����9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�AX]��V�1\�Qn�BJ�2W�EM!`5���)�#:�64��F�e50S�\��0 �=�PV���e���逕��E�����mw7shqQSH"U��)��9�!A��(����� ,+{9�ॲTR1!��&,�60e=�4F���2��2��	 R-��� ��������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2�"�2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D��� 5V��@2cVE����dT��pt갖�1L~E��#�F�Q��9E�#De1/��RT��59���	��A�EiR������9o\m20�20��+�-u�19r4�`�E1 �=`O9`�1"ae���O�2��_$W}am�41�4�3�/d1c_std��1)Ķ!�`_T��r�_ 4\jdg�a�q�PJ %!~`-�r�+bgB���#c300�Y�5j�QpQb1�bq��vB��v25�U������qm43� �Q<W�" PsA��e��� �t�i�P�W.��c��FX.�e�kE14��44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2-a��2A;_2��QW�2�bF�(�V11�2�3�`��X5�Ra21B�J*9�a:88rJ9X�l5�m1a�0���*���(85�&� ������P6���RB,52&A����,fA�9IfI50\u�z�O@V
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq� &ŦP1��vB)e�m�x����1p� �1�D6{�27�F�K�AREL Use{ S��FCTN��� J97�FA+�� (�Q޵�p%�)?��Vj9F?(�j�Rtk208 "Km�6Q�y�j��iæPr��9�s#��v�krcfp�RCFt3���Q~��kcctme�!�ME�g����6�ma�in�dV�� ��r!u��kDº�c���o�����J�dt�F �»�.vrT�f������E%�!��5�FRjK73B�K���UER��HJ�O  J�� (ڳF���F�q�Y��&T��p�F�z��19�tAkvBr���V�h�9p�E�y�<�k������8;�v���"CT��f ����)�
І��)�V 	�6���!��qFF�� �1q���=�����O�?� $"���$��je���TCP Aut�r~�<520 H5��J53E193��9V��96�!8��9���	 �B574��52��Je�(�� Se %!Y�����u��ma�Pqtool�ԕ�������conre�l�Ftrol Reliable�RrmvCU!��H51������ a551xe"�CNRE�I�c�&��it�l�\sfutst �"UTա��"X�\�u��g@�i�6Q]V0H�B,Eѝ6A� �Q �)C���X��Yf�Iȴ1|6s@6i��T�6IU��vR�d�
$e0%1��2�C58�E6���8�Pv�iV4OFH5�8SOeJ� mvBM6E~O58�I�0�E�# +@�&�F�0���F�P 6a���)/++�</N)0\tr1�����P� ,+{ɶ�rma;ski�msk�aA����ky'd�h	A	�P��sDisplay�Im�`v����J8�87 ("A��+He<ůצprds��I�T:���h�0pl�2�R�2��:�Gt�@��PRD�TɈ�r�C�@Fpm��D�Q�Asca��� V<Q&��bVvbrl�eې@��^S��8&5Uf�j8710��yl	��Uq���7 �&�p�p��P^@�P�firmQ����Pp� 2�=bk�6�r�3��6���tppl��PL ���O�p<b�ac�q	� �g1J�U�d�J��gait_9e��Y�&���Q���	�Shap���erationx�0��R67451tj9(`sGen� ms�42-f��r�p�50����2�rsgl�E���p�G���qF�205�p�5S���Ձ�ret�sap�BP�O�\s>� "GCR�ö?� �qngda�G ��V��st2axU�b�Aa]��bad�_|�btputl/��&�e���tplibB_��=�2.����5�Ό�cird�v�sl8p��x�hex��v��re?�Ɵx�key��v�pm��x�u9s$�6�gcr��F�������[�q27j92|�v�ollismq�Sk�9O�ݝ� (Gpl.���t��p!o���29$Fo8��cg7�no@�tptcls` CLS�o�b�\�#km�ai_
�s>�v�o	�t�b���ӿ�E��H��6�1en�u501�[m��u�tia|$calm�aUR��CalMa;teT;R51%�i=1]@-��/V� ��Z��� �fq1�9 "KA9E�L����2m��CLMTq�S#��et �LM3!} �:F�c�nspQ�cӞ��c_moq��� ���c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ����N�ve��C�clm��&Ao# �|$fin�de�0ST�D ter Fi?LANG���R��
��n3��z0gCen���r,�� ����J����� ��� K��Ú�=���_Ӛ����r� "FND�R�� 3��f��tguid�䙃N�."��J�tq�� ��������������J����_@������c��	m��Z��\fndr. ��n#>
B2p��Z�CP Ma�����C38A��� c��6� (���N�B����� �� 2�$�81��!m_���"ex�z 5�.Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$ �r*$��*$r*$%/s#�C�d/.,P�/0*ʲDPN��$���$�*�Gr�$k Ex�c�'IF�$MAS}K�%93 H5�%�H558�$548 H�$4-1�$��#21(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�4�9�0�4a�3�9j0"�M�49�4  �x�4�4tpsh��x�4�P�4- DQ� @�3�Q�4�R�4�pR%0 �2�r�4.b
E\���5�A�4��3adq\>�5K979":E�a~jO l "DQ^E^�3i�Dq ��4�R�O ?R�? ��q�5 ��T��3rAq�O�L#st�5~��7p�5��0REJ#�2�@av^Eͱ��F���4��.�5y �N� �2il(in8�4��31 JH1�2�Q4�251ݠ�4rmal� �3)�REo� Z_�æOx����4��^F�?onorTf��7_�ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4�REM���4yݱ"u@�RER5932fO��4�7Z��5lity,��U��e"Dil\��5��o ��798�7�?�25 �3hk9 10�3��FE�0=0|P_�Hl\mhm�5 ��qe�=$�^�
E���u�IAymptm`�U��BU��vste� y\�3��me�b�DvI� [�Qu�:F�Ub�*_��
E,�su��_ Er��ox���4�huse�E-�?�s�n�������FE��,�b#ox�����c݌," �������z��M�x�g��pdspw)� 	��9���b���(��1���c��Y� R�� �>�P���W��� �����'�0ɵ��[��͂���  ߤ ,+@� ��A�bum�pšf��B*�Bo!x%��7Aǰ60�BB�w���MC� (6�,�f�t I�s� ST��*��}B���z��w��"BBF
��>�`���)��\bbk968 "�X4�ω�bb�9vas69����etbŠb��X�����ed	��F��u�f� �seDa"������'�\��@,���b�ѽ�o6�$H�
�x�$�f���!�y���Q[�! tp�err�fd� T�Pl0o� Reco�v,��3D��R642 � 0��C@}s�� N@��(U�rr�o���yu2r���  �
  |����$$CLe�? �������������$z�_D�IGIT��������.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo�$j��+c:PRO�DUCTM�0\P_GSTKD��V&o�hozf99��D����$FEAT?_INDEX��xd���  �
�`ILECO_MP ;���#���`�cSETU�P2 <�e~�b�  N �a��c_AP2BCK� 1=�i  #�)wh0?{%&c����Q�xe%� I�m���8�� \�n����!���ȏW� �{��"���F�Տj� ��w���/�ğS���� �����B�T��x�� ����=�үa������ ,���P�߯t������ 9�ο�o�ϓ�(�:� ɿ^���Ϗϸ�G� ��k� �ߡ�6���Z� l��ϐ�ߴ���U��� y����D���h��� ���-���Q������ ���@�R���v���� )�����_�����* ��N��r��7 ��m�&�3�\�i
pP 2>#p*.VRc�*��� /���PC/1/OFR6:/].��/+T�`�/�/F%�/��,�`r/?�*.F�8?	H#&?e<��/�?;STM @�2�?�.K �?�=�iPendant Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OoO�O_:JPG  _J_�56_�O_�_��	PANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W �o�o�o)�Z4�o[��WI��
T�PEINS.XM)L��0\����qCustom Toolbar	���PASSWO�RDyFRS�:\L�� %P�assword ?Config��� ֏e�Ϗ�B0���T� f����������O�� s������>�͟b�� [���'���K��򯁯 ���:�L�ۯp����� #�5�ʿY��}��$� ��H�׿l�~�Ϣ�1� ����g��ϋ� ߯��� V���z�	�s߰�?��� c���
��.��R�d� �߈���;�M���q� �����<���`���� ��%���I������ ��8����n���! ��W�{"� F�j|�/� Se��/�/T/ �x//�/�/=/�/a/ �/?�/,?�/P?�/�/ �??�?9?�?�?o?O �?(O:O�?^O�?�O�O #O�OGO�OkO}O_�O 6_�O/_l_�O�__�_ �_U_�_y_o o�_Do �_ho�_	o�o-o�oQo �o�o�o�o@R�o v��;�_� ��*��N��G��� ���7�̏ޏm���� &�8�Ǐ\�돀��!� ��E�ڟi�ӟ���4� ßX�j��������į S��w������B�#���$FILE_D�GBCK 1=���/���� ( �)
�SUMMARY.�DGL���MD:����Dia�g Summar�y��Ϊ
CONSLOG�������D��ӱConsol�e logE�ͫ���MEMCHEC�K:�!ϯ���X�M�emory Da�ta��ѧ�{)}��HADOW���ϵ�J���Sha�dow Chan�gesM�'�-�?�)	FTP7Ϥ��3ߨ���Z�mme?nt TBD��ѧ�0=4)ETHERNET��������T�ӱEthe�rnet \�fi�guration�U�ؠ��DCSVR�F�߽߫�����%��� verif�y all��'�1�PY���DIFF������[���%��diff]�����1R�9�K��� ����X��CHGD������c��!r����2ZAS� ���GD���k��8z��FY3bI[� �/"�GD���s/�����/*&UPDA�TES.� �/���FRS:\�/�-�ԱUpdates� List�/��P�SRBWLD.C	M(?���"<?�/Y��PS_ROBOWEL��̯�?�?��? &�O-O�?QO�?uOO nO�O:O�O^O�O_�O )_�OM___�O�__�_ �_H_�_l_o�_�_7o �_[o�_lo�o o�oDo �o�ozo�o3E�o i�o���R� v���A��e�w� ���*���я`����� ����O�ޏs���� ��8�͟\�����'� ��K�]�쟁����4� ��ۯj������5�į Y��}������B�׿ �x�Ϝ�1���*�g� ����Ϝ���P���t� 	�ߪ�?���c�u�� ��(߽�L߶��߂�� ��(�M���q� ��� 6���Z������%��� I���B�����2������h����$FI�LE_� PR� ���������MDON�LY 1=.�� 
 ���q�� ��������~ %�I�m� 2��h��!/� ./W/�{/
/�/�/@/ �/d/�/?�//?�/S? e?�/�??�?<?�?�? r?O�?+O=O�?aO�? �O�O&O�OJO�O�O�O�_�O9_�OF_o_
VISBCKL6[*.VDv_�_.P�FR:\�_�^�.PVision� VD file �_�O4oFo\_joT_�o o�o�oSo�owo �oB�of�o�+ �������+� P��t������9�Ώ ]�򏁏��(���L�^� ������5���ܟk�  ���$�6�şZ��~������
MR_G�RP 1>.�L��C4  B���	 W������*u����RHB ��2� ��� ��� ���B�����Z� l���C���D��������Ŀ��J8�L��(�J���F��5U��R������ֿ Gn��E��.E88��-���:u��{@ ����@AߍA���f�?h?!A��fr���E�� F@ �������ھ��NJ�k�H9�H�u��F!��IP�s�?����(��9�<9��896C'�6<,6\b� �+�&�(�a�L߅�p�A��A��߲�v��� r������
�C�.�@� y�d��������������?�Z�lϖ�BH�� �Ζ��������
0�PJ��P�K}��ܿ� ��B���/ ��@�3�3:��.�gN�U�UU�U��q	>u?.�?!rX���	�-=[�z�=�̽=�V6<�=�=��=$q������@8�i7G���8�D�8?@9!�7��:����D�@ ?D�� Cϥ��+C������'/0- ��P/����/N��/r� �/���/�??;?&? _?J?\?�?�?�?�?�? �?O�?O7O"O[OFO OjO�O�O�O�O�г� ���O$_�OH_3_l_W_ �_{_�_�_�_�_�_o �_2ooVohoSo�owo �o�i��o�o�o�� );�o_J�j� ������%�� 5�[�F��j�����Ǐ ���֏�!��E�0� i�{�B/��f/�/�/�/ ���/��/A�\�e�P� ��t��������ί� �+��O�:�s�^�p� ����Ϳ���ܿ� � �OH��o�
ϓ�~Ϸ� �����������5� � Y�D�}�hߍ߳ߞ��� �����o�1�C�U� y��߉�������� ����-��Q�<�u�`� �������������� ;&_J\�� ��������ڟ� F�j4����� ����!//1/W/ B/{/f/�/�/�/�/�/ �/�/??A?,?e?,� �?P�q?�?�?�?�?O �?+OOOO:OLO�OpO �O�O�O�O�O�O_'_ _K_�o_�_�_�_l� �_0_�_�_�_#o
oGo .okoVoho�o�o�o�o �o�o�oC.g R�v����� 	���<�`�*< ��`�����ޏ�� )��M�8�q�\����� ��˟���ڟ���7� "�[�F�X���|���|? ֯�?�����3��W� B�{�f�����ÿ���� �����A�,�e�P� uϛ�b_�����Ϫ_�� ߀�=�(�a�s�Zߗ� ~߻ߦ�������� � 9�$�]�H��l��� ����������#��G� Y� �B�������z��� ����
ԏ:�C.g Rd������ 	�?*cN� r�����/̯ &/�M/�q/\/�/�/ �/�/�/�/�/?�/7? "?4?m?X?�?|?�?�? �?�?��O!O3O��WO iO�?�OxO�O�O�O�O �O_�O/__S_>_P_ �_t_�_�_�_�_�_�_ o+ooOo:oso^o�o �op��o�� ��$ ��o�o�~� ������5� � Y�D�}�h�������׏ ����
�C�.�/ v�<���8������П ����?�*�c�N��� r��������̯�� )��?9�_�q���JO�� ���ݿȿ��%�7� �[�F��jϣώ��� ��������!��E�0� i�T�yߟߊ��߮��� �o�o��o>�t� >��b��������� ��+��O�:�L���p� ������������' K6oZ�Z�|� ~�����5  YDi�z��� ���/
//U/@/ y/@��/�/�/�/���/ ^/???Q?8?u?\? �?�?�?�?�?�?�?O O;O&O8OqO\O�O�O �O�O�O�O�O_�O7_���$FNO ����VQ�
F0fQ} kP FLAG8��(LRRM_CHKTYP  WP���^P�WP��{QOM�P_MIN܇P����P� � XNPSSB_�CFG ?VU? ��_����S ooIUTP_�DEF_OW  ���R&hIRC�OM�P8o�$GE�NOVRD_DO�V�6�flTHR֨V d�edkd_E�NBWo k`RA�VC_GRP 19@�WCa X"_�o _1U<y� r�����	�� -��=�c�J���n��� �����ȏ����;��"�_�F�X���ibRO�U�`FVX�P��&�<b&�8�?��埘����>���  D?�јls���@@g�B�7��p�)�ԙ���`SMT
�cG�mM���� ��LQHOSTC�R19H���P��at��SM��f��\���	127.�0��1��  e ��ٿ�����ǿ@��R�d�vϙ�0�*�	a�nonymous������������0�([�� � ����� r����ߨߺ�����-� ��&�8�[�I�π� ������1�C� �W�y���`�r����� �ߺ�������%�c� u�J\n������ ���M�"4F X��i����� �7//0/B/T/� ��m/��/�/�/ ??,?�/P?b?t?�? �/�?��?�?�?OO e/w/�/�/�?�O�/�O �O�O�O�O=?_$_6_ H_kOY_�?�_�_�_�_ �_'O9OKO]O__Do�O hozo�o�o�o�O�o�o �o
?o}_Rdv ���_�_oo!� Uo*�<�N�`�r��o�� ����̏ޏ�?Q&��8�J�\���>�ENT� 1I�� P!\􏪟  ���� ՟ğ�������A�� M�(�v���^������ ���ʯ+�� �a�$� ��H���l�Ϳ����� ƿ'��K��o�2�h� �ϔ��ό��ϰ���� ���F�k�.ߏ�R߳� v��ߚ��߾���1����U��y�<�QUICC0��b�t����A1�����%���2&����u�!ROU�TERv�R�d���!?PCJOG�����!192.168.0.10���w�NAME !���!ROBOT�p�S_CFG �1H�� ��Auto-s�tarted�tFTP���� ��� 2D�� hz����U�`�
//./A�#�� ��~/����/�/ �/�/� ?2?D?V?h? �/?�?�?�?�?�?�? ���@O?dO�/�O �O�O�O�?�O�O__ *_MON_�Or_�_�_�_ �_	OO-O�_A_&ouO Jo\ono�o�o=o�o�o �o�oo�o4FX j|�_�_�_o� 7o��0�B�T�#x� ���������e���� �,�>�����ŏ ���Ο������ :�L�^�p�����'��� ʯܯ� �O�a�s��� ��l���������ƿؿ ����� �2�D�g�� zόϞϰ����#�5� G�I��}�R�d�v߈� ��iϾ��������)߀��<�N�`�r��XS�T_ERR J�5
���PDUSI�Z  ��^J�����>��WRD �?t��  �guest }��%�7�I�[�m�$�SCDMNGRPw 2Kt�������V$�K��� 	P01.�14 8��  � y����B    ;������ ���������
 �������������~����C.gR�|���  i�  �  
��������� +��������
����l .r�
��"�l��� m
�d������_G�ROU��L�� e�	����07EQUPD  	ղ��J�TYa �����TTP_A�UTH 1M��� <!iPen'dany��6�Y�!KAREL�:*��
-KC�///A/ VISION SETT�/v/�"�/�/�/ #�/�/
??Q?(?:?��?^?p>�CTRL� N����5�
��FFF9E�3�?�FRS:DEFAULT�<�FANUC �Web Server�:
�����<�kO}O�O�O�O�O��W�R_CONFIGw O�� �?���IDL_CPU�_PC@�B���7P�BHUMI�N(\��<TGNR_�IO������PN�PT_SIM_D�OmVw[TPMO_DNTOLmV �]_PRTY�X7RTOLNK 1P����_o!o3oEoWo|io�RMASTElP���R�O_CFG��o�iUO��o�bC�YCLE�o�d@_?ASG 1Q����
 ko,>Pb t�������p��sk�bNUM�����K@�`IPCH��o��`RTRY_�CN@oR��bSC�RN����Q��� �b�`�bR���Տ���$J23_D_SP_EN	�����OBPROC��U�iJOGP1�SY@��8��?�!�T�!�?*�P�OSRE�zVKANJI_�`��o_��$ ��T�L�6͕����CL_LGP<�_����EYLOGGI�N�`��L�ANGUAGE YYF7RD w����LG��U�?⧕��x� �����Z=P��'0��$� NMC:\RSCH\00\���LN_DISP V��
���������OC�R.RDzVT=�#�K@9�BOOK W
{��i��ii��X�����ǿٿ�����"��6	h�����e�?��G_BUFF 1%X�]��2	ա� ������������ !�N�E�W߄�{ߍߺ� �����������J�����DCS Z>r� =����^π+�ZE��������a�I�O 1[
{ ُ!� �!�1�C�U� i�y������������� ��	-AQcu@�������EfP/TM  �d�2 /ASew��� ����//+/=/�O/a/s/�/�/��S�EV����TYP�/??y͆��RS@"��×�F�L 1\
���� ��?�?�?�?�?�?�?�/?TP6��">>�NGNAM�ե��U`�UPS��GI�}�𑪅mA_LO{AD�G %��%DF_MOT�N���O�@MAXUALRM<��J��@sA�Q����WS ��@C �]m�-_���MPt2�7�^
{ رƭ	�!P�+ʠ�;_/��Rr�W�_�WU�W�_��R	o�_ o?o"ocoNoso�o�o �o�o�o�o�o�o; &Kq\�x�� �����#�I�4� m�P���|���Ǐ��� ֏��!��E�(�i�T� f�����ß��ӟ��� � �A�,�>�w�Z��� ����ѯ����د�� �O�2�s�^��������Ϳ���ܿ�'��BD�_LDXDISA�X@	��MEMO_{APR@E ?�+
 � *�~ϐπ�ϴ����������@I�SC 1_�+ ��IߨT��Q�c�� �߇��ߧ�����w�� ��>�)�b�t�[��� ��{����������:� ��I�[�/�������� ����o�����6!Z lS��s�� ��2�AS' �w����g���.//R/d/�_M?STR `�-w%�SCD 1am͠ L/�/H/�/�/?�/2? ?/?h?S?�?w?�?�? �?�?�?
O�?.OORO =OvOaO�O�O�O�O�O �O�O__<_'_L_r_ ]_�_�_�_�_�_�_o �_�_8o#o\oGo�oko �o�o�o�o�o�o�o" F1jUg�� �������B� -�f�Q���u�����ҏ�h/MKCFG �b�-㏕"LTA�RM_��cL�� σQ�N�><�METPUI�ǂ����)NDSP_CMNTh����|�  d�.���ς�ҟܔ|�POS�CF����PST�OL 1e'�4@�<#�
5�́5� E�S�1�S�U�g����� ��߯��ӯ���	�K� -�?���c�u�����|��SING_CHK�  ��;�ODA�Q,�f��Ç��D�EV 	L�	�MC:!�HSIZ�Eh��-��TAS�K %6�%$1�23456789� �Ϡ��TRIGw 1g�+ l6�%���ǃ�����8��p�YP[� ��EM_INF 1h3�� `)�AT&FV0E�0"ߙ�)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ������H������A���AI�q�,���|���� ���� ������J���n���� ��W�����������" ����X��/���� e������0� T;x�=�as ��/�,/c=/b/ �/A/�/�/�/�/� �?���^?p?#/ �?�/�?s?}/�?�?O �?6OHO�/lO?1?C? U?�Oy?�O�O3O _�?�D_�OU_z_a_�_�O�NITOR��G �?5�   	�EXEC1Ƀ�R2*�X3�X4�X5�X����V7�X8�X9Ƀ �RhBLd�RLd�RLd�R Ld
bLdbLd"bLd.b�Ld:bLdFbLc2Sh2�_h2kh2wh2�h2��h2�h2�h2�h2*�h3Sh3_h3�R��R_GRP_SV� 1in���(ͅ��
�Å���6�_MOx�_D=R^���PL_NAME� !6��p�!�Default� Persona�lity (from FD) ��RR2eq 1j)TUX)TX��q��X dϏ8�J�\� n���������ȏڏ� ���"�4�F�X�j�|������2'�П��� ��*�<�N�`�r��<��������ү������,�>�P�b� �R�dr 1o�y �\��, �3��~�� @D�  ��?�����?䰺�㱏A'�6����;��	lʲ	 �xJ����� ��< �"�� ��(pK�K� ��K=*�J����J���J�V���Z�����rτ́p@j��@T;f���f���ұ]�l��I��p������������b��3��´  �
`�>����b����z���ΐr�Jm��
�  B�H�˱]Ӂt�q�	�� p�  �P�pQ�p��p| � Ъ�g���c�	�'� � ���I� �  {����:�È
�?È=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁ryN���  '�������@2��@�c����/�C��}C�C�@ C�������
�AT�W�@<�P�R�%
h�B�b�A��j������:��Dz ۩��߹�����j���( �� -��C���'�7L�����q�Y������ �?�ff ���gy �����q:a��
�>+�  PƱj�( ����7	���^|�?����xZ��p<
6b<���;܍�<����<� <�&Jσ�AI�ɳ+�|���?fff?I��?&�k�@�.���J<?�` �q�.�˴fɺ�/ ��5/����j/U/�/ y/�/�/�/�/�/?�/0?q��F�?l? ?�?/�?+)�?�?ؿE�� E�I�G+� F��?)O �?9O_OJO�OnO�Of�BL޳B�?_h�.� �O�O��%_�OL_�?m_ �?�__�_�_�_�_�
��h�Îg>���_Co�_goRodo��o�GA�ds�q�C��o�o�o|���ؠ$]Hq���D���pC���pCHmZZ7t���6q�q���ܶN'�3A�A��AR1AO��^?�$�?��K�0±
=ç�>����3�W�
=�#�W��e��9�����{�����<���(�B�u���=B0��?����	L���H�F�G����G��H�U`�E���C�+����I#�I���HD�F���E��RC�j�=��
I���@H�!H�(� E<YD0 q�$��H�3�l�W� ��{��������՟� ��2��V�A�z���w� ����ԯ������� �R�=�v�a������� �����߿��<�'� `�Kτ�oρϺϥ��� �����&��J�\�G� ��kߤߏ��߳����� ��"��F�1�j�U�� y������������0��T�?�Q����(��1��3/E��<���5������q3�8�����q�4Mgs&I�B+2D�a���{�^^	�������uP2P7Q4_A��M0bt��R�������/   � /�b/P/�/t/�/ *�a)_3/�/�/�% 1a?�/?;?M?_?q?  �?�/�?�?�?��?O 2 F��$�vGb�/�A���@�a�`�qC��C@��o�O2���OF�� DzH@�� F?�P D���O�O�ys<O!_3_E_W_�i_s?���@@*pZ.t22!u2~
 p_ �_�_�_	oo-o?oQo couo�o�o�o�o��Q� ��+��1���$MSKCFM�AP  �5� �6�Q�Q�"~�cONREL  
q3�bEXCFENB?wq
s1uXqFNC_�QtJOGOVLI�M?wdIpMrd�bK�EY?w�u�bR�UN�|�u�bS?FSPDTY�av<Ju3sSIGN?Qt�T1MOT�Nq��b_CE_GRP� 1p�5s\ r���j�����T��� �������<��`�� U���M���̟��🧟 �&�ݟJ��C���7� ������گ��������4�V�`TCOM_�CFG 1q}иVp�����
P�_A�RC_\r
jyU?AP_CPL��nt�NOCHECK {?{ 	 r��1�C�U�g�y� �ϝϯ���������	���({NO_WAI�T_L�	uM�NT�X�r{�[m�_7ERRY�2sy3� &�������r��c� ��T_M�O��t��,  \��$�k�3�PARAuM��u{��V`[��!�u?�� =9@�345678901��&���E�W�3� c�����{������� �����=�U�M_RSPACE� �Vv��$OD�RDSP���jxO�FFSET_CAsRTܿ�DIS���PEN_FIL�E� �q��c֮�OPTION_IO���PWORK 5v_�ms �P(�R$0uj.j�	 ��Hj(6$�� RG_DSBL'  �5Js�\���RIENTTO�>p9!C��Pq=�#�UT_SIM_D
r�b� �V� LCT w�w�bc��U)+$_P�EXE�d&RAT�p �vju�p��2X�j�)TUX)TX�>##X d-�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?O�H2�/oO �O�O�O�O�O�O�O�O_]�<^O;_M___q_ �_�_�_�_�_�_�_o����X�OU[�o(��(���$}o�, ���IpB` @D�  &Ua?�[cAa?��]a�]�DWcUa쪋l;��	lmb�`��xJ�`������a�<; ��`� ��b, �H(��H3k7�HSM5G�22�G���Gp
��
�!��'|, KCR�>�>q�Gs�uaT�3���  �4spBpyr  ]�o�*SB_�����j]��t�q� ��rna ��,���6  U��PQ��|N�M�,k�!�	�'� � ���I� �  {��%�=��ͭ�迋ba	���I  �n @� �~���p�����& �N U�[�'!o�t:q�pC\�C�@@s�Bq�|��� m�
S�A\��h@ߐ�n�����Z�B\��A8���p� �-�qbz�P��t�_�������( �� -��恊�n�ڥ[A]Ѻ�b4�'!���(p �?�fAfo��
����O�Z�R��8��z���>N΁  Pia��(�� ��@���ک�a�c�dF#/?����x�����<
6b<߈�;܍�<�ê�<� <�&�o&�)�A�lcΐIƾ*�?fff?�?y&c���@�.u��J<?�`�� Yђ^�nd��]e��[g ��Gǡd<����1�� U�@�y�dߝ߯ߚ��� �߼�	���-�������&��"�E�� E���G+� F� ������������&���J�5��bB��A T�8�ђ��0�6���>� ��J�n�7��[mx�0��h��1��>�M�I`
�@��A�[��C-�)��?���� /�
YĒ��Jp��vav`#CH/�������}!@I�Y�'��3A�A�AR�1AO�^?�$��?����±�
=ç>�����3�W
=�#�����+e��ܒ������{�����<��.(��B�u��=�B0�������	�*H�F��G���G���H�U`E����C�+�-I#��I��HD��F��E���RC�j=U>
�I��@H��!H�( E<YD0/�?�?�? �?�?O�?3OOWOBO TO�OxO�O�O�O�O�O �O_/__S_>_w_b_ �_�_�_�_�_�_�_o o=o(oaoLo�o�o�o �o�o�o�o�o' $]H�l��� ����#��G�2� k�V���z���ŏ��� ԏ���1��U�g�R� ��v�����ӟ��������-��(���������a�����Q�c�,!3�8��}���,!4Mgs8����ɢIB+կ���a���{� ��A�/�e�S���w�J�P!�P��������7��ӯ�ϑ�R9�Kτ�oχϓϥ�  ���χ���� )��M����������{߉ߛ���ߒߤ�p������  )�G�q�_���2� F�$�&Gb	���n�[ZjM!C�s�@j/�A�S�~��F� Dz����� F�P DC��W����)������������x?̯��@@
9�RE�E��E��
 v��� ����*<pN`�*P �������1��$PA�RAM_MENU� ?-���  DEFPULSEl�	WAITTM�OUT�RCV�� SHEL�L_WRK.$CUR_STYL�;,OPT�/�PTB./("C�R?_DECSN��� ,y/�/�/�/�/�/�/ ?	??-?V?Q?c?u?��?�USE_PR_OG %�%�?\�?�3CCR������7_HOST !�!�44O�:AT̰�?PCO)ARC|�O�;_TIME��XB�  �GD�EBUGV@��3G�INP_FLMS�K�O�IT`��O�EP+GAP �L��#[�CH�O�HTYPE
����?�?�_�_ �_�_�_oo'o9obo ]ooo�o�o�o�o�o�o �o�o:5GY� }����������1�Z��EWOR�D ?	7]	�RS`�	PNS2�$��JOE!>��TEs@WVTRA�CECTL 1xv-�� ���Ӱ��ɆDT� Qy-����D � �� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� T�(�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_j��_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�_����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv��������//"#�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �#|"DEF�SPD |�,l!!J �8 IN �TRL }�-�" 8�%�!PE_C�ONFI� ~g%O�g!�$�%��$LID�#�-~74GRP 1�7�Q!�#!A ����&ff"!A+�33D�� D]�� CÀ A@+6�!�" d�$�9�9�*1*0� 	 �+9�(�&�"�? ´	C�?�;B@3AO�?�OIO3OmO"!>�T?�
5�O�O�N��O =��=#�
�O_�O_J_5_ n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_Roxoco�o �o�o�o�o�o�o�>)bM��;
�V7.10bet�a1�$  �A�E�rӻ��A " �p?!G�^�q>���r��0��q�ͻqBQ��qA\�p�q�4�q*�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏� ��4��1�j�U���y� ����֟������0� �T�?�x�c������� ү����!o�,�ۯP� ;�M���q�����ο�� �ݿ�(��L�7�p�x+9��sF@ �� �ͷϥ�g%������ +�!6I�[߆������� �ߠ���������!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ���=(aL ^������ �'9$]�Ϛ��� ��������/<� 5/`�r߄ߖߏ/>�/ �/�/�/�/?�/1?? U?@?R?�?v?�?�?�? �?�?�?O-OOQO<O uO`O�O�O�O�O���O _�O)__M_8_q_\_ n_�_�_�_�_�_�_o �_7oIot���o�o ���o�o�o(/!L/ ^/p/�/{*o��� ������A�,� e�P�b���������� Ώ��+�=�(�a�L� ��p������Oߟ񟠟 � �9�$�]�H���l� ~�����ۯƯ���#� No`oro�on��o�o�o �oԿ���8J\ ng����vϯϚ��� ����	���-��Q�<� u�`�r߫ߖ��ߺ��� ����;�M�8�q�\� ��������z������ %��I�4�m�X���|� ����������:�L� ^���Z�������� ���$�6�H�S wb����� ��//=/(/a/L/ �/p/�/�/�/�/�/? �/'??K?]?H?�?�� �?�?f?�?�?�?O�? 5O OYODO}OhO�O�O �O�O�O�O&8J4_ F_����_�_��_ �_"4-o�O*oco No�oro�o�o�o�o�o �o)M8q\ �������� �7�"�[�m��?���� R�Ǐ���֏�!�� E�0�i�T���x����� ���_$_V_ �2�l_�~_�_�����R�$P�LID_KNOW�_M  �T������SV� ��U͠�U��
��.� ǟR�=�O�����mӣ�M_GRP 1�T�!`0u��T@ٰ)o�ҵ�
���P зj��`���!�J� _�W�i�{ύϟϱ���`������߱�MR��Ņ��T��s�w�  s��ߠ޴߯߅��ߩ� ������A���'�� ����������� ��=���#����������}������S��ST^��1 1��U# ����0�_ A  .��,>Pb�� ������3 (iL^p���(��2*��'�<-/3/)/;/M/4f/x/�/�/�5�/�/�/�/6 ??(?:?7S?e?w?�?8�?�?�?�?~MAD  d�#`PARN_UM  w�\%OSCH?J ME�
�G`A�Iͣ�EUP�D`OrE
a�OT_CMP_��B@�P@�'˥TER_C;HK'U��˪?R�$_6[RSl�¯��_#MOA@�_�U_�_RE�_RES_G � �>�oo8o+o\o Oo�oso�o�o�o�o�o@�o�o�W �\�_ %�Ue Baf�S�  ����S0��� �SR0��#��S�0>� ]�b��S�0}������R�V 1�����rB@�c]��t�(@�c\����D@�c[�$���RTHR_INRl�DA��z˥d,�MASS9�� ZM�MN8�k�M�ON_QUEUE� ���˦��x� URDNPUbQN{�P[��END���_ڙ�EXE�ڕ�@BE��ʟ��OPTIO�Ǘ�[��PROGR�AM %��%�ۏ�O��TASK�_IAD0�OCFG� ���tO��ŠD�ATA���Ϋ@��27�>�P�b�t� ��,�����ɿۿ������#�5�G���INFOUӌ�������� �Ͽ���������+� =�O�a�s߅ߗߩ߻�@�������^�jč�� yġ?PDIT� �ίc���WE�RFL
��
RG�ADJ �n�A	����?����@���?IORITY{�QV}���MPDSPH������Uz����O�TOEy�1�R�� (!AF4�E��P]���!tc�ph���!ud|��!icm���ݏ6�XY_ȡ��R��ۡ)� *0+/ ۠�W :F�j���� ��%7[B��*��PORTT#�BC۠�����_CARTREP�
�R� SKSTA�z��ZSSAV����n�	2500H863���r�$!�U�R����q��n�}/�/�'� URGeE�B��rYWF� #DO{�rUVWV��$��A�WRUP_DELAY �R�>�$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?3A_QSKIP!�n�;l#x 	1/+O + OROdOvO9Hn��O �G�O�O�O�O�O_�O _D_V_h_._�_z_�_ �_�_�_�_
o�_.o@o Roovodo�o�o�o�o �o�o�o*<L�r`���n��$�RCVTM���]��pDCR!�L�ЈqC`N�C����C�Q?���>r��<�|�{4M�g�&���/��Z���t����l4��{�4Oi��O �<
6b<���;܍�>u.��?!<�&{�b�ˏݏ��8��� ��,�>�P�b�t��� ������Ο���ݟ� �:�%�7�p�S����� �ʯܯ� ��$�6� H�Z�l�~�������ƿ ���տ���2�D�'� h�zϽ��ϰ������� ��
��.�@�R�d�O� �ߚ߅߾ߩ������ ���<�N��r��� �����������&� 8�#�\�G�����}��� ��������S�4F Xj|����� ����0T? x�u����' //,/>/P/b/t/�/ �/�/�/�/�/�?�/ (??L?7?p?�?e?�? �?��?�? OO$O6O HOZOlO~O�O�O�?�? �O�O�O�O __D_V_ 9_z_�_�?�_�_�_�_ �_
oo.o@oRodovo��X�qGN_ATC� 1�� �AT&FV0E�0�kATDP�/6/9/2/9��hATA�n,�AT%G1%�B960�i+�++�o,�aH,��qIO_TYPE'  �u�sn_�o�REFPOS1 �1�P{ x�o�Xh_�d_�� ���K�6�o�
����.���R����{{2 1�P{���؏V��ԏz����q3 1� �$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����|<���S6 1�ѯ����/�����ѿO�S7 1�f�x���Ŀ�B�-�f��S8 1�����Y��������y�SMASK 1�P  
9�G��'XNOM���a~���ӁqMOTE  �hܗ�_CFG ᢥ����рrPL_RANG�ћQ����OWER ��e����SM_DRYPRG %i��%��J��TART� �
�X�UME_PRO'�9��~t�_EXEC_EN�B  �e��GS�PD������c��T3DB���RM��MT_!�T�ߓa�OBOT_NAM/E i���i�OB_ORD_N_UM ?
�\q�H863 � �T���������bPC_TIME�OUT�� x�`S�232��1��k� LTEAC�H PENDAN �ǅ�}���`�Mainten�ance Con�s�R}�m
"{�dKCL/Cg��Z ��n� No Use}�	��*NPO��х����(CH�_L���]���	��mMAVAI�L��{���SPACE1 2��| d��(>���&���p��M,8�?�ep/eT/ �/�/�/�/�W//,/ >/�/b/�/v?�?Z?�/ �?�9�e�a�=??,? >?�?b?�?vO�OZO�?��O�O�Os�2� /O*O<O�O`O�O�_��_u_�_�_�_�_[3 _#_5_G_Y_o}_�_ �o�o�o�o�o[4.o@oRodovo$�o �o����"�	�7�[5K]o��A� ���	�̏�?�&�T�[6h�z������� ^�ԏ���&��;�\�C�q�[7�������� ͟{���"�C��X�y�`���[8����Ư دꯘ��0�?�`�#��uϖ�}ϫ�[G ��i� �ϋ
G� ����$�6� H�Z�l�~ߐ��8 ǳ�@����߈��d(� ��M�_�q���� ��������?���2� %�7�e�w��������� �����������!�R E�W�����������?Q; `�� @0�@�ߖrz	�V_ �����
/L/^/ |/2/d/�/�/�/�/�/ �/?�/�/�/*?l?~? �?R?�?�?�?�?�?�?�?2O�?
��O[�_MODE  ��˝IS ���vO,*ϲ�O-_���	M_v_#dCWO�RK_AD�M7{��%aR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/D���d;2BaR��WY��^����^R^	r  P���� �  �8�P�	�D��GYk}� �������Qp/@/R//<)P;�o\T���Qpg-�t��_DiKT��[  � lv%����� �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OWW�# �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_olO ~Od+No`oro�o�o�o �o�o�o�o&8 J\n������u�  0�"0g�/ �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q�����$o�� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E����� Do��������ҿ��� ��,�>�P�b�tφ� �Ϫϼ���������w
�  58�J�\�n� �ߒߜկ��������� 	��-�?�Q�c�u��8���� ��- ����� �2�D�V�h� z�������������������& ���%	1234�5678�" 	��/� `r�������� (:L^p� ������ // $/6/H/Z/l/~/��/ �/�/�/�/�/? ?2? D?V?h?�/�?�?�?�? �?�?�?
OO.O@Oo? dOvO�O�O�O�O�O�O �O__*_YON_`_r_ �_�_�_�_�_�_�_o oC_8oJo\ono�o�o �o�o�o�o�oo" 4FXj|���������	��s�3�E�W�{�Cz�  Bp��   ���2���z�$�SCR_GRP �1�(�U8(ӿ\x^ �@  �	!�	 ׃��� "�$� ��-��+���R�w����D~�����#����O����M-10iAo 8909905 �Ŗ5 M61C �>4��Jׁ
� ���0�����#�1�	"�z�����h��¯Ҭ ��� c���O�8�J�� �����!�����ֿ.��B�y����������A��$�  @��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ�� ��������%��I�4� m��<�l߃ߕߧ���B���\����1� �U�@�R��v��� ��������;���*<=�
F���?�d��<�>HE����@��:��� B����ЗЙ���EL_�DEFAULT � �����B�MIPO�WERFL  ��$1 WFDO� $��ERV�ENT 1������"�pL!DUM_EIP���8��j!AF_�INE �=�!�FT���!���4 ��[!�RPC_MAI�N\>�J�nV�ISw=���!7TP�PU��	�d�?/!
PMON_PROXY@/��e./�/"Y/�f�z/�/!RDM_'SRV�/�	g�/#?G!R C?�h?�o?!
pM�/�i�^?�?!RLSY3NC�?8�8�?O�!ROS�.L�4�?SO"wO�#DOVO �O�O�O�O�O_�O1_ �OU__._@_�_d_v_ �_�_�_�_o�_?oo�coiICE_KL� ?%y (%�SVCPRG1@ho8��e���o�m3�oD�o�`4 �`5(D-�`6PU�`7x }�`���l9��{�d:?��a�o��a �oE��a�om��a�� �aB���aj叟a� ��a�5��a�]��a ����a3����a[�՟ �a�����a��%��aӏ M��a��u��a#����a K�ů�as���a��mo b�`�o�`8�}�w��� ����ɿ���ؿ��� 5�G�2�k�VϏ�zϳ� �����������1�� U�@�y�dߝ߯ߚ��� ��������?�*�Q� u�`��������� ���;�&�_�J��� n�����������sj_DEV y	��MC:(w!`OUT"�,REC �1�Z� d   	 	�������

 �Z�{0H6l Z�~����� � //D/2/h/z/\/ �/�/�/�/�/�/�/? �/,?R?@?v?d?�?�? �?�?�?�?�?OO(O NO<OrOTOfO�O�O�O �O�O�O_&__J_8_ Z_\_n_�_�_�_�_�_ �_�_"ooFo4oVo|o ^o�o�o�o�o�o�o�o 0TBxf� ���(���,� �P�>�`���h����� ����Ώ��(�:�� ^�L���p�������ܟ ���� �6�$�Z�H� ~���r�����دƯ� ���2��&�h�V��� z�����Կ�ȿ
��� ��.�d�RψϚ�|� �Ϭ���������<� �`�N�pߖ߄ߺߨ� ��������8�&�\��J�l��jV 1��w Pl�	}� � �F��
TYPEVF�ZN_CFG ��x�d�7�GRP 1��A�c ,B� A�� D;� B����  B4�RB21HEKLL:�(
� X����%RSR����E0i T�x�������/Sew_�  ��%w������#������A�2�#�d����HK 1��� ���m/ h/z/�/�/�/�/�/�/ �/
??E?@?R?d?�?��?�?�?��OMM �����?��FTOV_ENB ���+��HOW_REG_�UIO��IMWA�ITB�JKOU�T;F��LITIM�;E���OVAL|[OMC_UNITC��F+�MON_AL�IAS ?e�9 ( he�s_(_ :_L_^_��_�_�_�_ �_j_�_�_oo+o�_ Ooaoso�o�oBo�o�o �o�o�o'9K] n����t� ��#�5��Y�k�}� ����L�ŏ׏���� ��1�C�U�g������ ����ӟ~���	��-� ?��c�u�������V� ϯ������;�M� _�q��������˿ݿ ����%�7�I���m� ϑϣϵ�`������� ߺ�3�E�W�i�{�&� �߱������ߒ��� /�A�S���w���� X����������=� O�a�s���0������� ������'9K] ����b�� �#�GYk} �:������ /1/C/U/ /f/�/�/ �/�/l/�/�/	??-? �/Q?c?u?�?�?D?�? �?�?�?O�?)O;OMO _O
O�O�O�O�O�OvO��O__%_7_�C�$�SMON_DEF�PRO ����`Q �*SYSTEM*  d=OU�RECALL ?�}`Y ( �}�6copy fr�s:orderf�il.dat v�irt:\tem�p\=>192.�168.4�P46:3892>_�_�_vo}.�V*.d�_��^�_`oro�oe
x�yzrate 61 +o=oOo�o�oe�g�o�a�o�oc�u�b4�Rmd:�prgst�`.d�g�o�]U��
� �}3�uconslog�� �e�w����io�<�N�ߏ���f2�uerr?all.ls���_pՏf�x��� }9�_~�Xmpback<�pR���
� }0�t%b(`*��ǟ џb��t���c�_�_=�8736 W������o ��˩ϯ`�r����o�o ;�M�޿��'д ��ҿc�uχϚ���5� ͧ�������"���̨���b�t߆ߙtx��:\)ߪ�;�S�U�����.
� }5��a�ߺ� Φ��g�y��ϰ�9� T�����	�߷�@��� c�u�����-�?����� ������N�_q ����1����� �&��J�[m�� ��7�����" �F�i/{/����+/�=/O/�/�/?�)�8504 *?�/c?u? �?��567�?�?�? "�?58�?bOtO�O𙯫?��R�2164 WO�O�O�O��O�I �O`_r_�_�/��;_M_ �_�_o?'?�T�_�_ couo�o�?�?5O�G�o �o�oO"O�o�H�ob t���/�/QcU� �
�/��Nq�h� z���o�o:���� 
���Aӏd�v�������$SNPX_�ASG 1��������� P 0 '�%R[1]@1�.1����?���% ֟��&�	��\�?� f���u��������ϯ ��"��F�)�;�|�_� ������ֿ��˿�� �B�%�f�I�[Ϝ�� ���ϵ�������,�� 6�b�E߆�i�{߼ߟ� ����������L�/� V��e������� �����6��+�l�O� v��������������� 2V9K�o ������� &R5vYk�� ���/��<// F/r/U/�/y/�/�/�/ �/?�/&?	??\??? f?�?u?�?�?�?�?�? �?"OOFO)O;O|O_O �O�O�O�O�O�O_�O _B_%_f_I_[_�__ �_�_�_�_�_�_,oo 6oboEo�oio{o�o�o �o�o�o�oL/ V�e����� ���6��+�l�O��v�������PARAoM �����_ �	��P�����OFT_�KB_CFG  �ヱ���PIN_�SIM  ����C�U�g�����RV�QSTP_DSB�,�򂣟����SR� �/�� & � ULTIROBOTTASK������TOP_O�N_ERR  ����PTN �/�@��A	�RING_P�RM� ��VD�T_GRP 1�<ˉ�  	���� ��������Я���� �*�Q�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߣߠ߲����� ������0�B�i�f� x������������ �/�,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZ�~���� ���/ /G/D/V/ h/z/�/�/�/�/�/�/ ?
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_�8___\_��VPRG�_COUNT�q�@���RENBU��UM�S��__UP�D 1�/�8  
s_�oo*oSo No`oro�o�o�o�o�o �o�o+&8Js n������� ��"�K�F�X�j��� ������ۏ֏���#� �0�B�k�f�x����� ����ҟ������C� >�P�b���������ӯ�ί�����UYS�DEBUG�P�P��)�d�YH�SP_PwASS�UB?Z��LOG ��U��S)�#�0� � ��Q)�
MC�:\��6���_MPAC���U���Qñ�8� �Q�SAV ������ǲ&��ηSV;�TEM�_TIME 1���[ (m��&�����}YT1SVGgUNS�P�U'�U����ASK_OPTION�P�U�Q�Q���BCCFG 3��[u� n�A�a�`a�gZo��� �ߕ��߹������� :�%�^�p�[���� ������ �����6�!� Z�E�~�i���������&�������&8�� nY�}�?�� ԫ ��(L :p^����� ��/ /6/$/F/l/ Z/�/~/�/�/�/�/�/ �/�/2?8 F?X?v? �?�??�?�?�?�?�? O*O<O
O`ONO�OrO �O�O�O�O�O_�O&_ _J_8_n_\_~_�_�_ �_�_�_�_o�_ o"o 4ojoXo�oD?�o�o�o �o�oxo.TB x��j���� ����,�b�P��� t�����Ώ��ޏ�� (��L�:�p�^����� ��ʟ��o��6� H�Z�؟~�l������� د���ʯ ��D�2� h�V�x�z���¿��� Կ
���.��>�d�R� ��vϬϚ��Ͼ����� ��*��N��f�xߖ� �ߺ�8��������� 8�J�\�*��n��� ���������"��F� 4�j�X���|������� ������0@B T�x�d���� �>,Ntb ������/� (//8/:/L/�/p/�/ �/�/�/�/�/�/$?? H?6?l?Z?�?~?�?�? �?�?�?O�&O8OVO hOzO�?�O�O�O�O�O �O
__�O@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<o^o�oro �o�o�o�o�o�o  J8n$O��� ��X���4�"��X�B�v��$TBC�SG_GRP 2��B�� � �v� 
 ?�  ������׏ �������1��U�g��z���ƈ�d,� ���?v�	 H�C��d�>�����e�CL  B�p��Пܘ������\)��Y  A��ܟ$�B�g�B�Bl�i�X�ɼ���X��  D	J���r�����C����үܬ	���D�@v�=�W�j� }�H�Z���ſ���������v�	�V3.00��	�m61c�	*`X�P�u�g�p�>���2v�(:�� ��p���  O�����p�����z�JCFG� �B��� �����������=��=�c�q� K�qߗ߂߻ߦ����� ���'��$�]�H�� l������������ #��G�2�k�V���z� ������������ �p*<N���l� ������#5 GY}h��� �v�b��>�// / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?d? R?t?v?�?�?�?�?�? O�?*OO:O`ONO�O rO�O�O��O�O�O_ &__J_8_n_\_�_�_ �_�_�_�_�_�_�_o Fo4ojo|o�o�oZo�o �o�o�o�o�oB0 fT�x���� ���,��P�>�`� b�t�����Ώ����� ��&�L��Od�v��� 2�����ȟʟܟ� � 6�$�Z�l�~���N��� ��دƯ�� �2�� B�h�V���z�����Կ ¿����.��R�@� v�dϚψϪ��Ͼ��� ����<�*�L�N�`� �߄ߺߨ����ߚ�� �����\�J��n�� ���������"��� 2�X�F�|�j������� ��������.T Bxf����� ��>,bP �t�����/ �(//8/:/L/�/�� �/�/�/h/�/�/�/$? ?H?6?l?Z?�?�?�? �?�?�?�?O�?ODO VOhO"O4O�O�O�O�O �O�O
_�O_@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<oro`o �o�o�o�o�o�o�o &�/>P�/�� �������4� F�X��(���|����� ֏����Ə0��@� B�T���x�����ҟ�� ����,��P�>�t� b������������� ��:�(�^�L�n��� ����2d�����̿ �$�Z�H�~�lϢϐ� �������Ϻ� ��0� 2�D�zߌߞ߰�j��� �������
�,�.�@� v�d��������� ����<�*�`�N��� r������������� &J\�t�� B������ F4j|��^����/�  2 6# 6&J/6"��$TBJOP_�GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� ƞ6$ @2 �"	� �C�� �&b�  Cق'�!�!>ǌ��
559>��0+1�33=��CL� fff?>+0?�ffB� J1��%Y?d7�.��/>;��2\)?0��5���;��h{CY� �  @� ~�!B�  A�P?��?�3EC�  D��!�,�0*BO���?�3JB��
:�/��Bl�0��0�$��1�?O6!Aə�3AДC�1D�G6Ǌ=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__<�O�O>B�\JU�O�HH�1ts�A@g33@?1� C�� ��@�_�_&_8_>��D�UV_0�LP�Q30O<{�zR� @�0 �V�P!o3o�_<oRifo Po^o�o�o�oRo�o�o �o�oM(�ol��p~��p4�6&��q5	V3.0}0�#m61c�$�*(��$1!6�A�� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�IR�CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;S@;Q�U�|8�`rz@/&�8�6&<��1��w�^$ESTPAR�S  *({ _#H�R��ABLE 1%�p+Z�6#|�Q�Q � 1�|�|�|��5'=!|�	|�
|��|�˕6!|�|�:|���RDI��z!ʟܟ� ��$���O������¯ԯ�����S��x# V���˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���U-����ĜP�9� K�]�o��-�?�Q�c��u���6�NUM  ��z!� �>  Ȑ����_CF�G �����!@�b IMEBF_T�T����x#��a�VE�R��b�w�a�R {1�p+
 (3�6"1 ��  6!�� �������� �9�$�:� H�Z�l�~���������@������^$��_���@x�
b MI_�CHANm� x� >kDBGLV;0o��x�a!n ETHE�RAD ?�
� �y�$"�\&�n ROUT��!�p*!*�SN�MASK�x#�255.h�fx�^$OOLOFS_�DI��[ՠ	OR�QCTRL � p+;/���/+/=/ O/a/s/�/�/�/�/�/���/�/�/!?��PE?_DETAI���PON_SVOF�F�33P_MON� �H�v�2-9S�TRTCHK ����42VTCOMPATa8�24�:0FPROG �%�%MULTIROBOTTOx!O06�PLAY���L:_INST_M�P GL7YDUS8���?�2LCK�LPKQUICKMEt ��O�2SCRE�@}�
tps�@�2�A�@�I��@_Y����9�	SR_GR�P 1�� ���\�l_zZg_@�_�_�_�_�_�^�^� oj�Q'ODo/ohoSe ��oo�o�o�o�o�o �o!WE{i�������	1234567�h�!���X�E1�V[�
 �}ipn�l/a�gen.htmno��������ȏ�~�Panel� setup̌}��?��0�B�T�f� ��񏞟��ԟ� ��o����@�R�d�v� �����#�Я���� �*���ϯůr����� ����̿C��g��&� 8�J�\�n�����϶� ��������uϣϙ�F� X�j�|ߎߠ����;� ������0�B��*N�UALRMb@G ?�� [��� ���������� ��%� C�I�z�m�������v�SEV  �����t�ECFG CՁ=]/BaA$�   B�/D
 ��/C�Wi{� ������4 PRց; �To�\o�I�6?K0(%����0���� �//;/&/L/q/\/`�/�/�/l�D ��Q�/I_�@HIS�T 1ׁ9  �(  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1 Ec0p?�?�?�?/C�� >?P=962 n?�?
OO.O�?�?�136c?|O�O�O�OAO SO�?�O__0_�O�O _Lu_�_�_�_:_�/�_ �_oo)o;o�__oqo �o�o�o�oHo�o�o%7I~��a81�o u������o� ��)�;�M��q��� ������ˏZ�l��� %�7�I�[������� ��ǟٟh����!�3� E�W����������ï կ�v���/�A�S� e�Pb������ѿ� �����+�=�O�a�s� ϗϩϻ�������� ��'�9�K�]�o߁�� �߷��������ߎ�#� 5�G�Y�k�}���� �����������1�C� U�g�y���v������� ����	�?Qc u��(���� )�M_q� ��6���// %/�I/[/m//�/�/ �/D/�/�/�/?!?3? �/W?i?{?�?�?�?�� ���?�?OO/OAOD? eOwO�O�O�O�ONO`O �O__+_=_O_�Os_ �_�_�_�_�_\_�_o o'o9oKo�_�_�o�o �o�o�o�ojo�o# 5GY�o}�������?��$UI�_PANEDAT�A 1������  	�}�0�B�T�f�x��� )����mt� ۏ����#�5���Y� @�}���v�����ן�� �����1��U�g�N�\����� �1�� Ïȯگ����"�u� F���X�|�������Ŀ ֿ=������0�T� ;�x�_ϜϮϕ��Ϲ� �����,ߟ�M�� j�o߁ߓߥ߷���� ��`��#�5�G�Y�k� �ߏ���������� ����C�*�g�y�`� ��������F�X�	 -?Qc����߫ ����~; "_F��|�� ���/�7/I/0/ m/�����/�/�/�/�/ �/P/!?3?�W?i?{? �?�?�??�?�?�?O �?/OOSOeOLO�OpO �O�O�O�O�O_z/�/ J?O_a_s_�_�_�_�O �_@?�_oo'o9oKo �_oo�oho�o�o�o�o �o�o�o#
GY@ }d��&_8_�� ��1�C��g��_�� ������ӏ���^�� �?�&�c�u�\����� ��ϟ���ڟ�)�� M�����������˯ ݯ0�����7�I�[� m����������ٿ� ҿ���3�E�,�i�P� �ϟφ��Ϫ���Z�l�}���1�C�U�g�y���)߰�#�������  ��$�6��Z�A�~� e�w��������� ��2��V�h�O������v�p��$UI_P�ANELINK �1�v� � �  ���}1234567890����	 -?G ���o�� ���a��#5G�	����p&���  R��� ��Z��$/6/H/ Z/l/~//�/�/�/�/ �/�/�/
?2?D?V?h? z??$?�?�?�?�?�? 
O�?.O@OROdOvO�O  O�O�O�O�O�O_�O �O<_N_`_r_�_�_�0,���_�X�_�_�_  o2ooVohoKo�ooo �o�o�o�o�o�o� �,>r}����� �������/� A�S�e�w�������� я���tv�z��� �=�O�a�s������� 0S��ӟ���	��-� ��Q�c�u�������:� ϯ����)���M� _�q���������H�ݿ ���%�7�ƿ[�m� ϑϣϵ�D������� �!�3�Eߴ_i�{�
 �߂����߸������ /��S�e�H���~� ��R~'�'�a��:� L�^�p����������� ���� ��6HZ l~���#�5�� � 2D��hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?�/�?�?�?�? �?�?m?OO&O8OJO \O�?�O�O�O�O�O�O �O[�_��4_F_)_j_ |___�_�_�_�_�_�_ o�_0ooTofo��o ��o��o�o�o ,>1bt��� �K����(�:� ���{O������ʏ ܏�uO�$�6�H�Z� l���������Ɵ؟� ���� �2�D�V�h�z� 	�����¯ԯ����� �.�@�R�d�v���� ����п���ϕ�*� <�N�`�rτ��O�Ϻ� Io���������8�J� -�n߀�cߤ߇����� �����o1�oX��o |����������� ��0�B�T�f���� ����������S�e�w� ,>Pbt��' �����: L^p��#�� �� //$/�H/Z/ l/~/�/�/1/�/�/�/ �/? ?�/D?V?h?z? �?�?�???�?�?�?
O O.O��ROdO�߈OkO �O�O�O�O�O�O_�O <_N_1_r_�_g_�_7O�M�m�$UI�_QUICKME�N  ���_AobRESTORE 1��  ��|��Rto�o�im �o�o�o�o�o: L^p�%��� ���o����Z� l�~�����E�Ə؏� ��� �ÏD�V�h�z� ��7�������/���
� �.�@��d�v����� ��O�Я�����ß ͯ7�I���m������� ̿޿����&�8�J� �nπϒϤ϶�a��� ����Y�"�4�F�X�j� ߎߠ߲������ߋ����0�B�T�gSC�RE`?#m�u1sco`uU2��3��4��5��6��7��8��bUGSERq�v��Tp঑�ks����4��5*��6��7��8��`�NDO_CFG ��#k  n` �`PDATE ����Non�ebSEUFRA_ME  �TA��n�RTOL_AB�RTy�l��ENB�����GRP 1��ci/aCz  A�����Q�� $�6HRd��`U������MSK  ������Nv�%��U�%���bVI�SCAND_MA�X�I��FAIL_IMG� ��PݗP#��IM�REGNUM�
�,[SIZ�n`��A�,VONT�MOU��@����2��a���a����F�R:\ � �MC:\�\wLOG�B@F� !�'/!+/O/�U�z MCV��8#UD1r&E�X{+�S�PPO�64_��0'f�n6PO��LI�b�*�#V���,�f@�'�/� =	��(SZV�.�����'WAI�/ST�AT ����P@/�?�?�:$�?�?���2DWP  ���P G@+b=���� H�O_�JMPERR 1��#k
  �23�45678901 dF�ψO{O�O�O�O�O �O_�O*__N_A_S_x�_
� MLOWc>8
 �_TI�=��'MPHASOE  ��F��P�SHIFT�15 9�]@<�\� Do�U#oIo�oYoko�o �o�o�o�o�o�o6 lCU�y�� ��� ��	�V�-��e2����	VSwFT1�2	V�M�� �5�1G� ����%A�  BU8̀̀�@ pك�Ӂ˂�у��z�ME�@�?�{��!c>&+%�aM1��k�0��{ �$`0TDI�NEND��\�O � �z����S��w���P���ϜRELE�Q��Y���\�?_ACTIV��<:�R�A ��e���e�:�RD� ���YBOX �9��د�6��02����190.0m.�83���254��QF�	� �X�j��1�robot����   px�૿�5pc�� ̿�����7�����-�^f�ZABC�����,]@U��2ʿ�eϢ� �ϛϭϿ����� �� �V�=�z�a�s߰�E�	Z��1�Ѧ