��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 � �1��(�|UREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8GW�+0�$Y $DB\� 6COMW!2�MO� "0�A.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6*_�7_�8_�94F;CO�$ <� �o��o�hK3 1#`O_M|c@AC t � �E#6NGPvABA� �c1�Q8��`,���@nr1�� d�P��0e���axnp�UP&Pb26���p�"J��p_R�rPBC��J�rĘߜJV�@U� B���s}�g1�"YtP_�*0OFS&R @�� RO_K8T��aIyT�3T�NOM_�0��1p�34 >��DC �� Ќ@��hPV���mEX�p� �0g0xۤ�p�r
$TF��2C$MD3i�TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F�"F��40CP@�a2 6�@$�PPU�3N�)ύRևA�X�!DU��AI�3BUF�F=�@1� |pp���pPIZT� PP�M��M�y��F�SIMQSI�"ܢVAڤrT�=�w T�`�(zM��P�B�qFAkCTb�@EW�`P1�BTv?�MC�� �$*1JB8`p�*1DEC��F���ŤA��� ��H0CHNS_EMP1�$G��8��@!_4�3�p|@P��3�TCc�(r/�0-sx� �ܐ� MBi��!�����JR� i�SEGF�R��Iv �aR�TrpN�C��PVF��|?�bx &� �f{uJc!�Ja��� !2�8�ץ�AJ���SIZ�3S�c�B�TM���g�|��JaRSINFȑ b���q�۽�н�����L�3�B���CRC�e�3CCp��� �c��mcҞb�1J�c�P��.����D$ICb�Cq�5r�ե��@v�'����EV���zF��_J��F,pN��ܫ��?�4�0A�! � r���h�Ϩ��p�2��͕a�� �د�R>�Dx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�=M��CUR��Q�UA1  $@TITO1/S@S�!�����"0�DBPXWO���B0!5�$SKL���FDBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z���LB�)$�/���� %�/��$C�!&?�$ENE�q.'*?�Ú �RE�p2(H ���O�0#$L|3$$�#�B[�;�К�FO_D��ROSr�#������3�RIGGER�6P�ApS����ETUR�N�2�cMR_8�T�Uw��0EWM��M�GN�P���B#LAH�<E���P��O&$P� �'P@D�Q3�CkD{��DQฑ�4�11��FGO_oAWAY�BMO����Q#!�DCS�_�)  �PIS� I gb {s�C��A��[ �B$�S���AbP�@�EW-�TNTVճ�BV�Q.�C� (c`�UWr�P�J��P�<$0��SAFE���V�_SV�bEXCL�U��nONL�2��SY�*a&�OT<�a'�HI_V�'��(�D���_ *�P0� 9�_z��p ����ASG�� +nrr�@6Acc*b���G�#@E�V.iHb?fA�NNUN$0.$fdI%D�U�2�SC@�`��i�a��j�f�"�pO�GI$2,O�$F�ibW$}�OT9@�1� $DUMMY T��da��dn�� � ��E- ` ͑HE4(sg�*b�SAB���SUFFIW�V�@CA=�c5�g�6r �DMS�W�E. 8Q�KE3YI5���TM�10s��qA�vIN����D���/ D��HOST_P!�rT��t�a��tn��tsp�pEMpӰV��� SBLc �ULI�0  p8	=ȳ���DTk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&Q�DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F��!df�J� �ј�PC1�+6 H�bLL_DUs�~a3@{��3:���OTX"����s�r�0NOAUT5O�!7�p$)�$�*��c4�(�Cy�R8�C, �""�L�� 8H *8�LH <6����c"�` , `Ĭ�kª�q��q���sq��~q��7��8J��9��0����1��U1̺1ٺ1�1�U1 �1�1�2(ʩ2����2̺2ٺ2��2�2 �2�2*�3(�3��3��̺U3ٺ3�3�3 �U3�3�4(ʡ8T�?��!9 <�9�&�z��I��1���M��O�FE@'@� : y,6��Q? �@FP?9��5�9�E�@A�r���A� �;p$TP�$VARI:�ፂ6@P2�P< ���TDe���K`Q�縡�- ��BAC�"=# T�p��e$)_,�b8n�kp+ IFIG�kp��H  ��P����PF@`�!>t� ;E��sC�ST�D� D���c�<� 	C��{��_����l���R  ���F?ORCEUP?b���FLUS�`H�N�>�F ���RD_CM�@E������ ��@v\MP��REMr F�Q���1k@���7Q
Kr4	NJ�5EFFۓ�:�@IN2Q��OV�O�OVA�	TR3OV���DTՀ�DTMX� ��@ �
ے_PH"p��CL��_TpE�@�p2K	_(�Y_T��v*(��@A;QD� ������!0tܑ0RQ���_�a����M�7�CL�dρR�IV'�{��EAR6ۑIOHPC�@��2��B�B��CM9@����R �GCLF�e!DYk(M�ap#5TuDG��� ̑%/�SSD �s? �P�a�!�1���P_(�!�(�!1��E�3�!�3�+5�&�GRA���7�@��;�PW泅ONn��EBU�G_SD2HP�{�_/E A`��_�TERM`5Bi5���ORI#:e0C�9SM_�P��re0Di5�p�TA�9�Ei5�0UP\�F�� -�A{�A�dPw3S@B$SEG��:� EL{UUSE.�@NFIJ�B$��;1젎4�4C$UFlP=�$,�|QR@"��_G90Tk�D��~SNST�PATx����APTHJ��E�p%B`�'EC���AR$P�I�aSHFTy�A�A�H_SHORР꣦6% �0$�7PE��E�GOVR=��aPI�@��U�b �QAYLOW���IE"�r�A8��?���ERV��XQ �Y��mG>@�BN��U\��R2!P.uA�SYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC����EP;�uP;�6WOR�>@M`�!�GRSM5T6�G3�GR��13�aPAL@��P��q�u_H � ���'TOCA�`P	P�`$OP����pѡ�`0O��R%E�`R4C�AO�p��Be�`R�Eu�h|�A��e$PWR�3IMu�RR_�cN�\�q=B I&2H���p_ADDR��H_LENG�B�q�qT�q$�R��S�JڢSS��SKN��u\�0�u̳�uٳSE�A�n���HS��MN�!K�����b����OLX��p����`ACRO3pJ�@���X�+��Q��6�OSUP3�b_�IX��a�a1��}򚃳��� (��H��D��ٰ��X氋�IO2S鐁D������`�7��L $d��`Y!_O�FFr�PRM_���"�HTTP_�+�H:�M (|pOcBJ]"�p��$���LE~Cd���N � ��֑AB_�TqᶔS�`H�LVh�KR"uH�ITCOU��BG�LO�q���h�`����`��`SS� ����HW�#A:�O�ڠ<`INCPU>2VISIOW�͑���n��to��to�ٲ ��IOLN��P �8��R��p$S�Lob PUT_&n�$p��P& ¢���Y F_AS�"Q��$L������Q"  U�0	P4A��50��ZPHY��-��x���UOI �#R ` �K����$�u�"pPpk���$���,��a�UJ5�S-���;NE6WJOGKG̲'DIS���Kp���&�#T (�uAVF�+`��CTR�C
�FL�AG2�LG�dU� ���؜�13LG_SIZ����b�4�Xa��a�FDl�I`� w� m�_�{0a�^��c g���4�����Ǝ���x{0��� SCH_���a7�N�9�VW����E�"����4��U�M�Aљ`LJ�@�DAUf�EAU�p��d|Ҧr�GH�bĠ���B�OO��WL ?�6 IT�����wREC��SCR �ܓ�D
�\���MARGm�!��զ ��dH%�����S����W���U� �JGM[�M�NCHJ���FNK�EY\�K��PRGƂ�UF��7P��FW�D��HL��STP���V��=@��А�RES��HO`����C9T@��b ��7�[�UL����6�(RD� ����Gt��@PO��������MD�FOCU��RwGEX��TUI��	I��4�@�L� ����P����`���P��NE��CANAx��Bj�VAILI��CL !�UDCS_CHII4��s�O�D(!�S���S��灴 ��BUFF��!X�?PTH$m���v`��a���AtrY�?P��j�\3��`OS1Z2Z�3Z8�� Z � ��[aEȤ��Ȥ�IDX�dPSRrO����zA�STL�R�}�Y&�� Y$E�C���K�&�&z�� [ L Q��+00�	P���`#q�dt
�U�dw<���_ \ ?�4Г�\���Ѩ#\0C4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#b�D���'B�LD�%�$�%ORGڰ5�2��PVŇVY8�s�T�r�#}d^ ���$6��$�%S�`T� �B0��4�6RCLMC��4]?o?�9세�MI��p}d_ d=њR�Q��DSTB��p� ;F�HHA�X�R JHdLEXGCESra�BM!p�a`�/B�T�F��`5a�p=F_A7Ji���KbOtH� K�db q\Q���v$MBC��LI|�)SREQU�IR�R�a.\o�AXD�EBUZ� �MLt M��c�b�{Ph����2ANDRф�`�`d;�2�ȺSDC��N�INl�K�x`��X� N&��aZ�����RPST� �ezrLOC�RYIrp�EX<fA�px�9AAODAQ��7f XY�OND�rMF,Łf�s"��`}%�e/� ���FX3@�IGG�� g ��t"��ܓs#N�s$R�a%��iL��h�L�v�@�DATA#?pE�%�jq��Y��Nh t $+MD`qI}�)nv� ytq�ytHP`�Pxu��<(�zsANSW)�yt(@��yuD+�)\b��ܵ0o�i �@CU�w�V�p 0XeRR2��j Du�{Q��7B?d$CALIA@���G��2��RIN���"�<��INTE��Ck�r^�آXXb]���_N�qlk����9�D���Bm��DIVFDH�@���qnI$V,��S�;$��$Z�X��o�*����o�H �$BELT|�u!ACCEL�q.�~�=�IRC��� ���D�T�8�$SPS�@�"L��Ѐr��#^�S�Eы T�P�ATH3���I���3x�p�A_W��ڐ���2nC��4�_MG�$DD��T���$FW�Rp9���I�4��DE7�PP�ABN��ROTS�PEE�[g�� J���[�C@4���$OUSE_+�VPi�F�SYY���1 q�YN!@A�ǦOF�F�qǡMOU��N�G���OL����INC�tMa6��HB�<�0HBENCS+�8q`9Bp�4�FDm�IN��Ix�]��B��VE���#�y�23_UP�񕋳LOWL� ��p� B���Du�9B #P`�x ���BCv�r��MOSI��BMO�U��@�7PERCH  ȳOV��â
� �����D�ScF� @MP����� Vݡ�@y�j�LUk��Gj�p��UP=ó���ĶTR�K��AYLOA �Qe��A��x�����N`�F�RTI�A$��MOUІ�HB�BS0�p7D5���ë�Z��DUM2ԓS_BCKLSH_Cx� k����ϣ���=���ޡ �	ACLAL�"q��1м@��CH�K� �S�RTY@��^�%E1Qq_�N޴_UM�@�C#���SCL0�r�LM?T_J1_L��9@H�qU�EO�p�b�p_�e�k�e�SPC�0�u���N�PC�N�!Hz \P��C�0~"sXT��CN_:�1N9��I�SF!�?�V���U�/���x�T�2��CB!�SH�:� �E�E1T�T����y����T��PA ��_	P��_� =�����P�!����J6 L�@���OG�G�TO7RQU��ONֹ���E�R��H�E�g_W2���_郅����I�I�I��F�f`xJ�1�~1�VEC3�0BD:B�1p�@SBJRK�F9�0DBL_S�M��2M�P_DL2GRV������fH_��d����COS���LNH������@��!*,�aZ����fMY�_(�T�H��)THET0��NK23���"郶�CB�&CB�C AA�B�"��!��!�&�SB� 2�%GTS�Ar�CIMa������,4#97#$DU ���H\1� �:Bk62�r:AQ(rSf$NE�D��`I��B+5��$̀�!A�%�5�7���LPH�E�2���2SC%C%�2-&PFC0JM&̀V�8V�8T߀LVJV!KV/KUV=KVKKVYKVgIH�8FRM��#X!KUH/KH=KHKKHYKUHgIO�<O�8O�Y�NOJO!KO/KO�=KOKKOYKOM&F��2�!+i%0d�7SP�BALANCE_lo![cLE0H_�%SPc� &�b&�b&PFULC�h�b�gخb%p�1k%�UT�O_��T1T2�i/�2N��"�{�t�#�Ѱ`�0�*�.�T��OÀ<�v INSsEG"�ͱREV4v�Ͱl�DIF�ŕ�1�lzw��1m��OB0pq�я?�MI{���~nLCHWARY��_�AB��!�$MECH�!o ��q�AX��P����7Ђ�`n 
�d(�U�7ROB��CRr�H����s(�MSK�_f`�p P 
�`_��R/�k�z�����1S�~�|�z�{����z��qINUq�M?TCOM_C� �q  ���pO�?$NOREn��y��pЂr 8p �GRe�uSD�0A�B�$XYZ_�DA�1a���DEBaUUq������s z`�$��COD�� �L���p�$BUFINDX|�w  <�MORm�/t $فUA��ր����r�<��rG���u � $SIMUL  S�*�Y�<̑a�OBJE�`̖�ADJUS�ݐA'Y_IS�D�3�܎��_FI�=��Tu 7�~�6�'��p@} =�C�}p�@b�D���FRIr��T��RIO@ \�E}'�y��OPWOYq�v}0Y�SYSBU/@v�$SOPġd����ϪUΫ}pPRUN,����PA��D���r\ɡL�_OUo��q�$)�IMA�G��w��0P_qIM��L�INv�K�?RGOVRDt�梄X�(�P*�J�|��0L�_�`]��0�RB�1�0��M��E�D}��p ��N�PMdֲ��Uc�w�SL�`�q�w x $OwVSL4vSDI��DEX����#�$��-�V} *�N4�\@#�B�2�G�B�_�M��x� �q�E� �x Hw��p��AT+USW���C�0o��s���BTM�ǌ�I
�k�4��x�԰q�y Dw�E&���@E�r��7��жЗ�EXE��ἱ���8��f q�z @w���3UP'��$�pQ�XN����������� �PG΅{ h? $SUB�����0_���!�MPW�AIv�P7ã�LO�R�٠F\p˕$R�CVFAIL_C��٠BWD΁�v��DEFSP!p | Lw���Я�\���UNI+�����bH�R�+�}_L\p�P�� �P��p�}H�> �*�j��(�s`~�N�`KET�B�%�J�PE Ѓ~z��J0SIZE�����X�'���S�OR~��FORMAT�``��c ��WrEM�t��%�UX��G����LI��p�  �$ˀP_SWI��pq�J_PL��A�L_ �����AR��B��� C��D��$E��.�C�_�U�� � �� ���*�J3xK0����TIA4��u5��6��MOM��@������ˀB�ЃAD����������PU� NR��������m��� A$PI�6q��	� ����K4�)6��U��w`��SPEEDgPG������� �Ի�4T�� � 8@��SAMr`��p\�]��MOV_� _$�npt5��5���	1���2��������Ȣ'�S�Hp�IN �'�@�+�����4($4+T+GAMM�Wf�1'�$GETH`�p���Da���

pOLIBR>�II2�$HI=�_g�t��2�&E;��(A�.� �&LW�-6<�)56�&�]��v�p��V��?$PDCK���q"��_?�����q� &���7��4���9+�� �$IM_SR�pD�s�rF��r&�rLE���Om0H]��0�y��pq���PJqUR_S�CRN�FA���S_?SAVE_D��dE@�NOa�CAA�b� d@�$q�Z�Iǡs	�I � �J�K� ����H� L��>�"hq��� ���ɢ�� bW^U�S�A�2CM4� ��a��)q`��3�WW� I@v�_�q�3AMUAo��� � $PY�+�$W�P�vNG�{��P:��RA��RH��RO�PL�����qP� ��s'�X;�OI��&�Zxe ���m�� p��ˀ�3s�O�O��O�O�O�aa�_т� |��q�d@��.v��.v��d@��[wFv��E����%s�t;B�w�t|�tP���PMA��QUa ��Q�8��1٠QTH�H{OLW�QHYS��3ES��qUE�pZB���Oτ�  ـP�ܐ(�A����v�!�t�O`�q��u�"���8FA��IROG�����Q2���o�"��p�^�INFOҁ�׃hV����R�2AOI���� (�0SLEQ ������Y�3����Á��P0Ow0��5�!E0NU���AUT�A�COPAY�=�/�'��@Mg��N��=�}1������ ���RG��Á���X_�P�$;ख�`
��W��P��@��������EXT_CY�C b2A��RpÁ��r��_NAe!�А���ROv`	��� � ���P�OR_�1�E2�SReV �)_�I�DI��T_�k�}�'���dШ������5��6��7���8i�ME�PS�dB���2�$��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,��0FL`�o@YN���K�M��Ck��P�WR+�9ᘐ��D�ELA}�dY�pA�D�a� �QSK;IP4� �A�$�-OB`NT�} ��P_$�M�ƷF@\bIp ݷ�ݷ�ݷd���� 빸��Š�Ҡ�ߠz�9��J2R� n��� 4V�EX� TQQ����TQ������� ��`�#�RDCN�V� �`��X)�R�p�����r��m$�RGEAR_� I9OBT�2FLG��fi&pER�DTC����|����2TH2NS�}� 1���G: T\0 ���uЉM\Ѫ`I�d"�R�EF�1Á� l<�h��ENAB��cTPE�04�]���� Y�]��ъQn#��*��"P�������2�Қ��@����������3���'�9�K�]�o���4�Ҝ������������5�ҝ!�3�E�PW�i�{��6�Ҟ��@�����������7���-?Qcu�8�Ҡ��������SMSKÁ��l��a��EkA��M�OTE6����`�@�݂TQ�IO}5R�IS�tR�W@��� �pJ�����p����E�"$DSB_SIGN�1�UQ�x�C\�TPC_S�RS232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+�TQ��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�P%��S�0�����p�_XPE +�$FREEFROMS	p�na�GET�0��U�PD�A�2��SP|� :��� !$USAN�na&����ERI�0�Rp�RYq5*"_j@�P8m1�!�6WRK9K�D���6��QFRIgEND�Q�RUFg��҃�0TOOL�6M�Y�t$LENG�TH_VT\�FI!R�pC�@ˀE> +IOUFIN-RM���RGI�1ÐAIT�I�$GXñ3IvFG2v7G1���p3�BơGPR�p�1F�O_0n 0��!RE��p�53҅U�TC��3A�A��F �G(��":���e1n!��J�8�%����%]��%�� 74�OX O0�L��T�3H&��8���%b4J53GE�W�0�WsR�TD����T��M�����Q�T]�$V C2����1�а91�8��02�;2k3�;3 �:ifa�9-i�aQ���NS��ZR$V��2BVwEV�2AUQ�B;�����&�S�`��F`�"�k�@�2a�PS�E��$r1C��_g$Aܠ6wPR��7vMU�cS�t '�/8�9�� 0G�aV`��p�d`���50�@���-�
25S�� E��aRW����B��&�N�AX�!�A�:@LAh��rTHI�C�1I���X�d1T�FEj��q�uIF_CH�3�qI܇7�Q�pG1RxV���]�岺:�u�_JF~�P�RԀƱ�RVAT��� ��`���0�RҦ�DOfE��CO9UԱ��AXI����OFFSE׆TRIGNS���c����h����H�Y��IGGMA0PA�pJ��E�ORG_UNE9V�J� �S����?�d �$CА�=J�GROU�����TOށ�!��DSP���JOGӐ�#��_	Pӱ�"O�q����@n�&KEP�IR��dܔ�@M}R��AP�Q�^�Eh0��K�SY�S�q"K�PG2�B�RK�B��߄�p`Y�=�d����`AD_�<����BSOC����N��DUMMY1�4�p@SV�PDE�_OP�#SFSP_D_OVR-���1C��ˢΓOR٧3�N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1q"�LCHDL��REGCOVʤc0��Wq@1M������RO�#��rȐ_+��� @0��e@VER�$O�FSe@CV/ �2WD�}��Z2����TR�!���E_�FDO�MB_CiM���B��BL�bܒ#��adtVQR�$0�p���G$�7�AM�5��� eŤ��_M�;��"'����8$C�A��'�E�8�8$HcBK(1���IO<�q����QPPA�ʀ����
��Ŋ����DVC_DBhC;�� #"<Ѝ�r!S�1[ڤ��S�3[֪�ATIO"q 1q� ʡU�3���CABŐ�2�CvP ��9P^�B���_� �?SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW�_C��U��S@��SA��A�pl$UNITm�l_�AT���e��ƐCYCLq�NE�CA���FLTR_2_FIO�7(�ӌ)&B�LPқ/�.�_�SCT�CF_`�F0b�l���|�FS(!E�e�CHA�1��4�D��"3�RSD��$"}�����_Tb�PR�O����� EMi_䙰a�8!�a �!�a��DIR0�R�AILACI�)RM�r�LO��C���Q`q��#q�դ�PR=�%S�AC/�c =	��FUNCq�0rRINP�Q�0��2f�!RAC �B ��p[���[WARn�F��BL�Aq�A����DAk�\���LD0���Q�d�qeq�TI"rp��K�hPRIA�!r"AF��P@!=�;@��?,`�RK���Mǀ9I�!�DF_@B�l%1n�LM�FAq@OHRDY�4_�P@�RS�A�0� �MU�LSE@���aG ��ưt��m��$�1$�1$�1o����� x*�EG00�����!AR���Ӧ�09p�2,%� 7�AXE���ROB��WpA��_l-��SY[�W!‎&MS�'WRU�/-1��@�STR������Eb� 	�%��J��AB� ���&9�����kOTo0 	$��ARY�s#2��Ԓ��	ёFI@��$�LINK|�qC1��a_�#���%kqj2XYZ��t;rq�3��C1j2^8'0B��'�4����+ �3FI���7�q����'��_Jˑ���O3�Q'OP_�$;5���A#TBA�QBC��&��DUβ�&6��TURN߁"r�E11:�p��9GFL�`_���* Ȩ@�5�*7��Ʊ +1�� KŐM��&�8���"r��ORQ��a�(@#p=� j�g�#qXU�����mT'OVEtQ:�M��i�@��U��U��VW�Z �A�Wb��T{�, ��@ ;�uQ���P\�i��UuQ��We�e�SERʑe	��E� O���UdAas��4S�/7����AX��B� 'q��E1�e��i��i rp�jJ@�j�@�j�@�j P�j@ �j�!�f��i ��i��i��i��i �y�y�'y�7y�TqHyDEBU8�$32���qͲf2G + AB����رnS9VS�7� 
#�d� �L�#�L��1W��1W� JAW��AW��AW�QW��@!E@?D2�3LAB�29U4�Aӏ��Co  o�ERf�>5� � $�@_ mA��!�PO���à�0#�
�_MR}At�� d � 9T��ٔERR����;TY&���I��V8�0�cz�TOQ�d�PL[ �d�"�� ?�w��! � pp`T8)0���_V1Vr�a(Ӕ����2ٛ2�E�ĺ��@�H�E���$QW�����V!��$�P��o�cI��a�Σ	 HELL_�CFG!� }5��B_BASq��SR3��� �a#Sb���1�%���2��3��4��5*��6��7��8����RO����I0�0NL��\CAB+�����ACK4�����,�\@2@��&�?�_PU�CYO. U�OUG�P~ �����m�������TPհ_KAR�l�_�RE*��P���7QUE���uP�����CSTOPI_AL7�l�k0��h��]��l0SEM�4�(�Ml4�6�TYN�SO���DIZ�~�A������m_TM�MAN�RQ��k0E�����$KEYSWIT�CH���m���HE���BEAT��EF- LE~�����U���F!Ĳ���B�O_H�OM=OGREFUPPR&��y!� [��C��O��-ECO�C��Ԯ0_IOCMxWD
�a�%(k��� � Dh1���	UX���M�βgPgC�FORC��� 챒m�OM.  �� @�5(�U�#P�, 1��, 3��4�5��NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�� �� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E��VP���UPDs� � �`NЦ�5�YS�LOt�� � �L��d���A�aTAp�0d��|�ALU:eLd�~�CUѰjgF!a�ID_L�ÑeHI��jI��$FILE1_���d��$2�f;SA>�� hO��`?E_BLCK��b|$��hD_CPUy�M�yA��c�o�d��Y�����R �Đ
�PW��!� oqL�A��S=�ts�q~tRUN�qst�q~t����qst�q~t �TACCs���X -$�qLEN@;��tH��ph�_�I���ǀLOW_AXI��F1�q�d2*�M Z���ă��W�Im�ւ�aR�TOR��pg��D�Y���LACE�k�ւ�pV�ւ~�_M�A2�v�������TCV��؁��T��ي������t�V����V�J$j�R�MA�i�J��m�Ru�b����q2j�`#�U�{�t�K�JK��CVK;���H���3���J0����JJ��JJ��AAL��ڐ���ڐԖ4Օ5���NA1���ʋƀW�LP��_(�g����pr��� `�`GROU�w`��B��NFL�IC��f�REQUwIRE3�EBU�0�qB���w�2����p����q5�p�� \^��APPR��C}��Y�
ްEN٨CL9O7��S_M��H����u�
�qu�� ���MC�����9�'_MG��C�Co��`pM�в�N�BRKL�GNOL|�N�[�R���_LINђ�|�=�J����Pܔ�������� ���������6ɵ��̲8k�D����G� ��
��q)�<�7�PATH3�L�@B�L��H�wࡠ�J�CN�CA�Ғ�ڢ6B�IN�rUCV�4aZ��C!�UM��Y,���aE�p����������PAYLOAJ2L`R_A	N�q�Lpp����$�M�R_F2LS3HR��N�LOԡ��Rׯ�`ׯ�ACRL�_G�ŒЛ� ��H�j`߂$HM���FWLEXܣ�qJ�u� :���� ���������1�F1�V�j�@�R�d�v�������E����ȏ ڏ����"�4�q��� 6�M���~��U�g�y�$ယT��o�X��H� �����藕?����� ǟِݕ�ԕ�����%�7��P��J�� �� V�h�z���`A�T�採@�EL�� �S��J|�Ŝ�J�Ey�CTR��~�T�N��FQ��HAN/D_VB-���v`n�� $��F2M����ebSW�b�'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)�F�AW�Z`i�Aw�A���X X�'pi�Dw�Dʆ�Pf�G�p�)ST�k��!x��!N��DY �pנM�9$`%Ц�H� �H�c�׎���0� ��Pѵڵ����������J��� ����1��R�6��QA'SYMvř���v���J���cі�_SH >��ǺĤ�ED����������J�İ%��C��IDِ�_VI��!X�2PV_UNIX�FThP�J��_R�5 _Rc�cTz�pT�V��@�@��İ�߷��U �Ԓ�����Hqpˢ���aEN��`D	I����O4d�`J��� x g"IJAA ȱz�aabp�coc�`a��pdq�a� ��OMME��� �b�RqT(`PT�@� S��a7�;�Ƞ�@�h�a��iT�@<� $�DUMMY9Q�o$PS_��RFC�v�$v � 8���Pa� XƠ����STE���SB}RY�M21_VF�8$SV_ERF�qO��LsdsCLRJtEA��Odb`O�p� � D $�GLOBj�_LO ���u�q�cAp�r�@awSYS�qADR`�`�`TCH  �� ,��ɩb�W_NA���7�Ac��TSR���l ���
*?�& Q�0"?�;'?�I)?�Y) ��X���h���x����� �)��Ռ�Ӷ�;��Í�v�?��O�O�O�D�XOSCRE栘p�����ST��s}Hy`����/_H�A�q� TơgpTYP�b���G�a�G���Od0IS�_䓀d��UE�Md� ����ppS<�qaRSM_�q*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCOUx��S�Ԕ 1�!��UE&��Ubwr��PoROGM�FL@o$CUgpPO�Q\���UI_�`H�� � 8�� �_�HE�PS�#��`RY ?�qp�b�t�dp�OUS��� � @6p�v_$BUTTp�Rp>R�COLUMq�e���SERV5�P�ANEH�q� �; �@GEU����Fy��)$HELyPõ)BETERv�)ෆ���A � � ��0��0��0ҰSIN簪c�@N���IH�1��_� �֪�LN�rؓ �qpձ_ò=�s$H��TEXl�����FLA@��RELV��D`����j����M��?,�Š��m����"�U�SRVIEW�q�S <6p�`U�`��NFI@;�FOC�U��;�PRI@�m�`�QY�TRIP>�qm�UN<`Md�� #@p�*eWA�RN)e�SRTO�L%��g��ᴰO�NCORN��RAU䘠��T���w�VI�N�Le� $�גPATH9�גCwACH��LOG�!�LIMKR����v����HOST��!�b�R��OB�OT�d�IM>� �� ���Zq��Zq;�VCPU_A�VAIL�!�EX
	�!AN���q��10r��1r��1M�ѡ�.�p�  #`C����@$TOOL��$��_JMP� ����e$SS�����VSHIF��Nc�P�`ג��E�ȐR����OSU�R��Wk`RADILѮ��_�a��:�9a���`a�r��LULQ�$OUTPUT_3BM����IM�ABp �@�rTIL'SCO��C7� ������&��3 ��A���q���m�I�2G�o�y@Md��}��yDJU��N_�WAIT֖�}Ҵ�{�%! NE�u��YBO�� ��� $`�t�S�B@TPE��NE�Cp�J^FY�nB_T��R�І�a$�H[YĭcB��dM� ��F� �p�$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"�`�"��[���P?� �ZABC~%��  $�"�R��
ϐ�$$C�LAS�������!ϐ� � � VI�RT]��/ 0ABS�����1 5�� < �!F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZi{0�-�AXL�pl��!�n63  �{tIN��qztPRE�����v��p�uLARMRECOV 9l�rwtNG�� .;	 A   �|.�0PPLIC���?5�p��Handlin�gTool o� �
V7.50P�/23-�  �P�f��
��_S�Wt� UP�!�� x�F0��t���A�� v� 86-4�� �it�y�� r2 �7DA5�� ��� Qf@<ϐo�Noneisͅ�˰ ��T����!LAex>�_l�V�uT��s9�UTO�"�Њt��y��HGAPON�
0g�1��Uh�D [1581�����̟ޟry����Q 1���p�,� 蘦���;�@��q_���"�" �c�.�H���D�HTTHKYX� �"�-�?�Q���ɯۯ 5����#�A�G�Y�k� }�������ſ׿1��� ��=�C�U�g�yϋ� �ϯ�����-���	�� 9�?�Q�c�u߇ߙ߫� ����)�����5�;� M�_�q������� %�����1�7�I�[� m����������!�� ��-3EWi{ ������ )/ASew�� ��/��/%/+/ =/O/a/s/�/�/�/�/ ?�/�/?!?'?9?K? ]?o?�?�?�?�?O�?��?�?O#O]���TO��E�W�DO_CL�EAN��7��CNMw  � ��__/_A_S_�DS�PDRYR�O��H	Ic��M@�O�_�_�_ �_oo+o=oOoaoso��o�o���pB��v �u���aX�t������>9�PLUGG���G\��U�PRCvPB�@E��_�orOr�_7�SEGF}�K [mwxq�O�O���p��?rqLAP�_ �~q�[�m�������� Ǐُ����!�3�x�TOTAL�f yx�_USENU�p��� �H���B��RG_�STRING 1�u�
�M�n�S5�
ȑ_I�TEM1Җ  n 5�� ��$�6�H�Z� l�~�������Ưد����� �2�D�I�/O SIGNA�L̕Tryout Modeӕ�Inp��Sim�ulatedב�Out��OV�ERR�P = 1�00֒In c�ycl��בProg Abor���ב��Statu�sՓ	Heart�beatїMH� Faul��Aler'�W�E�W�iπ{ύϟϱ������� �CΛ�A����8� J�\�n߀ߒߤ߶��� �������"�4�F�X�8j�|���WOR{pΛ ��(ߎ����� ��$� 6�H�Z�l�~���������������� 2PƠ�X ��A{ ������� /ASew��p���SDEV[ �o�#/5/G/Y/k/ }/�/�/�/�/�/�/�/�??1?C?U?g?y?PALTݠ1��z? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�Op�O�O_�?GRI�` ΛDQ�?_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o2_l�R��a\_�o" 4FXj|��� ������0�B�<T��oPREG�>��  f���Ə؏����  �2�D�V�h�z��������ԟ���Z��$�ARG_��D ?�	���;���  	�$Z�	[O�]�O��Z�p�.�SBN�_CONFIG S;��������CII_SAVE  Z�����.��TCELLSET�UP ;�%HOME_IOZ�~Z�%MOV_��
�REP�lU�(�UTOBACKܠ���FRwA:\z� \�,z�Ǡ'`�z���\ǡi�INI�0z����n�MESS�AG���ǡC���ODE_D������%��O�4�n�PAUS�X!�;� ((O>��ϞˈϾϬ� ���������*�`߀N߄�rߨ߶�g�l TSK  wͥ�_��q�UPDT+��d�!�A�WSM_C5F��;���'�>-�GRP 2:�?�+ N�BŰA��%��XSCRD1�1
N7� �ĥĢ�� ��������*����� ��r�����������7� ��[�&8J\n���*�t�GROU�N�UϩUP_N5A�:�	t���_ED�17�
� �%-BCKEDT-�2�'K&�`���-t��z�q�q�z����2t1������q�k�(/��ED3/��/�.a/�/;/M/ED4�/t/)?��/.?p?�/�/ED5`??�?<?.�?O�?�?ED6O�?qO��?.MO�O'O9OED7�O`O_�O.�O\_�O�OED8L_,�_�^-�_ oo_�_�ED9�_�_]o�_	`-9o�oo%oCR _ 9]�oF�o�k�� � NO_DEL���GE_UNU�SE��LAL_?OUT �����WD_ABOR�ﰨ~��pITR_�RTN��|NO�NSk���˥C�AM_PARAM� 1;�!�
 8�
SONY X�C-56 234�567890 �ਡ@���?}��( А\��
���{����^�H�R5q�̹��ŏR5y7ڏ�Aff���KOWA SC�310M
�x��>��d @<�
� ��e�^��П\�� ��*�<��`�r�g��CE_RIA_I��!�=�F���}�z� ��_LeIU�]������<��FB�GP 1.��Ǯ�M�x_�q�0�C*  ��V��C1��9��@��iG���CR�C]��Ud��l��s��R��T���[Դm��v���������� C����(�����=�{HE�`ONFIǰ��B�G_PRI 1�{V���ߖπ�Ϻ����������C�HKPAUS�� ;1K� ,!uD� V�@�z�dߞ߈ߚ��� �������.��R�<�hb���O���������_MOR��� ���<�y����� 	 �� ���*��N�`����"���?��q?;�;�I���K��9�P����ça�- :���	�

��M����pU�ð��<��,,~��DB���튒�)
mc:cpm�idbg�f�:_�  5&'¥��p�/�  ����̟���� �s>�(���(��U�?�u�w�[g�/� 
� �f�M/w�O/~�
DEF l���s)�< buf.txts/�t/��ާ�)�	`���Λ�=L�T�'MC��1����?43���1��t�īC�z  BHH�CP�UeB�^&B����;��>C�?��CnY
K��E?{hDS��D���?r���D���D��^��=Fǁ,F�M�\F���Cm	�fF��F����:���'w�1�T��s���.�p�������BDw�M@x�8��1Ҩ����g@D��p@�0EY�1X��EQ�EJ�P F�E�F�� G��>^�F E�� FB�� H,- Ge���H3Y��:��  >�33 s���~  n8�~@��5Y�E>�ðyA��Y<#�
"Q� ���+_�'RS/MOFS�p�.8���)T1��DE ���F 
Q��;�(P  B_<_���R����	o�C4RP�Y
s@ ]AQ��2s@C�0B3�MaCR{@@*cw��UT�p�FPROG %�z�o�oigI�q���v���ldKEY_TB�L  �&S�#� ��	
�� �!"#$%&'(�)*+,-./0�1i�:;<=>?�@ABC� GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�������������������s���p`LCK�lx4�p`�`STAT ���S_AUTO_D�O���5�IND�T_ENB!���R��Q?�1�T2}�^�S�TOPb���TRL^r`LETE��Ċ�_SCREEN ��Zkcs�c��U��MMEN�U 1 �Y  <�l�oR�Y1� [���v�m���̟���� �ٟ�8��!�G��� W�i��������ïկ ��4���j�A�S��� w�����迿�ѿ��� �T�+�=�cϜ�sυ� �ϩϻ�������P� '�9߆�]�o߼ߓߥ� �������:��#�p� G�Y��������� ��$����3�l�C�U� ��y����������� ���	VY)�_MA�NUAL��t�DB;CO[�RIGڇ
��DBNUM� ���B1 e
�PXWO_RK 1!�[�_�U/4FX�_�AWAY�i�G�CP  b=�Pj_CAL� #�j�Y���܅ `�_�  1"��[ , 
�@od�&/~&lMZ��IdPx@P@#ON�TIMه� dɼ`&�
�e�MO�TNEND�o�R�ECORD 1(��[g2�/{�O� �!�/ky"?4?F?X? �(`?�?�/�??�?�? �?�?�?)O�?MO�?qO �O�O�OBO�O:O�O^O _%_7_I_�Om_�O�_  _�_�_�_�_Z_o~_ 3o�_Woio{o�o�_�o  o�oDo�o/�o S�oL�o���� @���+�yV,� c�u��������Ϗ>� P�����;�&���q� ��򏧟��P�ȟ�^� �����I�[�����  ���$�6��������jTOLEREN�CwB���L��͖ CS_CFG� )�/'d�MC:\U�L%0?4d.CSV�� �c��/#A ��CH
��z� //.ɿ���(S�RC_OUT� *���S�GN +��"���#�10-FE�B-20 17:�32015-JA�Np�0:51+? P/Vt�ɞ��/.��f�pa�m��PJPѲ���VERSION� Y�V2�.0.84,EFLOGIC 1,�/ 	:ޠ=��ޠL��PROG_�ENB��"p�UL�Sk' ����_WRSTJNK ��"�fEMO_OPT?_SL ?	�#�
 	R575/#=�����0�B�|���TO  ��صϗ��V_F EX�d�%��PAT�H AY�A\p�����5+ICT�-Fu-�j�#�egS�,�STBF_TTS�(@�	d���l#!w�� �MAU��z�^"MS%WX�.��<4,#�
Y�/�
!J�6�%ZI~m��$SBL_FAUL(�y0�9'TDIA[��1<�� ����1234567G890
��P�� HZl~���� ���/ /2/D/V/hh/�� P� ѩ�yƽ/��6�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�,�/�UMP���� �ATR���1OC@�PMEl�OOY_T�EMP?�È�3pF���G�|DUNI���.�YN_BRK �2_�/�EMGDI_STA��]��E�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�a�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��aDzr�A W�_BWD�p��xf�́t�_DI�� 9�5�d�T�asRֆSTEP��:P��OP_DOv��f�PFACTOR_Y_TUNwdM��EATURE �:�5̀rQ�Handling�Tool �� \�sfmEng�lish Dictionary���roduAA� Vis�� Ma�ster����
�EN̐nalog� I/O����g.�fd̐uto S�oftware �Update  �F OR�mat�ic Backu�p��H596�,�ground �Editޒ  1� H5Cam�era�F��OP;LGX�ell𜩐�II) X�omm�Րshw���com揭co���\tp����pane�� � opl��tyl�e select^��al C��nJ�~Ցonitor��gRDE��tr��?Reliab𠧒�6U�Diagno�s(�푥�552�8�u��heck �Safety U�IF��Enhan�ced Rob �Serv%�q )� "S�r�UserG Fr[�����a���xt. DIO 6�fiG� sŢ��wendx�Err�MLF� pȐĳr�r�� ����  !���FCTN Men�u`�v-�ݡ���T�P Inېfac��  ER J�GC�pבk E�xct�g��H55�8��igh-Sp�ex�Ski1�  �2
P��?���m�munic'�on1s��&�l�ur�ې���ST Ǡ��c�onn��2��TX�PL��ncr�s�tru����"FA�TKAREL Cmd. LE�{uaG�545\�ſRun-Ti��E{nv��d
!����ؠ++�s)�S/�W��[�Lic�enseZ��� 4�T�0�ogBook�(Syڐm)��H�54O�MACRO�s,\�/Offs�e��Loa�MH�������r, k�M�echStop �Prot���� l�ic/�MiвSh�if����ɒMixpx��)���xStS��Mode Swiwtch�� R5W��Mo�:�.�� 7#4 ���g��K��2h�ulti-T�=�M���LN (�Pos�Reg�iڑ������d�ݐtO Fun�ǩ�.�����Num~����Ï lne��ᝰ Adjup������  - W��ta�tuw᧒T��RDMz�ot��s�cove U�9����3Ѓ�uesOt 492�*�o������62;�SNP�X b ���8 Jy7`���Libr��FJ�48���ӗ� ����
�6O�� Pa�rts in VCCMt�32���x	�{Ѥ�J990��{/I� 2 P���TMILIB��Ht���P�AccD��L�
TE$TX܍ۨ�ap1S�Te<����pkey���wգ�d��Un�exceptx�motnZ��������3є�� O��΄� 90J�єSP CSXC<�f�l�Ҟ� Py�We}�Β�PRI�>vr\�t�men�� ��/iPɰa������vGrid�play��v��0�)��H1�M-10iA(B201 ��2\� 0\k/�A/scii�l�Т��ɐ/�Col��ԑG7uar� 
�� /�P-�ޠ"K��stN{Pat ��!S��Cyc�҂�or�ie��IF8�ata- quҐ�� ƶ���mH574��RML��am���Pb�HMI De3�(�b����PCϺ�P�asswo+!��"PE? Sp$�[���stp��� ven���Tw�N�p�YEL?LOW BOE	k$wArc��vis���3*�n0WeldW�cial�7�V#Mt�Op����1y�֠ 2F�a�pocrtN�(�p�T1�`T� �� ��xy]ֹ&TX��tw�ig�j�1� b� ct\��JPN ARC?PSU PR��ovݲOL� Sup�2fil� &PAɰא�cro�� "PM�(����O$SS� enвtex�� r����=�t�ssag$T��P��P@�Ȱ�锱�rtW��H'�>r�dpn��n1#
t�!� z ���ascbin4p�syn��+Aj�M� HEL�NCL� VIS PKG�S PLOA`�McB �,�4VW��RIPE GET_VAR FIEo 3\t��FL[��OOL: ADD� R729.FD/ \j8'�CsQ�Q�E��DVvQ�sQNO WTWTE��>}PD  �^��b�iRFOR ��EC�Tn�`��ALSE� ALAfPCPM�O-130  M�" #h�D: H�ANG FROM�mP�AQfr��R7�09 DRAM �AVAILCHE�CKSO!��sQVP�CS SU�@LIMCHK Q +P~d�FF POS��F��Q R593�8-12 CHA�RY�0�PROGR�A W�SAVE�N`AME�P.SV2��7��$En*��p�?FU�{�TRC|� �SHADV0UPD�AT KCJўRS�TATI�`�P M�UCH y�1��I�MQ MOTN-�003��}�ROB�OGUIDE DAUGH�a���*�Gtou����I� Š�hd�ATH�PepM�OVET�ǔVM�XPACK MA�Y ASSERT��D��YCLfqTA��rBE COR �vr*Q3rAN�pR�C OPTION�SJ1vr̐PSH�-171Z@x�tcǠSU1�1Hp^9R!�Q�`_T�P��'��j�d{tby app wa 5IҌ~d�PHI���p�aT�EL�MXSPD' TB5bLu 1��U�B6@�qENJ`CEV2�61��p��s	�may n�0� �R6{�R� �Rtr�aff)�� 40�*�p��fr��sy�svar scr� J7��cj`DJ�U��bH V��Q/��PSET ERR�`J` 68��PN�DANT SCR�EEN UNRE�A��'�J`D�pPA��pR`IO 1����PFI�pB�pG/ROUN�PD��G���R�P�QnRSVIP� !p�a�PDIGI?T VERS�r}B�Lo�UEWϕ P�06  �!��MA�Gp�abZV�DIx�`� SSUE��ܰ�EPLAN {JOT` DEL�p�ݡ#Z�@D͐CAsLLOb�Q ph���R�QIPND��I{MG�R719���MNT/�PES ��pVL�c��Holp�0Cq���tPG:�`:C�M�canΠ���pg.v�S: 3�D mK�view� d�` �p��eat7У�b� of �P�y���ANNOT �ACCESS M���Ɓ*�t4s a��lok��Fle�x/:�Rw!mo?�PA?�-�����`~n�pa SNBPJ AUTO-�0�6f����TB��PIA�BLE1q 636>��PLN: RG$��pl;pNWFMD�B�VI���tWIT� 9x�0@o��Qu�i#0�ҺPN RR�S?pUSB�� t� & removb�@ )�_��&AxEP7FT_=� 7<`�p�P:�OS-14;4 ��h s�g���@OST� � C�RASH DU �9��$P�pW�� .$��LOGI�N��8&�J��6b0�46 issue� 6 Jg��: �Slow �st~��c (Hos`��c���`IL`IMP�RWtSPOT:Wqh:0�T�STYW =./�VMGR�h��T0CAT��hosB��E�q��� �uO�S:+pRTU' �k�-S� ����E:���pv@�2�� t\�hߐ��m ��al�l��0�  $�H� �WA͐��3 CN�T0 T�� Wr}oU�alarm���0s�d � �0SE1����r R{�OMEpBp���K� 55��REàSEst��g�     �KoANJI�no����INISITA�LIZ-p�dn1we�ρ<��dr�� l�x`�SCII L��fails w��� ��`�YSTE�a���o��Pv� IItH���1W�Gro>P�m ol\wpSh�@�P��Ϡn cfslxL@АWRI ЏOF Lq��p?�F��up��de-r�ela�d "A�Po SY�ch�Ab�etwe:0INDc t0$gbDO����r� `�Gig�E�#operab[ilf  PAbHi�xH`��c�lead�\etf�Ps�r��OS 030�&: f{ig��GLA )P� ��i��7Np t�pswx�B��If��g������5aE>�a EXCE#dU��_�tPCLOS��"�rob�NTdpF�aU�c�!���PNIO V750�Q�1��Qa��DB Ė�P M�+P�QED��DET��-� \�rk��ONLINEhSBUGIQ ߔXĠi`Z�IB�S a�pABC JAR�KYFq� ���0MSIL�`� R�pNД� �p0GAR��D�*pR��P�"! jK�0cT�P�Hl#n��a�ZE V�� TwASK�$VP2(��4`
�!�$�P�`WI[BPK05�!FȐ�B/��BUSY oRUNN�� "��ȁ����R-p�LO��N�DIVY�CU9L��fsfoaBW�p���30	�V��ˠIT`�a5�05.�@OF�UGNEX�P1b�af�@��E��SVEMGN� NMLq� D0pCC_SAFEX �0c�08"qD �PE�T�`N@�#J87�����RsP�A'�M��K�`K�H G�UNCHG۔MEKCH�pMc� T� � y, g@�$ ORY LEAKA8�;�ޢSPEm�Ja:��V�tGRIܱ��@�CTLN�T�Rk�FpepR�j506�EN-`IN������p �`�Ǒk!��Tq3/dqo�STO�0)A�#�L�p �0�@�Q�АY�&�;pb1CTO8pP�s���FB�0@Yp`�`DU��a!O�supk�t4 � PЙF� Bnf�Q�PSVGN-1��V�S'RSR)J�UP��a2�Q�#D�q l �O��QBRKCTR5Ұ�|"-�r�<p�c�j!INVP�D ZO� ��T`h#�Q�cHset,|D��"DUAL� w�2*B�RVO117 A�]�TNѫt�+bTa2�473��q.?��sA�Uz�i�B�comp�lete��604�.� -�`haknc�U� F�Нe8��  ��npJ�tPd!q��`��� 5Nh596p�!5d��� "p�P�P�Q�0�P2@�p�A� xP��R(}\*xPe� aʰI����E��1��p� j � � xSt�^t ��A�AxP�q 5 siug��a��"AC;a���
�bCexPb_p��.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o`�dxP�b]o2�� �c�b�c�ixP�jupf�rm�dxP�o�`ex�e�a�oFdxPtpe�d}o��u`�cptlcibxzxP�lcr�xrxP\�blsazEdxP_fm�}gcxP�x@���o|sp�o�mc(�N�ob_jzop�uD6�wf��t��wms�1q��sld�)��jCmc�o\�n��nuhЌ���|st�e��>�p1l�qp�iwck����uvf0uߒ��lv�isn�Cgacu�lwQ
E F  ;! Fc.fd�Qv��� qw���Dat�a Acquis�i��nF�|1�RR6�31`��TR�QDM�CM �2�P75�H�1�P583xP1���71��59`�5�P57<PxP�Q����¨�(���Q��o p�xP!daq\�o�A��@�� ge/�e�tdms�"DMEsR"؟,�pgdD����.�m���-��qacq.<᡾xPmo��Dh���f{�u�`13���MACROs, Sksaff�@z�����03�SR�Q(��Q6���1�Q9ӡ�R�ZSxh��PxPJ643�@�7ؠ6�P�@�PRS��@���e �Q�UС �PIK�Q52 P�TLC�W��xP3 (��p/O��!�P�n �xP5��03�\sfmnmc "MNMCq�<��Qj��\$AcX�FM�� �ci,Ҥ�X����cd�pq+�
�sk�SKx�xP�SH560�,P��,�y�refp "REFp�d�A��jxP	�of�OF�c�<gy�to�TO�_����ٺ����+je�u��caxi�s2�xPE�\�e�q"�ISDTc��]�porax ��MN�x�u�b�isde܃�h�\�w�xP! is_basic��B�� P]��QAxes��R6������.�(sBa�Q�ess� �xP���2�D�@�z�atis���(�{������~��m��F�Mc�u�{�
ѩ�MNIS��ݝ����x�����ٺ��x� j7}5��Devic��� Interfa�c�RȔQJ7540��� xP�Ne`� �xP�ϐ2�б�����dn� "DNE����
tpdnu�i5UI��ݝ	b�d�bP�q_rs�ofOb
dv_aro��u����>�stchkc���z	 �(}onl��G!ffL+H�@J(��"l"/�n�bx��z�hamp���T�C�!i�a"�59`��S�q��0 (�+�P�o�u�!2��xpc�_2pcchm��C�HMP_�|8бpe�vws��2쳌pc�sF��#C SenxPacro�U·�-�R6�Pd�xPk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GE�M,\i(��Dgesnd�5���H{�}Ha��@sy���c�Isu�xD��Fmd��I��7��4���u���AccuCal�P�4� ��Rɢ7ޠB0��6+56f�6��99\aFF q�S(�U��2�
X�ap�!Bd��cb_��SaUL��  ��� ?�ܖto��ot�plus\tsr�nغ�qb�Wp��t����1��Tool (N. A.)�[K�7�Z�(P�m�����bfcls� k94�"K4p��qt�pap� "PS�9H�stpswo`��p�L7��t\�q ����D�yt5�4�q��@w�q��� �M�uk��rkey����s���}t�sfeatu�6�EA��� cf)t\�Xq�����d�h5���LRC0�md�!�C587���aR�(�����2V��8c?u3l\�pa3}H�&r-��Xu���t,�� �q "�q�Ot��~,���{@�/��1c�}����y�p �r��5���S�XAg��-�y���Wj874��- iRVis<���Queu�� �Ƒ�-�6�1���(����u���tӑ�����
�tpvtsn? "VTSN�3C�t+�� v\pRDV����*�prdq\�Q<�&�vstk=P�������nm&_�դ��clrqν���get�TX��Bd����aoQϿ�0qstr�D[� ��t�p'Z��Ɵ�npv��@�enlIP0��D!x�'�|����sc ߸��tv�o/��2�q���v b����q���!���h�]��(� Con�trol�PRAuX�P5��556�A�@59�P56.@5�6@5A�J69�$@982 J55?2 IDVR7�hq A���16�H���La��� ��Xe�f�rlparm.fn�FRL�am��C9�@(F������w6{���A��QJ6�43�� 50�0L�SE
_pVAR� $SGSYSC���RS_UNIT�S �P�2�4tA�T�X.$VNUM_OLD 5�1�xP�{�50+�"�` Funct���5tA�� }��`#@�`3�a0��cڂ��9���@HA5נ� �P���(�A ����۶}����ֻ}��bPRb�߶~p{pr4�TPSPI0�3�}�r�10�#;A � t�
`���1���96�����%C�� A�ف��J�bIncr �	����\���1o�5qni4�MNINp	xP�`���!���Hour  �� 2�21� �AAVM����0 ��T�UP ��J5�45 ��616�2�VCAM � (�CLI{O ��R6�<N2�MSC "�P �STY�L�C�28~ 13�\�NRE "FwHRM SCH^��DCSU%O�RSR {b�04� �EIOC��1 j 542 �� os| � eg�ist�����7��1�MASmK�934"7 ���OCO ��"3�8��2���� C0 HB��� 4�";39N� Re�� ��LCHK
%OP�LG%��3"%MH�CR.%MC  ; 4l? ��6 dPI�s54�s� DSW%�MD� pQ�K!63!7�0�0p"�1�Р"�4 �6<27 CgTN K � 5 ��%�"7��<25�%/�=T�%FRDM� ��Sg!��930 FB( NBA�P� ( �HLB  Men��SM$@jB( PV3C ��20v��2�HTC�CT�MIL��\@PAC� 16U�hAJ`SA�I \@ELN��<29�s�UECK <�b�@FRM �b�sOR���IPL��}Rk0CSXC ���VVFnaTg@H�TTP �!26� ��G�@ob�IGUI"%IPG�S�r� H863 �qb�!�07r�!34 |�r�84 \so`0! Qx`CC3 Fb�291�!96 rb!g51 ���!53R%� 1!s3!��~�.rp"9js VATFU�J775"��pLR6�^RP�WSMjUCTO�@xT58 F!s80���1XY ta�3!770 ��8�85�UOL  GTS�o
�{` LCM ��r| TSS�EfP6� W�\@CPE �`��0VR� l�QN�L"��@001 i7mrb�c3 =�b0�0���0�`6 w�b^-P- R-�b8n@75EW�b9 �Ґa�� ���b�`ׁ�b2 O2000��`3��`4*5�`5!�c��#$�`7.%�`8 h�605? U0�@B�6E"aRp7� !Pr8 t�a@�tr�2 iB/�1vp3L�vp5 Ȃtr9Σʐa4@-p�r3 	F��r5&�re`u�&�r7 ��r8�U�p9 \h738�a��R2D7"�1�f��2&�7� �3� 7iC��4>w58Ip�Or60 C�L��1bEN�4 I�py�L�uP��@N�-PJ8d�N�8NeN�9 H�(r`�E�b7]�|�⠂8�Вࠂ9 2H��a`0�qЂ5�%?U097 0��@q1�0���1 (�q�3 5R���0 ���mpU��0�0��7*�H@(q�\P"wRB6�q124�b`;��@���@06� 6x�3 pB/x�u ���x�6 H606�a1� ��7 6� ���p�b15�5 ����7jUU1g62 �3 g���4*�65 2ec "_��P�4U1`����B1���`0'�1�74 �q��P�E1�86 R ��P�7� ��P�8&�3 (��90 B/�s1q91����@202��6 3���A�R�U2� d��2 bI2h`��4�᪂2�L4���19v Q�2�*�u2d�Tpt2� ��EH�a2hP�$�5��F�!U2�p�p
�2�p���@5�0-@��84 @�9��TX@�� :�e5�`rb26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0`@�gqGA���a52ѐ��Ḳ6�60ہ5�� ׁ2��8�E��9��EU5@ٰ\�q5�hQ`S�2ޖ5�p\�w�۲�pJ �-P��5��p1\t�H�4��PeCH�7j��phiw��@��P�x��559 ldu� P�D���Q �@������� �`.���P>��8�581l�"�q58�!AM۲�T�A iC�a58�9��@�x����5 �a��12׀0.�1����,�2����,�!P\�h8��Lp ��,�7z��6�0840\� ANRS 0C}A`��p��{��ran���FRA��Д�� ����A%���ѹ�� ������(����Ќ� ��З���������������$�G��1���⨂��������� xS�`q� � �����`64��M���iC/50T-�H������*��)p46��� C��N�����m75s֐� Sp��b46��v��༌ГM-71?�70�З����42�������C��-�а�70H�r�E��/h����O$��rD���c7c7C�q���ą���L��/��2\?imm7c7�g� ������`���(� ��e�����"��������a r��c�T,�Ѿ�"��,�� ��xx�Ex�m77t����k���5�����v)�iC��-HS -� B
_�>���+�Т�7U�]���M*h7�s��7������-9?�/260L_������QB�������]�9p�A/@���q�S��х���h6k21��c��92�������.�)92c 0�g$�@�����)$p��5$���pylH"O"
�21���t?�350����p���$�
�� �350!���0��9�U/�0\m9��M9AA3��4%� s��3M$��X%u���"him98J3����� �i d�"m4~�103�p�� ����h794̂�&R���H�0���� \���g�5AU��՜� �0���*2��00��#06�АՃ���!07{r ����� ���kЙ@����EP�#������?�p�#!�;&07\;!�B1P�߀A��/��CBׂ2�!�:/��?8�ҽCD25L�����0�"l�2BAL
#��B��\20�2 _�r�re���X��1@��N����A@��z��`C�pU��`��#04��DyA�\�`fQ��sU���\��5  ���� p�^t��<$8�5���+P=�ab1l��1LT��lA�8�!uDnE(�20�T��J�1 e�bH8�5���b�Ռ�5[�16Bs��������d�2��x��m6t !`Q����bˀ���b#�(�6iB;S�p�! ��3� ��b�s��-`�_�W8�_���&�6I	$�X5�1�Uc85��R�p6S� ���/�/+q�!�q��`񈓃6o��5m[o)�m�6sW��Q�?��set06p ��3%H�5��10p$����g�/�JrH�� � ��A�856�����F�� ���p/2��h�܅�✐)�5��̑v��(��m6��Y�H�ѝ̑�m�6�Ҝ��a6�DM�����-S�+��H 2�����Ҽ�� �r ̑��✐��l����p1���F���2�\wt6h T6H�� ��Ҝ�'Vl���� ���V7ᜐ/����;3A7��p~S��������4�`圐�V�T��!3��2�PM[�p�%ܖO�chn��vel5����Vq���_arp#��̑�.�~��2l_hemq$8�.�'�6415��� 5���?����F������5g�L�ј[���1���𙋹1����M7NU�М��eʾ����uq$D;��-�!4��3&H�f�c�Ĝ� h������u�� �㜐��ZS�!ܑ4�&��M-����S�$̑�ք �� 0��<������07shJ�H �v�À�sF��S*� ����̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(UL� &�(�,���0�\�?����̑�a�� xS�t���a�e�w�2ȫ�(�	�2�C��A/����\�+p�����2�1 (ܱ�CL S ����B̺��7F��h�?�<�lơ1L� ���c� ���u9�0����e/q��O���98�K��r9 (��,��Rs�ז�5�G�m20c��i��w�A2��:�0`�$��2�2 l�0�k�X�S� ,�ι�2��O���1!4�1w���2T@� _std��G�y� �ң�<H� jdgm���� w0\� �1L���	�P��~�W*�b��t 5P������3�,����E{������LL��5\L��3��L�|#~���~!���4��#��O����h�L6 A�������2璥���44�����[6\j4s��·��@�#��ol�E"w�8P k�����?0xj�H1�1`Rr�>��]�2a�#2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l��0`�&�"��|�`Am1�2@��ػ��3�HqB ��K�R��ˑb�W� ��Fs���)�ѐ�!����a�1����5��16�16C��C<����0\imBQ���d����b��\B5�-���DiL���O�_�<ѠPEtL�E�RH��ZǠPgω�am1l ��u���̑�b�<����<�$�T�̑�F�����Ȋ�Dpb��X"x�ᒢ��p� ����^t��9�0\� �j971\kckrcfJ�F�s������c��e "CTM�E�r�����!�a�`main.[��g�`Grun}�_vc�# 0�w�1Oܕ_u����bctme��Ӧ�`�ܑ�j735�-� KAREL U�se {�U���J���1���p� U ̑�9�B@��L�9����7j[�atk208 "K��Kя��\��9��a��̹�����cKRC�a�o ��kc�qJ�&s��� ��Grſ�fsD��:y�0�s��A1X\j|хr�dtB�, ��`.	v�q�� �sǑIf��Wfj52�TKQu�to Set��J�� H5K536�(�932���91�5�8(�9�BA�1(�7�4O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v���! conre;a�#�Controlw Re�ble��CNRE(�T�<�4��2���D�)���S�55i2��q(g�� (����4X�cOux�\s�futs�UTS `�i�栜���t�棈���? 6�T�!�S#A OO+D6����������,!��6�c+� igt�t6iB��I0�TW8 �0��la��vo58�o�b@Få򬡯i�Xh���!Xk�0Y!8\m6e�!6EC���v��6���������<1!6�A���A�6s��ƀ�U�g�T|ώ���rE1�qR��˔Z4�T������,#�eZp)g ����<ONO0���uJ���tCR;��F�a� �xSt�f��prdsuchk �1���2&&?���t��*D %$�r(�✑�娟:r���'�s�qO��<s�crc�C�\At�trldJ"o�\�V�|���Paylo�nfirm�l�!�87��7��A�3ad�! �?ވI�?hplQ��3��3"�q��x pl�`���d87��l�calC�u�Du���;��movx�����initX�:s8O��a�r4 ���r67A4|�e GeneratiڲĐ��7g2q$��g =R� (Sh��c ,|�bE��$ԒA\�:�"��4���4�4�. sg��5��F$d6"e�!p? "SHAP�T�Q ngcr pGC��a(�&"� ��"G3DA¶��r6�"�aW�/�$dataxX:s�"tpad��<[q�%tput;a__�O7;a�o8�1�yl+s��r�?�:�#�?�5x$�?�:c O�:y O�:H�IO�s`O%g�q�ǒ�?�@0\��"o�j�92;!�Ppl.C�ollis�QSkip#��@5��@J��D ��@\ވ�C@X��7��7�|s2��potcls�LS��DU�k?�\_ et1s�`�< \�Q䜐�@���`dcKqQ�F�C;��J,�n��` (��4eN����T�{���'j(�c�q����/IӸaȁ��̠GH�����зa��e\mcclmt "CLM�/��� �mate\��lmpALM�?>p7qCmc?����2vm�qp��%�3s��_sv90<�_x_msu�2L�^v_� K�o�{in��8(3r<�c_lo�gr��rtrcW� �v_3�~yac��d�<�ten��der$cCe�' Fiρ�R��Q��?�l�enteAr߄|��(Sd��V1�TX�+fK�r�a�99sQ9+�5�r�\tq\� "FN�DR���S�TDn$LAN]G�Pgui��D�`���S������sp�!ğ֙uf�ҝ�s����$�����e+�=�� �������������w�H�r\fn_�ϣ��|$`x�tcpma��- TCP�����?R638 R�Ҭ���38��M7p, ���Ӡ�$Ӡ�8p0Р��VS,�>�tk��99 �a��B3���PզԠ��0D�2�����UI��t� ��hqB���8��������p���re�ȿ��exe@4φ�B���pe38�ԡG�rmpWXφ�var@�φ�@3N�����vx�!ҡ���q�RBT �$cOPTN ask E0��1��R MAS0�H5�93/�96 H5�0�i�480�5�H0��m�Q�K��7�0�g�Pl�h0ԧ�2�ORDP��@"��_t\mas��0�a@��"�ԧ�����k�� �R����ӹ`m��bL��7�.f��u�d���r��splay�D�E���1w�UPD�T Ub��887 M(��Di{���v�� ��Ԛ⧔��#�B���|����o  ��� �a�䣣��60q��B�����qscan0��B���ad@�������q`�䗣��#��К�`2�� vl v��Ù�$�>�b����! S��Easyy/К�Util��|룙�511 J������R7 ��Nor|֠��inc),<6Q�� �`c��"4�[���986FVRx� So����q�nd 6����P��4�a\ (�@�
  �������d���K�bdZ���men�7���- Me`t!yFњ�Fb�0�T�Ua�577?i 3R��\�5�u?��!� n���f���<���l\mh�Ц�pűE|hmn�	���<\O���eD�1�� l!��y��Ù�\|p����B���Ћmh�@��:. aG!���/�t��55�6�!X�l�.u�s��Y/k)ensu)bL���eK�h��  �B\1;5g?y?�?�?D��?*rm�p�?Ktbox O2K|?0�G��C?A%ds���?1ӛ#� �TR��/� �P�4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?�Ă�Q3t.�P׀al���P+OP51�7��IN0a��Q(8}g��PESTf3u�a�PB�l�ig�h�6��aq��P � sxS��`  n��0mbumpP�Q969g�69�Qq��P�0�baAp�@Q� �BOX��,>vchqe�s�>vetu㒼�=wffse�3� ��]�;u`aW��:z#ol�sm<ub�a-��]D�K�ibQ�c���p�Q<twaǂ tp�Q�҄Taror ROecov�b�O�P�642����a�0q��a⁠QErǃ�QCry�з`�P'�T�`��aar������	{'�p�ak971��71���m���>�pjo@t��PXc��C�1�adb� -�ail��na�g���b�QR629��a�Q��b�P  ?�
  �P���$$CL[q O����������$�PS_DI�GIT���"�!�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����*�璬1:PROD�UCT�Q0\PGSTK�bV,n��99�\����$FEAT_I�NDEX��~��� 搠I�LECOMP ;��)��"���SETUP2 �<��� � N !�_AP2BCK 1=�?  �)}6/"E+%,/i/��W/ �/~+/�/O/�/s/�/ ?�/>?�/b?t??�? '?�?�?]?�?�?O(O �?LO�?pO�?}O�O5O �OYO�O _�O$_�OH_ Z_�O~__�_�_C_�_ g_�_�_	o2o�_Vo�_ zo�oo�o?o�o�ouo 
�o.@�od�o� ��M�q�� �<��`�r����%� ��̏[�������!� J�ُn�������3�ȟ W������"���F�X� �|����/���֯e� �����0���T��x� �����=�ҿ�s�π��,ϻ�9�b�� P�/ 2) *.cVRiϳ�!�*�����������PC��7�!�FR6:D"�c��χ��T� �߽�Lը��ܮx���*.F��>� �	N�,�k��ߏ��STM �����Q������!�iPe�ndant Pa'nel���H��F����4������GIF�������u����JPG&P��<�����	PAN?EL1.DT�́������2 �Y�G��
3w�����//�
4�a/�O///��/�
TPEIN�S.XML�/����\�/�/�!Cus�tom Tool�bar?�PA?SSWORD/�?FRS:\R??� %Passw�ord Config�?��?k?�?O H�6O�?ZOlO�?�OO �O�OUO�OyO_�O�O D_�Oh_�Oa_�_-_�_ Q_�_�_�_o�_@oRo �_voo�o)o;o�o_o �o�o�o*�oN�or ��7��m� �&���\����� y���E�ڏi������ 4�ÏX�j�������� A�S��w�����B� џf�������+���O� ��������>�ͯ߯ t����'���ο]�� ���(Ϸ�L�ۿpς� Ϧ�5���Y�k� ߏ� $߳��Z���~�ߢ� ��C���g�����2� ��V����ߌ���?� ����u�
���.�@��� d������)���M��� q�����<��5r �%��[� &�J�n� �3�W���"/ �F/X/�|//�/�/ A/�/e/�/�/�/0?�/ T?�/M?�??�?=?�? �?s?O�?,O>O�?bO �?�OO'O�OKO�OoO �O_�O:_�O^_p_�O �_#_�_�_Y_�_}_o�_�_Ho)f�$FI�LE_DGBCK� 1=��5`��� (� �)
SUMM?ARY.DGRo�\OMD:�o�o
`�Diag Su�mmary�o�Z
CONSLOG�o��o�a
J�aCo�nsole lo�gK�[�`MEMCHECK@'�o��^qMemor?y Data��W߁)�qHADOW���P��s�Shadow ChangesS��-c-��)	F�TP=��9����w�`qmment T�BD׏�W0<�)�ETHERNE�T̏�^�q�Z��a�Ethernet� bpfigura�tion[��P��DCSVRFˏ��Ï�ܟ�q%�� v�erify alylߟ-c1PY���DIFFԟ��̟a���p%��dif!fc���q��1X�?�Q�� ����{X��CHGD��¯ԯi��px��� �¤�2`�G�Y�� 1��� �GD��ʿ�ܿq��p���Ϥ�F�Y3h�O�a��� 1��(�GD���ψ��y��p�ϡ�0��UPDATES.��Ц��[FRS:�\�����aUpd�ates Lis�t���kPSRBW�LD.CM.��\���B��_pPS_R?OBOWEL���_ ����o��,o!�3��� W���{�
�t���@��� d�����/��Se �����N�r � =�a�r �&�J���/ �9/K/�o/��/"/ �/�/X/�/|/�/#?�/ G?�/k?}??�?0?�? �?f?�?�?O�?OUO �?yOO�O�O>O�ObO �O	_�O-_�OQ_c_�O �__�_:_�_�_p_o �_o;o�__o�_�o�o $o�oHo�o�o~o�o 7�o0m�o� � �V�z�!��E� �i�{�
���.�ÏR� ���������.�S�� w������<�џ`��� ���+���O�ޟH��� ���8���߯n����$FILE_��{PR��������� ��MDONLY 1�=4�� 
 ���w�į��诨�ѿ �������+Ϻ�O�޿ sυ�ϩ�8�����n� ߒ�'߶�4�]��ρ� ߥ߷�F���j���� ��5���Y�k��ߏ�� ��B�����x����1� C���g������,��� P���������?���Lu�VISBC�KR�<�a�*.V�D|�4 FR:�\��4 Vi�sion VD file� :L bpZ�#��Y �}/$/�H/�l/ �/�/1/�/�/�/�/ �/ ?�/1?V?�/z?	? �?�???�?c?�?�?�? .O�?ROdOO�OO�O ;O�O�OqO_�O*_<_ �O`_�O�__%_�_��MR_GRP 1�>4�L�UC4�  B�P	 �]�ol`�*u����RHB� ��2 ���� ��� ��� He�Y�Q`orkbIh�o�Jd�o�Sc�o�oM�6�M�D�Kc�F�5U�a�S��0�o�o �E��D�
�(D�#�-����9j>>�}A�uAf��!lq?�W�A�f��xq0~�� F@ �r�d�a}�J��NJk��H9�Hu���F!��IP�s�}?�`�.9��<9�8�96C'6<,6\b�1�,�.�g�R���^x�PA� ����|�ݏx���%� �I�4�F��j����� ǟ���֟��!��E��`r�UBH�P A�~�������W
6��P=��PJ��0˯�o�oB��P5����@�33@���x4�m�,�@UUU���U�~w�>u.�?!x�^��ֿ����3��=[z�=��̽=V6<��=�=�=�$q��~��@8��i7G��8��D�8@9!�7ϥ�@Ϣ����cD�@ D��g Cϫo��C��P��P'�6��_V� m �o��To��xo�ߜo�� ����A�,�e�P�b� ������������ �=�(�a�L���p��� ������^�������* ��N9r]��� �����8# \nY�}���� ���/ԭ//A/� e/P/�/p/�/�/�/�/ �/?�/+??;?a?L? �?p?�?�?�?�?�?�? �?'OOKO6OoO�OH� �Ol��ߐߢ��O�� _ ��G_bOk_V_�_z_�_ �_�_�_�_o�_1oo Uo@oyodovo�o�o�o �o�o�oN u������ ���;�&�_�J��� n�������ݏȏ�� %�7�I�[�"/�描� ����ٟ�������3� �W�B�{�f������� կ�������A�,� e�P�b��������O�O �O��O�OL�_p� :_�����Ϧ������ ��'��7�]�H߁�l� �ߐ��ߴ�������#� �G�2�k�2��Vw� ����������1�� U�@�R���v������� ������-Q� u���r��6� �)M4q\ n������/ �#/I/4/m/X/�/|/ �/�/�/�/�/?ֿ� B?�f?0�BϜ?f��? ���/�?�?�?/OOSO >OwObO�O�O�O�O�O �O�O__=_(_a_L_ ^_�_�_�_���_��o �_o9o$o]oHo�olo �o�o�o�o�o�o�o# G2kV{�h �������C� .�g�y�`��������� �Џ���?�*�c� N���r��������̟ ��)��M�_�&?H? ���?���?�?�?��� �?@�I�4�m�X�j��� ��ǿ���ֿ���� E�0�i�Tύ�xϱϜ� ��������_,��_S� ��w�b߇߭ߘ��߼� ������=�(�:�s� ^��������� �'�9� �]�o���� ~������������� 5 YDV�z� �����1 U@yd��v�� ���/Я*/��
/� u/��/�/�/�/�/�/ �/??;?&?_?J?�? n?�?�?�?�?�?O�? %OOIO4O"�|OBO�O >O�O�O�O�O�O!__ E_0_i_T_�_x_�_�_ �_�_�_o�_/o��?o eowo�oP��oo�o�o �o�o+=$aL �p������ �'��K�6�o�Z�� ����ɏ��폴� � �D�/ /z�D/��h/ ş���ԟ���1�� U�@�R���v�����ӯ ������-��Q�<� u�`���`O�O�O��� ޿��;�&�_�J�o� �πϹϤ�������� %��"�[�F��Fo�� �����ߠo��d�!�� �W�>�{�b���� ����������A�,� >�w�b����������������=��$�FNO ����\��
F0l q  oFLAG>�(R�RM_CHKTY/P  ] ��d ��] ��OM�� _MIN� 	����� �  X�T SSB_CFG� ?\ �����OTP_DEF�_OW  	�|�,IRCOM� �>�$GENOV�RD_DO���<�lTHR� dz�dq_ENB]� qRAVC_?GRP 1@�I X(/ %/7/ /[/B//�/x/�/�/ �/�/�/?�/3??C? i?P?�?t?�?�?�?�? �?OOOAO(OeOLO�^O�OoROU�F\\� �,�|B,�8�?����O�O�O	__��� � DE_�Hy_�\@@m_B�=�vR/��I\�O�SMT�G��SUoo&oRHO7STC�1H�I� ���zMSM��l[bo��	127.0�`1�o  e�o�o�o #z�oFXj|��l60s	anonymous������ao�&�&��o�x��o�� ����ҏ�3��,� >�a�O���������� Ο�U%�7�I��]�� ��f�x��������ү ����+�i�{�P�b� t����������� �S�(�:�L�^ϭ�o� �Ϧϸ������=�� $�6�H�Zߩ���Ϳs� ���������� �2� ��V�h�z��߰��� ������
��k�}ߏ� �ߣ���߬������� ��C�*<Nq�_ ������-�?� Q�c�eJ��n�� �����/"/ E�X/j/|/�/�/� %'/?[0?B? T?f?x?��?�?�?�? �??E/W/,O>OPObO��KDaENT 1I��K P!�?�O  �P�O�O�O�O �O#_�OG_
_S_._|_ �_d_�_�_�_�_o�_ 1o�_ogo*o�oNo�o ro�o�o�o	�o-�o Qu8n��� �����#��L� q�4���X���|�ݏ�� �ď֏7���[����B�QUICC0 ��h�z�۟��1ܟ��ʟ+���2,���{��!ROUTER�|�X�j�˯!PC�JOG̯��!�192.168.�0.10��}GNA�ME !�J!�ROBOT�vNS_CFG 1H�I� �A�uto-star�ted�$FTP�/���/�?޿#?� �&�8�JϏ?nπϒ� ��ǿ��[������"� 4ߵ&����������� �����������'�9� K�]�o������� ������/�/�/G��� k��ߏ����������� ��1T���Py �����"�4�	 H-|�Qcu�V D����/� ;/M/_/q/�/��� �/
/�/>?%?7?I? [?*/?�?�?�?�/�? l?�?O!O3OEO�/�/ �/�/�?�O ?�O�O�O __�?A_S_e_w_�O 4_._�_�_�_�_oVO hOzO�O�_so�O�o�o �o�o�o�_'9 Kno�o����� o*o<oNoP5��oY� k�}�����pŏ׏� ���0���C�U�g�y����_�T_ERR �J;�����PDU�SIZ  ��^�P����>ٕWR�D ?z��� � guest���+�=�O�a��s�*�SCDMNG�RP 2Kz�Ð��۠\���K�� 	P0�1.14 8�q _  y���B    �;����{ �����������������������~ �ǟI�4��m�X�|��  �i  �  k
���� �����+�������_
���l�.x�+���"�l�ڲ۰s�d�������__GROU��L��� ��	��۠0�7K�QUPD  ����PČ�TY�g�����TTP�_AUTH 1M��� <!iP�endan����<�_�!KAR�EL:*������KC%�5�G��V�ISION SE!TZ���|��Ҽ� ����������
�W��.�@��d�v���CTRL N��������
 �,FF�F9E3���F�RS:DEFAU�LT�FAN�UC Web S_erver�
�� ����q��������������WR_CON�FIG O�� ����IDL_�CPU_PC"���B��= �BH�#MIN.�BGNR_IO��� ����% NPT_SI�M_DOs}T�PMODNTOL�s �_PRTY��=!OLNK 1P���'�9K]o�MAS�TEr �����O_gCFG��UO��|��CYCLE����_ASG 19Q���
 q2/ D/V/h/z/�/�/�/�/��/�/�/
??y"N�UM���Q�I�PCH��£RTRY_CN"�u���SCRN������� ���R���?��$J2�3_DSP_EN������0OBP�ROC�3��JO�GV�1S_�@��8�?�';ZO'?}?0CPOSREO~�KANJI_� Ϡu�A#��3T ����E�O�ECL_L�M B2e?�@EYLO�GGIN��������LANGUA�GE _�=�� }Q��LG�2U������ �x������PC � �'0������MC�:\RSCH\0�0\˝LN_DISP V��������TOC�4D�z\A�SOGBOOK W+��o�0��o�o���Xi�o@�o�o�o�o~}	x(y��	ne�i�e�kElG_BUFF� 1X���}2 ����Ӣ���� ��'�T�K�]����� ������ɏۏ����#�P��ËqDCS �Zxm =��� %|d1h`���ʟܟg�IO 1[+# �?'����'�7� I�[�o��������ǯ ٯ����!�3�G�W� i�{�������ÿ׿��El TM  ��d ��#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߈tN�SEV�0m�TYP�� ��$�}�ARS"�(_�s>�2FL 1\��0��������������5�TP<P����DmNGNAMp�4�U�f�UPS`�GI�5�A�5s�_�LOAD@G �%j%@_MO�V�u����MAXUALRMB7�P8��y���3�0]&q��Ca]s�3�~�� t8@=@^+ طv�	��V0+�P�A5d�r���U������ E(iTy�� �����/ /A/ ,/Q/w/b/�/~/�/�/ �/�/�/??)?O?:? s?V?�?�?�?�?�?�? �?O'OOKO.OoOZO lO�O�O�O�O�O�O�O #__G_2_D_}_`_�_ �_�_�_�_�_�_o
o oUo8oyodo�o�o�o��o�o�o�o�o-��D�_LDXDISA�^�� �MEMO_{APX�E ?��
 �0y�����������I�SC 1_�� �O����W�i� ����Ə�����}�� ߏD�/�h�z�a���� ����������@� ��O�a�5��������� ���u��ׯ<�'�`� r�Y������y�޿� ۿ���8Ϲ�G�Y�-� ��}϶ϝ�����m������4��X�j�#�_M?STR `��}տSCD 1as}� R���N��������8� #�5�n�Y��}��� ���������4��X� C�|�g����������� ����	B-Rx c������ �>)bM�q �����/�(/ /L/7/p/[/m/�/�/ �/�/�/�/?�/"?H? 3?l?W?�?{?�?�?�?�n�MKCFG �b���?��LTA�RM_�2cRuB �3WpTN>BpMETPUOp�2�����NDSP_CMNTnE@F��E�� d���N��2A�O�D�EPOS�CF�G�NPST�OL 1e-�4@�<#�
;Q�1;U K_YW7_Y_[_m_�_�_ �_�_�_�_o�_oQo 3oEo�oio{o�o�a�A�SING_CHK�  �MAqODA�Q2CfO�7J�eD�EV 	Rz	�MC:'|HSIZ�En@����eTAS�K %<z%$1�23456789� ��u�gTRIGw 1g�� l<u%���3���>s�vvYPaq��kEM_INF 1h9G� `)�AT&FV0E�0(���)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ���ڄH������G�ֈAO�w�2�������џ ������ ��͏ߏP��t����� ��]�ί�����(� ۟�^��#�5����� k�ܿ� ϻ�ů6�� Z�A�~ϐ�C���g�y� �������2�i�C�h� ό�G߰��ߩ��ߙ� ���������d�v�)� ���߾�y������ ��<�N��r�%�7�I� [������9�&��J[�g��>O�NITOR�@G �?;{   	�EXEC1�3�2*�3�4�5��p��7�8�9�3 �n�R�R�R RRR(R4�R@RLR2Y2�e2q2}2�2��2�2�2�2*�3Y3e3��a�R_GRP_SV� 1it��q(�5�
�3�8��"��۵MO~q_�DCd~�1PL_N�AME !<u�� �!Defa�ult Pers�onality �(from FD�) �4RR2k! �1j)TEX)TsH��!�AX d�? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO@^OpO�O�O�Ox2-? �O�O�O__0_B_T_f_x_�b<�O�_�_�_ �_�_�_o o2oDoVotho&xRj" 1o�)�&0\�b, ��9��b�a @D��  �a?��c�a?x�`�a�aA'�6�e�w;�	l�b	� �xJp��`�`	p� �< ��(p� �.r� K��K ��K=�*�J���J���JV��kq`�q�P�x�|� @j�@T;f�r��f�q�acrs��I�� ��p���p�r�ph}�3���´  ��>���ph�`z��w꜖"�Jm�q� H�N��ac��$��dw��  ��  P� Q� �>� |  а�m��Əi}	'� �� �I� ��  ����:��È�È=����(��#�a	���I�  �n @@H�i~�ab�Ӌ�b�$�w���"N0��  �'Ж�q�p@2��@����r�q5��C�pC0C�@� C����`
��A1]w@B�*V~X�
nwB0h�A��p�ӊ�p@����aDz���֏����Я	�pv�( ?�� -��I�`�-�=��A�a�we�_q�`�p �?�ff ��m��� ����Ƽ�!�1!ݿ�>1�  P�apv(�`ţ� �=��qst��?���`x`�� <
6b�<߈;܍��<�ê<� �<�&P�ό�A�O��c1��ƍ�?ff�f?O�?&��qt@��.�J<?�`��wi4����d ly�e߾g;ߪ�t�� p�[ߔ�߸ߣ������ ����6�wh�F 0%�r�!��߷�1�������E�� E��O�G+� F� !���/���?�e�P���Xt���lyBL�cB�� Enw4�������+�� R��s����x�����h�Ô�>��I�`mXj���A�y�weC��������#/*/c/N/wim�����v/C�`�� CHs/`
=$�p��<!�!��ܼ�'�3�A�A�AR1�AO�^?�$��?���±
�=ç>�����3�W
=�#�\]�;e��?������{����<��>(�B��u��=B�0�������	R��zH�F�G����G��H��U`E���C��+��}I#��I��HD��F��E��R�C�j=�>
�I��@H�!�H�( E<YD0w/O*OONO 9OrO]O�O�O�O�O�O �O�O_�O8_#_\_G_ �_�_}_�_�_�_�_�_ �_"oooXoCo|ogo �o�o�o�o�o�o�o 	B-fQ�u� ������,�� P�b�M���q�����Ώ ���ݏ�(��L�7� p�[������ʟ��� ٟ���6�!�Z�E�W�t��#1( ��9��K���ĥ ������Ư!3�8�x��!4Mgs���,�IB+8�J��a���{�d� d�����ȿ���ڼ%%P8�P�=:G����S�6�h�z���R��Ϯ����������  %�� ��h�Vߌ� z߰�&�g�/9�$�������7����A�8S�e�w�  ��������������2 �F�$�&Gb���������!C���@���8������F� DzN��� F�P D�!������)#B�'�9K]o#?��W�@@v
4$8��8��8�.
 v���! 3EWi{�����:� ��ۨ��1��$MSK�CFMAP  ���� ����(.�ONR�EL  ��!9��EXCFE�NBE'
#7%^!F�NCe/W$JOGO/VLIME'dO S"]d�KEYE'�%]�RUN�,�%��SFSPDT�Y0g&P%9#SIG�NE/W$T1MOT��/T!�_CE_�GRP 1p��#\x��?p��?�? �?�?�?O�?OBO �?fOO[O�OSO�O�O �O�O�O_,_�OP__ I_�_=_�_�_�_�_�_�oo�_:o�TC�OM_CFG 1�q	-�vo�o�o
�Va_ARC_b"��p)UAP_CP�L�ot$NOCHE�CK ?	+ �x�%7I [m���������!�.+NO_?WAIT_L 7%6S2NT^ar	+��s�_ERR_129s	)9�� ,ȍޏ��x���&��d�T_MO��t��,� ��*oq�9�P�ARAM��u	+��a�ß'g{��� =?�345678901��,�� K�]�9�i�������ɯۯ��&g������C��cUM_RSP�ACE/�|����$ODRDSP�c�#6p(OFFSET�_CART�o��D�ISƿ��PEN_FILE尨!�ai���`OPTION_�IO�/��PWOR�K ve7s# ��V�ؤ��p�4�p�	 ���p���<���RG_DS�BL  ��P#���ϸ�RIENTkTOD ?�C�� �!l�UT_SIM_D$�"����V��LCT w�}�h�iĜa[�1�_P�EXE�j�RAT�vШ&p%� ��2^3j�)TEX)TH�>)�X d3��� ����%�7�I�[�m� ������������ �!�3�E���2��u� ��������������c�<d�ASew ���������Ǎ�^0OUa0o(��(����}u2, ����O H @D�  &[?�aG?��c�c�D][�Z�;��	ls���xJ���������<; ��� ��2��H(��H3k7�HSM5G�22�G���Gp
͜�'f�/-,2�KCR�>�D!�M#�{Z/��3�����4y H "�c/�u/�/0B_�����jc��t�!�/ �/�"t3�2����/6  U��P%�Q%��%��|T��S62�q?'e	�'� � �2�I� �  {��+==��ͳ?��;	�h	�0�I  �n @�2 �.��Ov;��ٟ?r&gN�]O  ''��uD@!� C�C�@�F#H!�/�O�O sb
S���@�@���@�e`0B�QA8�0Yv: �13Uwz$oV_�/z_e_�_��_	��( �� -�2�1�1ta�Ua�c���:A-����.  �?�fAf���[o"o�_Uʈ`oXÜQ8���o�j>N�1  Po�V(�� �eF0�f�Y���L�/?����xb�P�<
6b<߈�;܍�<�ê�<� <�&�,/aA�;r�@Ov�0P?fff?�0?y&ip�T@�.{r�J<?�`�u #	�Bdqt�Yc�a �Mw�Bo��7�"� [�F��j�������ُ ����3�����,���(�E�� E���3G+� F� �a��ҟ�����,���P�;���B�pA Z�>��B��6�<OίD� ��P��t�=���a�s�x����6j�h��7o��>�S��O�`����Fϑ�A�a�_��C3Ϙ�/�%?��?���������
#	Ę��P �N||#CH���Ŀ����ރ�@I�_�'��3A�A�AR�1AO�^?�$��?��� �±�
=ç>�����3�W
=�#�� U��e���B���@��{�����<���(��B�u��=�B0�������	�b�H�F��G���G���H�U`E����C�+��I#��I��HD��F��E���RC�j=[�
�I��@H��!H�( E<YD0߻���� ����� �9�$�]�H� Z���~����������� ��#5 YD}h ������� 
C.gR��� ����	/�-// */c/N/�/r/�/�/�/ �/�/?�/)??M?8? q?\?�?�?�?�?�?�? �?O�?7O"O[OmOXO �O|O�O�O�O�O�O�O��O3_Q(�������b��gUU���W_i_2�3�8���_�_2�4Mgs8�_�_�RIB+�_�_��a���{� miGo5okoYo�o}lJ��P'rP�nܡݯ��o=_�o�_�[R?Q�u���  �p���o�� /��S��z
uүܠ�������ڱ������p�����  /��M�w�e��������l2� F�$��Gb	��t��a�`�p�S�C�y�@p�5�G�Y�~۠F� Dz���� F�P DC��]����پ���ʯܯ� ��~�?̯��@@�?�RK�K���K���
 �|������� Ŀֿ�����0�B�pT�fϽ�V� ���{���1��$PA�RAM_MENU� ?3���  DEFPULSEr��	WAITTM�OUT��RCV��� SHEL�L_WRK.$CUR_STYL��;	�OPT�ߧPTB4�.�C�R?_DECSN���e ��ߑߣ��������� ��!�3�\�W�i�{�����USE_PR_OG %��%��\���CCR���e�����_HOST !��!��:���AT�`�V��/�X�|����_TIME���^��  ��GD�EBUG\�˴�G�INP_FLMS�K����Tfp����P+GA  ����)�CH����TYPE
�������� ��� -?h cu������ �//@/;/M/_/�/ �/�/�/�/�/�/�/?�?%?7?`?��WOR�D ?	=	�RSfu	PNS2UԜ2JOK�DR�TEy�]TRA�CECTL 1xv3��� �`_� &�`�`|�>�6DT Qy3��%@�0D � ��c�aa:@V�@BR�2O DOVOhOzO�O�O�O�O@�O�O�O
__.Z<TDT,Sb_t_�_�Z]_�SM �R._@_RXN\L�
o�["c P_�_�VJ�PbF��WJ`UNd	Nd
NdNdNd5of@oRodovo �o�o�o�o�o�o (:L^p�����r�t^��r�t��t�t�|��r*�t�t�t�|j�
�r�t�tҀ�r���z"�t#�t��r%��t&�|(�t)�t*��t+�t,�|.�t/
�t0�t1�YJ�\�n� ��������ȟڟ��� �"�4�F�X�.Iv��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p��j�� ��� $6H Zl~����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o� �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ����������*��$PGTRA�CELEN  �)�  ���(��>�_UP z���mљu�Y�n�>�_�CFG {m�)W�(�n���P���� ��DEFSP/D |��'�P���>�IN��TR�L }��(�8���IPE_CON�FI��~m��mњ��Ԛ�>�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�8��1��� ´�����B�9����O��9�s�(�>�T?��
5�������� �=��=#�
 ����P;t_�������� G Dz (�
 H�X~i��� ���/�/D///�h/S/�/��
V7�.10beta1���  A��E�"ӻ�A �(�� ?!G��!>����"����!{���!BQ��!�A\� �!���!2p
����Ț/8?J?\?�n?};� ���/� �/�?}/�?�?OO:O %O7OpO[O�OO�O�O �O�O�O_�O6_!_Z_ E_~_i_�_�_�_�_�_ �_'o2o�_VoAoSo �owo�o�o�o�o�o�o .R=v1�/�#F@ �y�}� �{m��y=��1�'� O�a��?�?�?������ ߏʏ��'��K�6� H���l�����ɟ��� ؟�#��G�2�k�V� ��z��������o� �ίC�.�g�R�d��� �������п	���-� ?�*�cώ���Ϯ� �����B�;�f� x�������DϹ��߶� �������7�"�[�F� X��|��������� ��!�3��W�B�{�f� �������� ����� /S>wbt� �����= OzόϾψ����� �� /.�'/R�d�v� �߁/0�/�/�/�/�/ �/�/#??G?2?k?V? h?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O���O�O�O__ ?_*_c_N_�_r_�_�_ �_�_�_o�_)oTf x�to���/�o />/P/b/t/m o�|����� ��3��W�B�{�f� x�����Տ������ �A�S�>�w�b����O ��џ������+�� O�:�s�^�������ͯ ���ܯ�@oRodo�o `��o�o�o��ƿ�o� ��*<N�Y��}� hϡό��ϰ������� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�c�N�ﲟ��� l��������;�&� _�J���n��������� ��,�>�P�:L�� ���������� (�:�3��0iT� x�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?a?s?��?�?X?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O *\&_8_r����_�_��$PLI�D_KNOW_M�  ��� Q�TSV ���P��?o"o4o�OXo�CoUo�o R�SM_?GRP 1��Z'U0{`�@�`uf
�e�`
�5� �gpk 'Pe] o�������X���SMR�c��m1T�EyQ}? yR�� ��������폯���ӏ �G�!��-������� ����韫���ϟ�C� ��)������������寧���QST�a1W 1��)���P;0� A 4��E 2�D�V�h�������߿ ¿Կ���9��.�o� R�d�vψ��ϬϾ�����2�0� Q�	<3��3�/�A�S߂�4l�~ߐߢ��5 ���������6
��.�@��7Y�k�}���8��������M_AD  )���PARNUM  !�}o+��WSCHE� S�
��pf���S��UPDf��x��_CM�P_�`H�� �'��UER_CHK-���ZE*<�RSr��_�Q_MO�G���_�X�_R/ES_G��!��� D�>1bU� y�����/�	/����+/� k�H/g/l/��Ї/�/ �/�	��/�/�/�X� ?$?)?���D?c?h?�����?�?�?�V �1��U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_�INRr�J�b�Ud�2FMASS?O Z�SGMN>OqCMON�_QUEUE a��U�V P~P X�N$ UhN�FV�@�END�A��IEX1E�O�E��BE�@�O>�COPTIO�G���@PROGRAM7 %�J%�@�?����BTASK_I�G�6^OCFG ኤOz��_�PDATuA�c��[@Ц2=�DoVohozo�j2o �o�o�o�o�o)x;M jINFO[��m��D��� �����1�C�U� g�y���������ӏ����	�dwpt�l �)�QE DIT ��_i��^WERF�LX	C�RGADoJ �tZA���¿�?נʕFA��IOORITY�GW���MPDSPNQ�����U�GD��OTO�E@1�X� (/!AF:@E� c�~Ч!tcpn�>��!ud����!icm���?<��XY_�Q�X�=��Q)� *�1�5��P��]�@�L� ��p��������ʿ� �+�=�$�a�Hυϗ�=*��PORT)QH���P�E��_C?ARTREPPX�>�SKSTA�H�
�SSAV�@�tZ	�2500H86A3���_x�
�'��X�@�swPtS��x�ߧ���URGE�@�B��x	WF��DO�F"[W\��������WRUP_DEL�AY �X���RO_HOTqX	B%��c���R_NORM�ALq^R��v�SE�MI�����9�QS�KIP'��tUr�x 	7�1�1�� X�j�|�?�tU������ ��������$J \n4����� ���4FX |j������ �/0/B//R/x/f/�/�/�/tU�$RCgVTM$��D�� �DCR'������!A���BX�KC31d?�<��:�.��:����u� ��������%��:�o?�� �<
6b<߈�;܍�>u.��?!<�& �?h?�?�?�@>��?O  O2ODOVOhOzO�O�O �O�O�O�?�O�O__ @_+_=_v_Y_�_�_�? �_�_�_oo*o<oNo `oro�o�o�o�_�o�o �o�o�o8J-n ��_������ �"�4�F�X�j�U�� ����ď���ӏ�� �B�T��x������� ��ҟ�����,�>� )�b�M����������� �ïկ�Y�:�L�^� p���������ʿܿ�  ����6�!�Z�E�~� ��{ϴϗ�����-��  �2�D�V�h�zߌߞ� ����������
���.� �R�=�v��k��� �������*�<�N� `�r������������ ����&J\? �������� "4FXj|���!GN_ATC �1�	; �AT&FV0E0��ATDP/6/9/2/9��ATA�,�AT%G1%B�960�++U+�,�H/,�!�IO_TYPE � �%�#t�R�EFPOS1 1}�V+ x�u/�n�/j�/
=�/ �/�/Q?<?u??�?4?�?X?�?�?�+2 1�V+�/�?�?\O�?x�O�?�!3 1�O�*O<OvO�O�O_�OS4 1��O�O�O_��_t_�_+_S5 1�B_T_f_�_o	oBo>�_S6 1��_�_��_5o�o�o�oUoS7 1�lo~o�o�oH�3l�oS8 1� %_����SMASK 1��V/  
?�M��XNOS/�r�����~�!MOTE  n���$��_CFG ᢫��q���"PL_�RANG�����POWER ������SM_DRYPRG %o��%�P��TART� ��^�UME_PRO-�?����$�_EXEC_EN�B  ���GS�PD��Րݘ��T3DB��
�RM�
��MT_'�T�����OBOT_NA_ME o�����OB_ORD_�NUM ?��b!H863�  �կ����PC_TIMoEOUT�� x�oS232Ă1��� LTEA�CH PENDA1N��w��-���Mainte�nance Co#ns���s�"���?KCL/Cm��
�
���t�ҿ ?No Use-��8Ϝ�0�NPO�򁮋���.�C7H_L������q�	��s�MAVA#IL�����糅���SPACE1 2��, j�߂�D��s�߂� �{S�?8�?�k�v� k�Z߬��ߤ��ߚ�  �2�D���hߊ�|�� `����������  �2�D��h��|����`���������y���2����0�B���f� ����{���3);M_ ������/� /44FXj| */���/�/�/?(??=?5Q/c/u/�/ �/G?�/�/�?O�?$OEO,OZO6n?�?�? �?�?dO�?�?_,_�O A_b_I_w_7�O�O �O�O�O�_�O_(oIo@o^oofo�o8�_ �_�_�_�_�oo6oE�f){���Gw �o� �:��
M� ��� *�<�N�`�r������� w���o�収���d.��%�S�e�w��� ��������Ǐَ��� Θ8�+�=�k�}����� ��ůׯ͟����%� '�X�K�]��������� ӿ������#�E��W� `� @ �������x�����\�e����������� R�d߂�8�j߬߾߈� �ߤ����������0� r���X�������@������8����
�����_MODE � �{��S �"�{|�2�0��ψ��3�	S|)CWORK_AD���k�|+R  ��{�`� �� _?INTVAL���d����R_OPTI[ON� ��H �VAT_GRP �2��up#(N�k| ��_����� /0/B/��h�u/T�  }/�/�/�/�/�/�/? !?�/E?W?i?{?�?�? 5?�?�?�?�?�?O/O AOOeOwO�O�O�O�O UO�O�O__�O=_O_ a_s_5_�_�_�_�_�_ �_�_o'o9o�_Iooo �o�oUo�o�o�o�o�o �o5GYk-� ��u����� 1�C��g�y���M��� ��ӏ叧�	��-�?� Q�c������������ ���ǟ�;�M�_�����$SCAN_GTIM��_%}��R �(�#(�(�<04+d d 
!AD�ʣ��u�/X�����U���25���@�d5�P�g��]	�������p��dd�x�  P����� �� � 8� ҿ�!���D��$�M�_�qσ� �ϧϹ��������ƿv��F�X�x�/� ;�ob���pm��t�_DiQ̡  � l�|�̡ĥ �������!�3�E�W� i�{���������� ����/�A�S�e�] �Ӈ������������� );M_q� ������ r���j�Tfx�� �����//,/ >/P/b/t/�/�/�/�/8�/�%�/  0��6 ��!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O* �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo�O �OJ�o�o�o�o�o�o �o 2DVhz �������
�7?  ;�>�P�b� t���������Ǐُ� ���!�3�E�W�i�{�p������ß �ş 3�ܟ��&�8�J�\�@n�������������ɯ����,� ��+�	123�45678�� +	� =5���f� x����������� ��
��.�@�R�d�v� �Ϛ�៾�������� �*�<�N�`�r߄߳� �ߺ���������&� 8�J�\�n�ߒ��� ���������"�4�F� u�j�|����������� ����0_�Tf x������� I>Pbt� ������!/ (/:/L/^/p/�/�/�/�/�/�/�2�/?��#/9?K?]?�iC�z  Bp˚  � ��h2��*��$SCR_GRP� 1�(�U8(�\xd��@ � ��'�	 �3�1�2 �4(1*�&�I3�F1O�OXO}m��D!�@�0ʛ)���HUK��LM-10i�A 890?�90�;��F;�M61CA D�:�CP��1
\&V�1	�6F��CW�9)A7Y	(R�_�_Ф_�_�_�\�� �0i^�oOUO>oPo #G�/���o'o�o�o\�o�oB�0��rtAA�0*  !@�Bu&Xw?��ju��bH0{UzAF@ F�`�r��o �����+��O� :�s��mBqrr����������B�͏b���� 7�"�[�F�X���|��� ��ٟğ���N���AO�0�B�CU
L���E��jqBq>g�#H@��@pϯ B����G�I
E�0EL_�DEFAULT � �T���E��MIPO�WERFL  �
E*��7�WFDO�� *��1ERV�ENT 1����`(�� L!DUM_EIP���>��j!AF_�INE�¿C�!�FT������!�o:� ��a�!�RPC_MAI�Nb�DȺPϭ�t�V�IS}�Cɻ����!7TP��PU�ϫ��d��E�!
PMON_PROXYF߂��e4ߑ��_ߧ�f�����!RDM_'SRV�߫�g��)�G!R�Iﰴh�u�!
v�M�ߨ�i�d���!RLSY3NC��>�8����!ROS��4��4��Y�(�}���J�\� ������������7 ��["4F�j| ����!�E�io�ICE_KL� ?%� (%�SVCPRG1@n>���3��3�D��4//�5./D3/�6V/[/�7~/ �/��D�/�9�/�+�@��/��#?� �K?��s?� /�? �H/�?�p/�?��/ O��/;O��/cO� ?�O�9?�O�a?�O ��?_��?+_��? S_�O{_�)O�_� QO�_�yO�_��Os ����>o�o}1�o �o�o�o�o�o�o ;M8q\��� ������7�"� [�F��j�������ُ ď���!��E�0�W� {�f�����ß���ҟ ���A�,�e�P��� t��������ί�y_DEV ���MC:�w�_!�OUT���2��REC �1�`e�j� �	 �����˿඿�ڿ��
 � `e���6�N�<�r�`� �τϦ��Ϯ������� &��J�8�n߀�bߤ� ���߶�������"�� 2�X�F�|�j����� ���������.�T� B�x�Z�l��������� ����,P>` bt����� �(L:\�d ����� /�$/ 6//Z/H/~/l/�/�/ �/�/.��/?�/2? ? V?D?f?�?n?�?�?�? �?�?
O�?.O@O"OdO RO�OvO�O�O�O�O�O �O__<_*_`_N_�_ �_x_�_�_�_�_�_o o8oo,ono\o�o�o �o�o�o�o�o�o  "4jX���� ������B�$� f�T�v���������� ��؏��>�,�b�P�xr���p�V 1�}�� P
�	!��^��� ���TY�PE\��HELL_CFG �.�<F��  	�����RSR������ ӯ�������?�*� <�u�`��������������  �%�3�E��Q�\��ҰM�o�p��d��2Ұd]�K�:��HK 1�H� u�������A�<� N�`߉߄ߖߨ����� ������&�8��=�?OMM �H����9�FTOV_EN�B&�1�OW_R�EG_UI���I_MWAIT��a�.��OUT������wTIM������VAL����_UN�IT��K�1�MON�_ALIAS ?�ew� ( he �#����������Ҵ�� );M��q�� ��d��% �I[m�<� �����!/3/E/ W//{/�/�/�/�/n/ �/�/??/?�/S?e? w?�?�?F?�?�?�?�? �?O+O=OOOaOO�O �O�O�O�OxO�O__ '_9_�O]_o_�_�_>_ �_�_�_�_�_�_#o5o GoYokoo�o�o�o�o �o�o�o1C�o gy��H��� �	��-�?�Q�c�u�  �������ϏᏌ�� �)�;��L�q����� ��R�˟ݟ����� 7�I�[�m��*����� ǯٯ믖��!�3�E� �i�{�������\�տ �����ȿA�S�e� wω�4ϭϿ����ώ� ���+�=�O���s߅� �ߩ߻�f������� '���K�]�o���>� ����������#�5� G�Y��}����������n��$SMON_�DEFPRO ������� *SY�STEM*  d�=��RECAL�L ?}�� (� �}4copy� frs:ord�erfil.da�t virt:\�tmpback\�=>inspir�on:11828���s��  }+�.mdb:*.*�CUZ���/x.:\�8R�Po���0.a6 H__�//�- ?�b/t/�/�/�F/ �a/�/??)�M �/p?�?�?�8?J?� �? OO%/7/�/�/lO ~O�O�/�/PO�/�O�O _!?3?�?W?h_z_�_ �?�?B_�?�_�_
oO /OAOSOdovo�oo�O Ho�O�o�o+_�_ O_�or���_:L _���'o9o�o�o n������o��o[�� ���#5�Yj�|� ����D������ �1���U�f�x����� ��J�ӏ������-� ��Q�b�t�������<� ϟa����)�;�į ߿pςϔϧ���˯]� �� ��%���ʿ[�l� ~ߐߣ���F�ٿ���� �!�3ϼ�W�h�z�� �ϱ�L�������
�� /���S�d�v������ >�������+�=� ����r����D�� _�'�����]� n����6H�����/#
xyzrate 61 �@��n/�/�/%.'>R3304 H/Z/�/�/?"3.@�- a?s?�?�?* *�I?��$Y?�?�?O!�$�SNPX_ASG 1����9A�� P �0 '%R[1]@1.1O 	?�#%dO�OsO �O�O�O�O�O�O __ D_'_9_z_]_�_�_�_ �_�_�_
o�_o@o#o doGoYo�o}o�o�o�o �o�o�o*4`C �gy����� ��	�J�-�T���c� ������ڏ����� 4��)�j�M�t����� ğ������ݟ�0�� T�7�I���m������� �ǯٯ���$�P�3� t�W�i��������ÿ ����:��D�p�S� ��wω��ϭ��� ��� $���Z�=�dߐ�s� �ߗߩ������� �� D�'�9�z�]���� �����
����@�#� d�G�Y���}������� ������*4`C �gy����� �	J-T�c ������/� 4//)/j/M/t/�/�/ �/�/�/�/�/?0?4�,DPARAM �9ECA ��	��:P�4�0�$HOFT_KB_?CFG  p3?E��4PIN_SIM  9K�6�?�?��?�0,@RVQST_P_DSB�>�2�1On8J0SR ���;� & MU�LTIROBOT�TASK=Op3��6TOP_ON_?ERR  �F�8~�APTN �5��@A�BRING_PRM�O� J0VDT_G�RP 1�Y9�@  	�7n8_(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2Dkhz �������
� 1�.�@�R�d�v����� ����Џ�����*� <�N�`�r��������� ̟ޟ���&�8�J� \�����������ȯگ ����"�I�F�X�j� |�������Ŀֿ�� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�tߛߘߪ� ����������(�:� a�^�p������� ���� �'�$�6�H�Z� l�~���������������3VPRG_CO7UNT�6��A�5NENB�OM=��4J_UPD 1}��;8  
 p2������  )$6Hql~� ����/�/ / I/D/V/h/�/�/�/�/ �/�/�/�/!??.?@? i?d?v?�?�?�?�?�? �?�?OOAO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_��_�_YSDEBSUG" � �Pdk	��PSP_PASS�"B?�[LOG� ��mr�P�X�_  �g~�Q
MC:\d<�_b_MPCm�H�o�o�Qa�o �~vfSAV �m�:dUb�U\gS�V�\TEM_TI�ME 1�� �() �%��o	T1SVGUNS} �#'k�spAS�K_OPTION�" �gospBC?CFG ��|� �b�{�}` ����a&��#�\�G� ��k�����ȏ����� �"��F�1�j�U��� y���ğ���ӟ��� 0��T�f��UR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz�ʠrBrv�x����z� �%�� I�4�m�X���|����� ���֏���3��W� B�g���x�����՟�� ������S�>�w� b�����'2A ��ʯܯ ������E�0�i�T� ��x���ÿտ翢�� ��/��?�e�1�/�� �/�ϜϮ�������� ,��P�>�`߆�tߪ� ���߼�������� L�:�p�^����� ������� �6�H�>/ `�r������������ ���� 0Vhz 8������
 .�R@vd� ������// </*/L/r/`/�/�/�/ �/�/�/�/�/?8?&? \?J?�?n?�?�?�?�? ���?OO�?FO4OVO XOjO�O�O�O�O�O�O __�OB_0_f_T_v_ �_�_�_z_�_�_�_o o>o,oboPoroto�o �o�o�o�o�o( 8^L�p��� ����$��H�6� l�~�(O����f�d�� ؏���2� �B�D�V� ������n����ԟ
� ��.�@�R�d����v� �������Я���*� �N�<�^�`�r����� ̿���޿��$�J� 8�n�\ϒπ϶Ϥ��� ����ߊ�(�:�L��� |�jߌ߲ߠ������� ���0�B�T��x�f� ������������� ,��P�>�t�b����� ����������: (JL^���� �� �6$Z H~l��^��� dߚ //D/2/h/V/ x/�/�/�/�/�/�/�/ ?
?@?.?d?v?�?�? T?�?�?�?�?�?OO <O*O`ONO�OrO�O�O �O�O�O_�O&__6_ 8_J_�_n_�_�_�_�_ �_�_�_"ooFo�� po�o,oZo�o�o�o�o �o0Tfx� H������� ,�>��b�P���t��� ������Ώ��(�� L�:�p�^�������ʟ ���ܟ� �"�$�6� l�Z���~�����د� �o��&�ЯV�D�z� h�������Կ¿��
� �.��R�@�v�dϚ�΄�  ���� ��������$TB�JOP_GRP �2ǌ��?  ?������������xJBЌ���9� �<� �X���� �@���	 �C��� t�b  C�x���>��͘�̐դ�>̚йѳ33=�CLj��fff?��?�ffBG��ь�����t޽ц�>�(��\)�ߖ�E噙��;��hCYj���  @h��B� � A����f��C�  Dhъ�1����O�4�N�����
:���Bl^��j�i�l�l����?Aə�A�"��sD��֊=qH����нp�h�Q�;�A�j��ٙ�@L��D	�2�������$�6�>BÏ\��T���Q�ts}x�@33@���C���y�1����>��Dh�����������<{�h�@i� �� t��	���K &�j�n|�� �p�/�/:/k/��ԇ���!��	�V3.00J�m761cI�*� I�����/�' Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,I�!C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^��;Q�T,8�4E` *�ϴ?�2����3\�X/O��ES�TPARS  ظ�	���HR@AB_LE 1����0��
H�7 8��9
G�
H
H����
G	�
H

H
HYE���
H
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_ P_b_t_�^:BS _� �JGoYoko}o�o�o �o�o�o�o�o1 CUgy����` #oRL�y�_�_�_�_�O��O�O�O�OX:B�rN�UM  ��*�P��� V@P�:B_CFG �譋Z�h�@��IMEBF_TT%AU��2@�VERS�q���R 1���
' (�/����b� ����J�\���j�|� ��ǟ��ȟ֟���� �0�B�T���x��������2�_���@�
���MI_CHAN��� � ��DBGLV����������ETHERAD �?��O���ಯ��h�����ROUmT�!��!�������SNMASK�D��U�255.����#�����OOL�OFS_DI%@��u.�ORQCTRL �����}ϛ3 rϧϹ��������� %�7�I�[�:���h�z����APE_DET�AI"�G�PON_�SVOFF=���P_MON �֍��2��STRTC_HK �^������VTCOMPA�T��O�����FPR�OG %^�%�MULTIROB�OTTݱ���9�P�LAY&H��_IN�ST_Mް �������US�q��L�CK���QUIC�KME�=���SC�REZ�G�tps� ���u�z�����_��@@n�.�S�R_GRP 1о^� �O� ���
��+O=sa�쀚�
m�� ����L/C 1gU�y��� ��	/�-//Q/?/�a/�/	1234�567�0�/�/@X�t�1���
 �}�ipnl/� g?en.htm�?� ?2?D?V?`P�anel setupZ<}P�?�?�?�?�?�? �??,O >OPObOtO�O�?�O!O �O�O�O__(_�O�O ^_p_�_�_�_�_/_]_ S_ oo$o6oHoZo�_ ~o�_�o�o�o�o�o�o so�o2DVhz� 1'���
�� .��R��v��������ЏG���UALR�M��G ?9� �1�#�5�f�Y��� }�������џן����,��P��SEV � ����E?CFG ������A��   BȽ�
 Q���^� ���	��-�?�Q�c�@u�������������C �����I��?���(%D�6� � $�]�Hρ�lϥϐ��� ��������#��G����� �߿U�I_�Y�HIST 1վ�  (��� ��3/SOF�TPART/GE�NLINK?cu�rrent=editpage,��,1���!�3���� ����menu��962�߆���0��K�]�o�36u�
� �.�@���W�i�{��� ������R����� /A��ew��� �N��+= O�s��������f��f//'/ 9/K/]/`�/�/�/�/ �/�/j/�/?#?5?G? Y?�/�/�?�?�?�?�? �?x?OO1OCOUOgO �?�O�O�O�O�O�OtO �O_-_?_Q_c_u__ �_�_�_�_�_�_�� )o;oMo_oqo�o�_�o �o�o�o�o�o%7 I[m� �� �����3�E�W� i�{������ÏՏ� ������A�S�e�w� ����*���џ���� �ooO�a�s����� ����ͯ߯���'� ��K�]�o��������� F�ۿ����#�5�Ŀ Y�k�}Ϗϡϳ�B��� ������1�C���g� yߋߝ߯���P����� 	��-�?�*�<�u�� ������������ )�;�M���������� ������l�%7 I[������ �hz!3EW i������� v////A/S/e/P����$UI_PA�NEDATA 1������!�  	�}�w/�/�/�/�/?? )?>?��/i?{?�? �?�?�?*?�?�?OO OAO(OeOLO�O�O�O��O�O�O�O�O_&Y� b�>RQ?V_h_ z_�_�_�__�_G?�_ 
oo.o@oRodo�_�o oo�o�o�o�o�o�o *<#`G��}�-\�v�#�_�� !�3�E�W��{��_�� ��ÏՏ���`��/� �S�:�w���p����� џ������+��O� a���������ͯ߯ �D����9�K�]�o� �������ɿ���Կ �#�
�G�.�k�}�d� �ψ����Ͼ���n��� 1�C�U�g�yߋ��ϯ� ��4�����	��-�?� ��c�J������ ���������;�M�4� q�X����������� %7��[�� �����@� �3WiP�t �����/�// A/����w/�/�/�/�/ �/$/�/h?+?=?O? a?s?�?�/�?�?�?�? �?O�?'OOKO]ODO �OhO�O�O�O�ON/`/ _#_5_G_Y_k_�O�_ �_?�_�_�_�_oo �_Co*ogoyo`o�o�o �o�o�o�o�o-`Q8u�O�O}��@������)� >��U-�j�|������� ď+��Ϗ���B� )�f�M���������������ݟ�&�S�K��$UI_PANELINK 1�U�  ��  ��}1�234567890s���������ͯդ �Rq����!�3�E�W� �{�������ÿտm��m�&����Qo�  �0�B�T�f�x�� v�&ϲ���������� ��0�B�T�f�xߊ�"� �����������߲� >�P�b�t���0�� ����������$�L� ^�p�����,�>�����`�� $�0,&� [gI�m��� ����>P3 t�i��Ϻ�  -n��'/9/K/]/o/ �/t�/�/�/�/�/�/ ?�/)?;?M?_?q?�? �UQ�=�2"��?�? �?OO%O7O��OOaO sO�O�O�O�OJO�O�O __'_9_�O]_o_�_ �_�_�_F_�_�_�_o #o5oGo�_ko}o�o�o �o�oTo�o�o1 C�ogy���� �B�	��-��Q� c�F�����|������ �֏�)��M���= �?��?/ȟڟ��� �"�?F�X�j�|��� ��/�į֯����� 0��?�?�?x������� ��ҿY����,�>� P�b��ϘϪϼ��� ��o���(�:�L�^� �ςߔߦ߸������� }��$�6�H�Z�l��� ����������y��  �2�D�V�h�z���� -���������
��. RdG��}� ���c���<�� `r������� �//&/8/J/�n/ �/�/�/�/�/7�I�[� 	�"?4?F?X?j?|?� �?�?�?�?�?�?�?O 0OBOTOfOxO�OO�O �O�O�O�O_�O,_>_ P_b_t_�__�_�_�_ �_�_oo�_:oLo^o po�o�o#o�o�o�o�o  ��6H�l~ a������� �2��V�h�K����� ��1�U
��.� @�R�d�W/�������� П������*�<�N� `�r��/�/?��̯ޯ ���&���J�\�n� ������3�ȿڿ��� �"ϱ�F�X�j�|ώ� �ϲ�A��������� 0߿�T�f�xߊߜ߮� =���������,�>� ��b�t�����+ ������:�L�/� p���e�����������  ��6���ۏ���$UI_QU�ICKMEN  }���}���RESTOR�E 1٩�  �
�8m3\n ���G���� /�4/F/X/j/|/' �/�/�//�/�/?? 0?�/T?f?x?�?�?�? Q?�?�?�?OO�/'O 9OKO�?�O�O�O�O�O qO�O__(_:_�O^_ p_�_�_�_QO[_�_�_ I_�_$o6oHoZoloo �o�o�o�o�o{o�o  2D�_Qcu�o �������.� @�R�d�v��������xЏ⏜SCRE� �?�u1�sc� u2�3��4�5�6�7��8��USER�����T���ksT'���4��5��6���7��8��� NDO_CFG ڱ�  �  � PD�ATE h���None�S�EUFRAME � ϖ��RTOL_ABRT�����ENB(��G�RP 1��	�?Cz  A�~�|��%|�������į֦��X�� UH�X�7�?MSK  K�S��7�N�%uT�%������VISCA�ND_MAXI��I�3���FAILO_IMGI�z �% �#S���IMREG�NUMI�
���S�IZI�� �ϔ�,�ONTMOU4'�K�Ε�&�����a��a���s�FR:\��� � M�C:\(�\LOGnh�B@Ԕ !{��Ϡ�����z �MCV����7UD1 �EX	��z ��PO64_t�Q��n6��PO!�LI�Oڞ�re�V�N�f@`��I�� =	_�SZ�Vmޘ��`�WA�Imߠ�STAT �k�% @��4�F��T�$#�x �2D�WP  ��P� G��=��������_JMP�ERR 1ޱ
�  �p2345678901��� 	�:�-�?�]�c����� ������������$�MLOW�ޘ�����g_TI/�˘'���MPHASE  �k�ԓ� ��SH�IFT%�1 Ǚ��<z��_� ���F/| Se������ �0///?/x/O/a/��/�/�/�/�/�����k�	VSFT1�\�	V��M+3 S�5�Ք p���ſA�  B8[0�[0�Πpg3a1Y2�_3Y�7ME��K�͗q	6e���&%���M���b��	���$��TDINEND3�4��4OH�+�G�1�OS2OIV I�{��]LRELEv�I��4.�@��1_AC�TIV�IT��B��A �m��/_��B�RDBГOZ�YBO�X �ǝf_\���b�2�TI�190.0.�P8�3p\�V254tp^�Ԓ	 �S��_�[b��r�obot84q_   p�9o\�pc�PZoMh�]�Hm�_Jk@1�o�ZA+BCd��k�,���P \�Xo}�o0); M�q����� ���>��aZ�b��_V