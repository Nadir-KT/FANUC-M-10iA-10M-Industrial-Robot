��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  V � �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1��GPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|~GRG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"GSB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5H UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8�GW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3��B�2���AXD��#
 d $�CARD_EXI�ST4$FSS�B_TYP!AH�KBD_SNB�1A�GN Gn $�SLOT_NUM��APREV4D�EBU� g1(��;1_EDIT1� � 1G=�� S�0%$EP<�$OP��U0LETE_O�K�BUS�P_CR�A$;4AV� 0/LACIw1�Rp�@k �1$@MEN�@$D�V�Q`Pv�VA{G BL� OU&R ,A�0��!� B� LM_O��
eR�"CAM_�;1 xr$ATTR4�@� �ANNN@5IMG?_HEIGH�AXc�WIDTH4VT�� �UU0F_ASwPEC�A$M�0gEXP�.@AX�f��CF�D X O$GR� � S�!z.@B�PNFLI�`<�d� UIRE 3T�!GITCH+C�`N�� S�d_LZ`ACL�"�`EDp�dL� J�4S�0� <za�!�p;G0 � 
$WARNM�0�f�!�@� -s�pNS=T� CORN�"a1�FLTR{uTRA�T� T}p  $ACCa1�p��|{�rORI�P�C�k�RT0_S~B\qHuG,I1 [ �T�`�"3I�pTYPD�@*2 3`#@�� �!�B*HDDcJ�* Cd�2_�3_�4�_�5_�6_�7_�8r_�94�@�CO�$ <� �o�o�hK3� 1#`O_Mc@AC/ t � E#63NGPvABA� �c�1�Q8��`,��@nr1�� d�P�0e�]p,� cvnpUP&P�b26���p�"J�p_)R�rPBC��J�rĘߜJV�@U� B��s}��g1�"YtP_*0O�FS&R @� RcO_K8T��aIT�3�T�NOM_�0�1�p�34 >��D Ԑ� Ќ@��hPV��mE!X�p� �0g0ۤ�p��r
$TF�2C$7MD3i�TO�3�0yU� F� ��)Hw2tC1(�Ez�g0#E{"F�"F�40�CP@�a2 �@�$�PPU�3Nc)ύRևAX�!�DU��AI�3B�UF�F=�@1 �|pp���pPITV� PP�M�M��y��F�SIMQ�SI�"ܢVAڤT��=�w T�`(zM��P�B�qFACTb�@EW�P1��BTv?�MC�5 �$*1JB`p�*1DEC��F��ů���� �H0CHNS_EMP1�G$G��8��@_4��3�p|@P��3�TC c�(r/�0-sx��ܐ�� MBi��!����JR|� i�SEGFR���Iv �aR�TpN�C��PVF4>�bx &��f{u Jc!�Ja��� !28�ץ8�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb��Ӏq�۽�н����Lp�3�B���CRC�e�3CCp����c� �mcҞb�1J�cѿ�.�T���D$ICb�Cq��5r�ե��@v�'���E�V���zF��_��FR,pN��ܫ�?�84�0A�! �r�� �h�Ϩ��p�2�͕a��� �د�R�Dx Ϗ��o"2�7�!ARV�O`C�$LG�pV�B�1�P��@�t�aA�0'�|�+01Ro�� MEp`"1� CRA 3 A�ZV�g6p�O �FCCb�`�`F�`K������ADI��a� A�bA'�.p��p�`��c�`S4PƑ�a�AMIP��-`Y�3P�M��]pUR��QUA1  ]$@TITO1/S�@S�!����"0�DBOPXWO��B0!5�O$SK���28@�DBq�!"�"�PR�� 
� =���΁!# S q1$�2�$z���L�)$��/���� %�/�$Cr�!&?�$ENE�q�.'*?�Ú RE|�p2(H ���O�0#$L|3$�$�#�B[�;���FO�_D��ROS�r�#������3RIoGGER�6PApS|����ETURN�2n�cMR_8�TUw���0EWM���M�GN�P���BLA�H�<E���P��&$P� �'P@�Q3�CkD{��DQ���4��11��FGO_AWAY�BMO�ѱQ#!�� CS_�)  �PIS� I g�b {s�C��A��[  �B$�S��AbP�@�E9W-�TNTVճ�BV�Q[C�(c`�UWr��P�J��P�$0��SAsFE���V_SV�b�EXCLU��NnONL2��SY��*a&�OT�a'�HI�_V�4��B���_G *P0� 9�_z���p ��ASG�� +nrr�@6A@cc*b��G�#@E�V.i|Hb?fANNUN$0,.$fdID�U�2�SC@�`�i�a��j�f��!�pOGI$2,�O�$FibW$}�O�T9@�1 $DUMMYT��da��d�n�� � �E- ` ͑HE4(sg��*b�SAB��SUFFmIW��@CA=��c5�g6�abM�SW�E. 8̀KgEYI5���TM�100s�qA�vIN��#���b��/ D��H7OST_P!�r�`��ta��tn��tsp�pE�MӰV��� SBL�c ULI�0  A8	=ȳ�ј Tk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&�`DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F��!df�J� �q�C1�+6 H�bLL_DUs�~a3@{��3:���OTX"����s�"�0NOAUT5O�!7�p$)�$�*��c4�(�Cy��8�C, ��q&�L��� 8H *8�LH <6����c"� �`, `Ĭ�kª�q��@q��sq��~q��7���8��9��0����1���1̺1ٺ1�1��1 �1�1�2R(�2����2̺2ٺU2�2�2 �2�U2�3(�3��3���̺3ٺ3�3�3* �3�3�4(��a8��?��!9 <�9�&�z��I��1���M���QFE@'@� : y,6��Q? �@FP?9��5�9�E�@A�q�A� ;�p$TP�$�VARI:�Z���U�P2�P< ���TDe���K`Q���ܖ!��BAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�(H  ��P�Y�@|`�!>t ;E�4�sC�ST�D� D���c�<� 	 C��{��_���l����R  ���FORC�EUP?b��FLUS�`H�N>�F ��^�RD_CM�@E������� ��@vMP��REMr F�Q��1�`P���7Q
K4	NJ��5EFFۓ:�@I�N2Q��OVO�O{VA�	TROV���DTՀ�DTMX� ��@�
ے_P`H"p��CL��A_TpE�@�pK	_(�FY_T��v(��@%A;QD� �����`�!0tܑ0RQ��"�_�a����M�7�sCL�dρRIV'��{��EARۑIOFHPC�@����B�Bƅ�CM9@���R ��GCLF�e!DaYk(M�ap#5Tu�DG��� �%�aFsSSD �s? P�a(�!�1���P_�!�(J�!1��E�3�!3�+=5�&�GRA��7��@��;�PW��OyNn��EBUG_S�D2H�P{�_E �A �p����TERM`5Bi5U?��ORI#e0C�9SM_�P��e0�D�9TA�9E�9U}P\�F� -�A�{�AdPw3S@B$gSEG�:� EL{UwUSE�@NFIJ�B$�;1젎4�4C�$UFlP=�$,�|QR@��_G90qTk�D�~SNST��PAT����APTHJ3Q�E�p%B�`�'EC���ARx$P�I�aSHFTy��A�A�H_SHOR(Р꣦6 �0$�7P9E��E�OVR=��aRPI�@�U�b �Q�AYLOW���I�E"�r�A��?���ERV��XQ�Y��mG>@@�BN��U�a�R2!=P.uASYMH�.uFAWJ0G�ѡEq��A�Y�R�Ud>@��EC���EP;�uP;��6WOR>@M`��0SMT6�G3�G1R��13�aPAL@����`�q�uH � :���TOCA�`yP	P�`$OP����p�ѡ�`0O,��RE�`R4C�A�O�p낎Be�`R��Eu�h�A��e$P�WR�IMu�RR�_�cN��q=B I�&2H���p_ADD�R��H_LENG��B�q�q�q$�R��S��JڢSS��SK�N��u\��u̳�uٳS�E�A�jrS��MN�!K�����b����OLX��p�<���`ACRO3pJ� �@��X�+��Q��6�OUP3�b_�IX��a�a1��}򚃳� ��(��H��D��ٰ���氋�IO2S��D�����	�7��L $d��`Y!_O�FFr�PRM_���3�aTTP_�+�H:�M (|pOcBJ]"�p��$���LE~Cd���N � ��֑AB_�TqᶔS�`H�LVh�KR"uH�ITCOU��BG�LO�q���h�`����`��`SS� ����HW�#A:�O�ڠ<`INCPU>2VISIOW�͑���n��to��to�ٲ ��IOLN��P �8��R��p$S�Lob PUT_&n�$p��P& ¢���Y F_AS�"Q��$L������Q"  U�0	P4A��^���ZPHY��-��WP��UOI �#R ` �K����$�u�"pPpk���$���,���!UJ5�S-���;NE6WJOGKG̲'DIS����Kp���&�#T (�uAVF�+`��CTR�C
�FL�AG2��LG�dU� ���؜�13LG_SIZ����b�4�Xa��a�FDl�I`� w� m�_�{0a�^��c g���4�����Ǝ���x{0��� SCH_���a7�N�d�VW����E�"����4��U�M�Aљ`LJ�@�DAUf�EAU�p��d|��r�GH�ba���BO}O��WL ?��6 IT��y0�R;EC��SCR ܓ��D
�\���MARGm�!��զ ��d%�$����S����W����U� �JGM[�MN�CHJ���FNKEuY\�K��PRG���UF��7P��FWDv��HL��STP���V��=@��А�RS"��HO`����C9T�� b ��7�[�UL���@6�(RD� ����Gt��@PO��������M�D�FOCU��RG�EX��TUI��I��4�@�L� ����P����`��Pr��NE��CANA���Bj�VAILI�C�L !�UDCS_H!II4��s�O�(!"�S���S�缳!��BUFF�!Xj�?PTH$m�@��v`��D���AtrY�?P��j�3��`WOS1Z2Z3Z���� Z � ���[aEȤ��ȤID%X�dPSRrO��ԬzA�STL�R}�Y�&�� Y$E��C���K�&&8z�� [ LQ�� +00�	P���`#qdt
��U�dw<���_ \ �`4Г�\��Ѩ#�\0C4�] ��C�LDPL��UTRQ�LI��dڰ�)�$F�LG&�� 1�#�D���'B�LD�%�$�%ORGڰ5�2�PVŀ�VY8�s�T�r�$}d^� ���$6��$�%SB�`T� �B0�4�6RCLMC�4]?o?��9�9MI�p}d_� d=њRQ���DSTB�p� �;F�HHAX�R �JHdLEXCESHrD�BM!p�a`���/B�T�PC��`a�p=F_A7Ji��K�bOtH� K�db \�Q���v$MBC�L�I|�)SREQUI�R�R�a.\o�AXDESBUZ�ALt M���c�b�{P����2FANDRѧ`�`d;Ҙ2�ȺSDC��N�I�Nl�K�x`��X� N�&��aZ���UPS�T� ezrLO�C�RIrp�EX�<fA�p�9AAOD�AQ��f XY�OND�rMF,Łf �s"��}%�e/� ��A�FX3@IGG�� g ��t"��ܓhs#N�s$R�a%���iL��hL�v�@�D'ATA#?pE�%��tR��Y�Nh t_ $MD`qI}�A)nv� ytq�ytHP`��Pxu��(�zsANSAW)�yt@��yuD+��)\b���0o�i �@CUw�V�p 0XewRR2��j Du��{Q��7Bd$CALIIA@��G��2���RIN��"�<B:��INTE��Ck��r^�آXb]���_N�qlk���9�D���B�m��DIVFDH�@���qnI$V�,��S�$��$AZ�X�o�*�����oH �$B�ELT�u!ACC�EL�.�~�=�ICRC�� ���D�T��8�$PS�@�"L�@�r��#^�S�E�<� T�PATH3����I����ж�RO�A_@W��ڐ���2nC���4�_MG�$D�D��T���$FW��Rp9��I�4��D}E7�PPABN��ROTSPEE�[g�� J��[�C@�4��@$USE_d+�VPi��SYY����1 �aYN!@A��ǦOFF�qǡM�OU��NG���O9L����INC�tMa�6��HB��0HBENCS+�8q9Bp�4�FDm�IN�IԒ]�ౌB��VE��#�y�2�3_UP񕋳LOWL���p� B���Du�9B�``�x ����BCv�r�MOSI���BMOU��@�7P�ERCH  ȳOV��â
ǝ���� D�ScF�@MP����B� Vݡ�@y�j�LU0k��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A���Ԓ����N`�F�RT1I�A$��MOUЖЀHB�BS0�p7D5����ë�Z�DUM2�ԓS_BCKLSH_CԒk���� ϣ���=���ޡ �	ACLAL"q��1М�@��CHK� �S�RTY��^�%�E1Qq_�޴_UM��@�C#��SCL�0�r�LMT_J1_L��9@H�qU�EO�p�b�_�e�k�e�SPC��u���N�PC�N�Hz \P�2�C�0~"XT��CN_:�N9��I�SF!�?�V���U� /���ԒT���CB!�SH�:��E�E1TрT����y���T��P�A ��_P��_ � =������!�����J6 L�@��OG|�G�TORQU��ONֹ��E�R��H�LE�g_W2���_郠����I�IJ�I��Ff`xJ�1X�~1�VC3�0BD:B�1�@SB�JRKF9�0D�BL_SM��2M��P_DL2GR�V����fH�_��d���COS���LNH� �������!*,��aZ���fMY��_(�TH��)T�HET0��NK2a3���"��CB�&CB�CAA�B�"�0�!��!�&SB� 2N�%GTS�Ar�CI Ma�����,4#97#$DU���H\1�  �:Bk62�:AQ(rSf'$NE�D�`I��HB+5��$̀�!A�%��5�7���LPH�E�2���2SC% C%�2-&FC0JM&̀EV�8V�8߀LVJUV!KV/KV=KVKKVYKVgIH�8FRPM��#X!KH/KH=KUHKKHYKHgIO�<�O�8O�YNOJO�!KO/KO=KOKKO
YKOM&F�2�!+i%�0d�7SPBALA�NCE_o![cLE60H_�%SPc� &��b&�b&PFUL�C�h�b�g�b%p�1=k%�UTO_���T1T2�i/�2N ��"�{�t#�Ѱ`�0(�*�.�T��OÀ<�>v INSEG"�ͱ�REV4vͰl�DI�F�ŕ�1lzw��1m�0OBpq�я?��MI{���nLCHgWARY�_�AB��~!�$MECH�!�o ��q�AX��P�����7Ђ�`n 
p�d(�U�ROB���CRr�H���1(��MSK_f`�p� P �`_��R /�k�z�����1S�~��|�z�{���z��qIN�Uq�MTCOM�_C� �q  ����pO�$NO�REn����pЂ7r 8p GRe�u�SDZ�AB�$?XYZ_DA�1a���DEBUUq�������s z`$��COD�� L���p��$BUFIwNDX|��<��MORm�t $فUA��֐����r�<��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p} =�C�}pt�@b�D��FRIrӚ�T��RO@ \�E�}'���OPWO�Yq�v0Y�SY�SBU/@v�$SO!Pġd���ϪUΫ}p�PRUN����PA�D���rɡL�_O�Uo顢q�$^)�IMAG��w���0P_qIM��L�I�Nv�K�RGOVCRDt��X�(�P*�J�|��0L_�`]�L�0�RB1�����M��ED}��p J��N�PMֲ��c��w�SL�`q�w x $OVSL4vwSDI��DEX�@���#���-�V} *�N4�\#�B�2�G�4B�_�M�+��q|�E� x Hw���p��ATUSW����C�0o�s���BT�M�ǌ�I�k�4p��x�԰q�y Dw�!E&���@E�r��p7��жЗ�EXE���ἱ�����f q�z3 @w���UP'��3$�pQ�XN����������� �PG�΅{ h $S#UB����0_���!��MPWAIv�PL7ã�LOR�٠F\p�˕$RCVFA�IL_C��٠BW�D΁�v�DEFS}P!p | Lw����Я�\���UN!I+�����H�R�+�V}_L\pP����	P��p�}H�> �*��j�(�s`ȢN�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��G���PLI��p� � $ˀP_S�WI�pq�J_PL~��AL_ ���J��A��B��� C���D�$E���.�C_�U�� � � ���*��J3K0����TIA�4��5��6��MOM��������ˀB��AD��������6��PU� NR�������H��m��� A$PI�6 q��	�����K4��)6�U��w`��S/PEEDgPG�� ������Ի�4T��� � @��SA�Mr`��\�]��MOV_�_$�npt5�H�5���1���2��@������'�S�Hp�IN�'�@�+�����4($4+T+G�AMMWf�1'�$GGET`�p���Da�z��

pLIBR>ѺII2�$HI=�_�g�t��2�&E;��(A�.� �&LW�-6<��)56�&]��v�p��V���$PDCK���q��_?�����q�&���7��4����9+� �$_IM_SR�pD�s0�rF��r�rLE���aOm0H]��0�-ܬpq��PJqUR_SCRN�FA����S_SAVE_DX��dE@�NOa�CA A�b�d@�$q�Z�Iǡ s	�I� �J�K� ��� �H�L��>�"hq� �����ɢ�ɡ @bW^US�A�,M4���a��)q`��3�W@W�I@v�_�q�.MUA�o�� � $P9Y+�$W�P�vNG�{��P:��RA�0�RH��RO�PL������q� ��s'�X;�O�I�&�Zxe ���m��# p��ˀ�3s�O@�O�O�O�O�aa�_т� |��q�d@��.v ��.v��d@��[wFv��E���% ,r;B��E�|�tP����PMA�QUa ŉ�Q8��1٠QT�H�HOLW�QH�YS��ES��qU�E�pZB��Oτ�  ��Pܐ(�A�����v�!�t�O`�q���u�"���FA��IROG�����Q2���o��"��p��INFOBҁ�׃V����R�H�OI��� (�0SLEQ������Y��3����Á��P0O�w0���!E0N9U��AUT�A�COPY�=�/�'�
�@Mg�N��=�}1��4���� ��RG��Á͏��X_�P�$P;ख�`��W��P���@�������EXT/_CYC bHᝡ�RpÁ�r��_NA�e!А���RO�v`	�� � ���POR_�1�E.2�SRV �)_�I�DI��T_�k�}�@'���dЇ�����5���6��7��8i�H�S�dB���2�$��F�p��GPLeAdA
�TAR�Б@����P�2�裔d� ,��0FL`�o@YN���K�M��Ck��P�WR+�9ᘐ��D�ELA}�dY�pA�D�a� �QSK;IP4� �A�$�-OB`NT����P_$�M�ƷF@\bIp ݷ�ݷ�ݷd���� 빸��Š�Ҡ�ߠz�9��J2R� n��� 4V�EX� TQQ����TQ������� ��`�#�RDCN�V� �`��X)�R�p�����r��m$�RGEAR_� I9OBT�2FLG��fi&pER�DTC����|����2TH2NS�}� 1���G: T\0 ���uЉM\Ѫ`I�dG�R�EF�1Á� l<�h��ENAB��cTPE�04�]���� Y�]��ъQn#��*��"P�������2�Қ��@����������3�ҁ�'�9�K�]�o�� +��4�Ҝ������������5�ҝ�!�3�E�W�i�{��6�Ҟ������������
�7�ҟ-?Q(cu�8�Ҡ�������SMS�KÁ�l��a��E�kA��MOTE6�����@�݂TQ��IO}5�IS�tRr�W@��� �pJ���NU�������E�"$DSB_SIGN�1UQ�x��C\�TP��S23�2���R�iDEVICEUS�XRSR�PARIT��4!O�PBIT�QI�O?WCONTR+�TQX��?SRCU� MpS�UXTASK�3Nx�p�0p$TATU�PK��S�0������p_XPC)�$F�REEFROMS8	pna�GET�0��WUPD�A�2%F"�P� :��� !>$USAN�na8&����ERI�0�&RpRYq5*"_j@�qPm1�!�6WRK9�KD���6��QFR�IEND�Q�RUFxg�҃�0TOOL�6�MY�t$LEN�GTH_VT\�FCIR�pC�@ˀE> �+IUFIN-RM�ΕRGI�1ÐAITI�$GXñ3IvFG2v7G1���p3��B�GPR�p�1F�Oa_n 0��!RE��0p�53҅U�TC��3A�A�F �G(��":���e1n!��J�8 �%���%]��%�� 74��X O0�L
��T�3H&��8���%�b453GE�W�0�WsR�TD����T��M�����Q�T]�$V �2����1�а91T�8�02�;2k3�;3�:ifa�9-i�aQ0��NS��ZR$V��2B�VwEV�	V�B;�����&�S�`��F�"��k�@�2a�PS�E���$r1C��_3$Aܠ6wPR��7vMU�cS�t '�/89�G� 0G�aV`��p�d`���50�@��-��
25S�� �"�aRW����B�&�MN�AX�!�A:@�LAh��rTHIC¤1I���X�d1TF�Ej��q�uIF_C	H�3�qI܇7�Q�pG1RxV���]��:��u�_JF~�PR|ԀƱ�RVAT��� ��`���0R�榀DOfE��COU�Ա��AXI���O�FFSE׆TRIGNS���c����h������H�Y��IG#MA0PA�pJ�E��ORG_UNEV��J� �S������d �$CА��J�GROU����TqOށ�!��DSP���JOGӐ�#��_Pӱ�"O�q����@�&7KEP�IR��ܔ2�@M}R��AP�Q^��Eh0��K�SYS��q"K�PG2�BRAK�B��߄�pY�0=�d����`AD_������BSOC���N���DUMMY14�p@SV�PDE_�OP�#SFSPD�_OVR-���C���ˢΓOR٧3N�]0ڦF�ڦ��OV���SF��p���F�+�r!���CC��1q"L�CHDL��REC�OVʤc0��Wq@M������RO�#��Ȑ9_+��� @0�e@�VER�$OF�Se@CV/ �2WD��}��Z2���T�R�!���E_F�DO�MB_CM4���B��BL�bܒ#��adtVQR�$0pd���G$�7�AM5�`�� eŤ��_M;��"'����8$CA�'�E�8�8$HB�K(1���IO<�8����QPPA�������
��Ŋ����DVC_DBhC;��#"<Ѝ�r!S�1[ڤ�S�y3[֪�ATIOq 1q� ʡU�3���CABŐ�2�CvP���9P^�B���_� �S�UBCPU""ƐS �P �M�)0NS�c�M�"r�$HW_AC��U��S@��SA�A~�pl$UNITm�l_�AT���e�Ɛ�CYCLq�NEC�A���FLTR_2_FIO�7(��)&�B�LPқ/�.�_S[CT�CF_`�Fb�l���|�FS(!E�e�CHA�1��4�D°"3�RSD��$"}���#!�_Tb�PROX����� EMi_��ra�8!�a !�̹a��DIR0�RAOILACI�)RMr�CLO��C���Qq���#q�դ�PR=�S��A�pC/�c 	���FUNCq�0rRINP�Q�0��2�!3RAC �B ��[8���[WARn���#BL�Aq�A�����DAk�\���LD0���Q��q2eq�TI"r8��K�hPRIA�!r"AF��Pz!=�;���?,`�RK���MǀI�!�DF_@B�%1�n�LM�FAq@H�RDY�4_�P@R�S�A�0� �MUL�SE@���a ���ưt��m�m$�1$�1$1�o����� x*�EG� ����!cAR���Ӧ�09�2�,%� 7�AXE��RKOB��WpA��_l-���SY[�W!‎&S&�'WRU�/-1��@��STR������Eb� 	�%��J��A�B� ���&9�����O�To0 	$��A�RY�s#2��Ԓ�	�ёFI@��$LGINK|�qC1�aI_�#���%kqj2XYZ��t;rq�3�RC1j2^8'0B���'�4����+ �3FI���7�q����'���_Jˑ���O3�QO�P_�$;5���AT�BA�QBC��&�D�Uβ�&6��TURN߁"r�E11:�p��9GFL�`_���* �@�5�*7��Ʊ 1��� KŐM��&8����"r��ORQ ��a�(@#p=�j��g�#qXU�����mTOVEtQ:�M��i�� �U��U��VW�Z�A �Wb��T{�, ��@;� uQ���P\�i��UuQ�W`e�e�SERʑ
e	��E� O���UdAas��4S�/7����AX��B�'q ��E1�e��i��irp �jJ@�j�@�j�@�jP �j@ �j�!�f��i� �i��i��i��i� y�y�'y�7yTq�HyDEBU8�$ 32���qͲf2G �+ AB����رnSVS�7� 
#�d�� L�#�L��1W��1W�JA W��AW��AW�QW�@!�E@?D2�3LAB��29U4�Aӏ��C 7 o�ERf�5�� � $�@_ A6��!�PO��à��0#�
�_MRA�t�� d � T��ٔERR��=�;STY&���I��V�0��cz�TOQ�d�PL [ �d�"�� ?�w�!_ � pp`T)0���_V1Vr�aӔ����2ٛ2�E�����@�H�E���$W������V!��$�P��o�cI��aΣ�	 HELL_C�FG!� 5���B_BASq�SqR3��� a#QSb���1�%��U2��3��4��5���6��7��8���RaO����I0�0NL��\CAB+�����ACK4�����,��2@��&�?�_PU�CO,. U�OUG�P~ ��`��m�������TPհ�_KAR�l�_�R�E*��P���7Q�UE���uP����C�STOPI_AL 7�l�k0��h��]�l0GSEM�4�(�M4�66�TYN�SO���DIZ�~�A�����m�_TM�MANR�Q��k0E����$�KEYSWITCaH���m���HE��OBEAT��E- �LE~�����U��F�!Ĳ���B�O_HOuM=OGREFUP�PR&��y!� [�Cr��O��-ECOC�|�Ԯ0_IOCMWD<
�a�(k���� � Dh1���U�X���M�βgPgCFgORC��� ���m�OM.  � Q@�5(�U�#P, Q1��, 3��45�	�NPX_AS�t�� 0��ADD|���$SIZ���$VAR���TKIP/�.��A���M�ǐ��/�1�+ U"�S�U!Cz���FRIF��J�S���5Ԇ��NF�Ѝ� �� xp`SI��TE��C���CSGL��TQ2�@&����� ��OSTMT��,�P �&BWuP��SHO9W4���SV�$߻� �Q�A00�@Ma}���� ��P���&���5��6��U7��8��9��A�� O ���Ѕ�Ӂ���0��F��� G��0G�� �0G���@G��PG���1	1	1	1�+	18	1E	2��2���2��2��2��2���2��2��2��2���2	2	2	2�+	28	2E	3��3���3��3��3��3���3��3��3��3���3	3	3	3�+	38	3E	4�4���4��4��4��4���4��4��4��4���4	4	4	4�+	48	4E	5�5���5��5��5��5���5��5��5��5���5	5	5	5�+	58	5E	6�6���6��6��6��6���6��6��6��6���6	6	6	6�+	68	6E	7�7���7��7��7��7���7��7��7��7���7	7	7	7�+	78	7E��VP���UPDs� � �`NЦ�
��Y�SLOt�� � �L��d���A�aT�A�0d��|�ALU�:ed�~�CUѰjgF�!aID_L�ÑeH�I�jI��$FILcE_���d��$2��
�cSA>�� h�O��`E_BLCK���b$��hD_CPUyM�yA��c�o�dxb����R �Đg
PW��!� oqLA��S=�ts�q~tRUN�qst�q~t����qst�q~t ��T��ACCs���X -$�qLE�N;��tH��ph�_�I���ǀLOW_AXMI�F1�q�d2*�AMZ���ă��W�Im�8ւ�aR�TOR��p�g�D�Y���LAC�Ek�ւ�pV�ւ~�_�MA2�v�������T#CV��؁��T��ي �����t�V����V�IJj�R�MA�i�J���m�u�b����q2�j�#�U�{�t�K�JK���VK;���H���3f��J0����JJ��;JJ��AAL��ڐ(��ڐԖ4Օ5����N1���ʋƀW�L�P�_(�g����pr��� `�`GROU�w`��B��NFL�IC��f�REQUwIRE3�EBU�0�qB���w�2����p����q5�p�� \^��APPR��C}��Y�
ްEN٨CL9O7��S_M��H����u�
�qu�� ���MC�����9�'_MG��C�Co��`pM�в�N�BRKL�GNOL|�N�[�R���_LINђ�|�=�J����Pܔ�������� ���������6ɵ��̲8k����q���G� ��
��q)�<�7�PATH3�L�@B�L��H�wࡠ�J�CN�CA�Ғ�ڢ6B�IN�rUCV�4aZ��C!�UM��Y,���aE�p����������PAYLOAJ2L`R_A	N�q�Lpp����$�M�R_F2LS3HR��N�LOԡ��Rׯ�`ׯ�ACRL�_G�ŒЛ� ��H�j`߂$HM���FWLEXܣ�qJ�u� :���� ���������1�F1�V�j�@�R�d�v�������E����ȏ ڏ����"�4�q��� 6�M���~��U�g�y�$ယT��o�X��H� �����藕?����� ǟِݕ�ԕ�����%�7��JJ�� �� V�h�z���`A�T�採@�EL�� �S��J|�Ŝ�J�Ey�CTR��~�T�N��FQ��HAN/D_VB-���v`n�� $��F2M�X���ebSW�q��'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aDM)F�AW�Z`i�Aw�AA��X X�'pi�Dw��D��Pf�G�p�)S�Tk��!x��!N��DY�pנM�9$`%Ц� H��H�c�׎���0� ��Pѵڵ������������� ����1��R�6��QA'SYMvř���v���J���cі�_SH >��ǺĤ�ED����������J�İ%��C��IDِ�_VI��!X�2PV_UNIX�FThP�J��_R�5 _Rc�cTz�pT�V��@�@��İ�߷��U �Ԓ�����Hqpˢ���aEN�3�D)I����O4dD�`NJ�� x g"IJAAȱz�aabp�coc�`pa�pdq�a� ��/OMME��� �b4�RqAT(`PT�@� S��a7�;�Ƞ�@�h��a�iT�@<� $DUMMY9Q��$PS_��RF�C��$v p�p���Pa� XƠ����STE���S�BRY�M21_V�F�8$SV_ER�F�O��LsdsCLR�JtA��Odb`O��p � D �$GLOBj�_LO���u�q�cAp�r�@�aSYS�qADR�``�`TCH  �� ,��ɩb�W7_NA���7���SR���l ���
*?�&Q� 0"?�;'?�I)?�Y)�� X���h���x������) ��Ռ�Ӷ�;��Ív��?��O�O�O�DD�XS�CRE栘p��f��ST��s}y`�����/_HAΗq� TơgpTYP�b���G�aG�j��Od0IS_�䓀d�UEMd�# ����ppS�qa�RSM_�q*eUNEXCEP)fW�`S_}pM�x���g�z�8����ӑCOU��S��Ԕ 1�!�UE�&��Ubwr��PRO�GM�FL@$CUgpPO�Q��5��I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp��OUS�� �� @6p�v$BU�TTp�RpR�CO�LUMq�e��SE�RV5�PANE|H�q� � �@'GEU���Fy��?)$HELPõ)B/ETERv�)ෆ� ��A � ��0`��0��0ҰIN簊�c�@N��IH�1��_� �v��LN�r� �qprձ_ò=�$H���TEXl����F�LA@��RELVB��D`��������M��?,�ű�m�����"�USRVwIEW�q� <6p�`U�`�NFI<@;�FOCU��;�7PRI� m�`�Q�Y�TRIP�qm��UN<`Md� x#@p�*eWARN)e�6�SRTOL%���g��ᴰONCOR�N��RAU����T����w�VIN�Le�� $גPA�TH9�גCACH���LOG�!�LI�MKR����v���HwOST�!�bz�R��OBOT��d�IM>� �� ����Zq�Zq;�V�CPU_AVAIYL�!�EX	�!AN���q��1r��1r���1�ѡ�p� � #`C����@$�TOOL�$��_wJMP� ���e$SS�����VSHIF��Nc߃P�`ג�E�ȐR�����OSUR��Wk`RADILѮ��_�a��:�9a��`a�r���LULQ$OUTPUT_BM����IM�AB �@�r�TILSCO��C7����� ��&��3��A��@�q���m�I�2G�#�'��pLe�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM���F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? ��ZABC%��  $�"R���
ϐ�$$CLA}S������!�ϐϐ � VI�RT]��/ 0ABS�����1 5�� < �!F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZi{0�-�AXL�p��"�n63  �{tIN��qztPRE�����v��p�uLARMRECOV 9l�rwtNG�� .;	 A   �|.�0PPLIC���?5�p��Handlin�gTool o� �
V7.50P�/23-�  �P�f��
��_S�Wt� UP�!�� x�F0��t���A�0v� 86-4�� �it�y�� r2 �7DA5�� ��� Qf@<ϐo�Noneisͅ�˰ ��T����!LAex>�_l�V�uT��s9�UTO�"�Њt��y��HGAPON�
0g�1��Uh�D [1581�����̟ޟry����Q 1���p�,� 蘦���;�@��q_���"2 �c�.�H���D�HTTHKYX� �"�-�?�Q���ɯۯ 5����#�A�G�Y�k� }�������ſ׿1��� ��=�C�U�g�yϋ� �ϯ�����-���	�� 9�?�Q�c�u߇ߙ߫� ����)�����5�;� M�_�q������� %�����1�7�I�[� m����������!�� ��-3EWi{ ������ )/ASew�� ��/��/%/+/ =/O/a/s/�/�/�/�/ ?�/�/?!?'?9?K? ]?o?�?�?�?�?O�?��?�?O#O]���TO��E�W�DO_CL�EAN��7��CNMw  � ��__/_A_S_�DS�PDRYR�O��H	Ic��M@�O�_�_�_ �_oo+o=oOoaoso��o�o���pB��v �u���aX�t������>��PLUGG���G\��U�PRCvPB�@E��_�orOr�_7�SEGF}�K [mwxq�O�O���p��?rqLAP�_ �~q�[�m�������� Ǐُ����!�3�x�TOTAL�f yx�_USENU�p��� �H���B��RG_�STRING 1�u�
�M�n�S5�
ȑ_I�TEM1Җ  n 5�� ��$�6�H�Z� l�~�������Ưد����� �2�D�I�/O SIGNA�L̕Tryout Modeӕ�Inp��Sim�ulatedב�Out��OV�ERR�P = 1�00֒In c�ycl��בProg Abor���ב��Statu�sՓ	Heart�beatїMH� Faul��Aler'�W�E�W�iπ{ύϟϱ������� �CΛ�A����8� J�\�n߀ߒߤ߶��� �������"�4�F�X�8j�|���WOR{pΛ ��(ߎ����� ��$� 6�H�Z�l�~���������������� 2PƠ�X ��A{ ������� /ASew��p���SDEV[ �o�#/5/G/Y/k/ }/�/�/�/�/�/�/�/�??1?C?U?g?y?PALTݠ1��z? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�Op�O�O_�?GRI�` ΛDQ�?_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o2_l�R��a\_�o" 4FXj|��� ������0�B�<T��oPREG�>��  f���Ə؏����  �2�D�V�h�z��������ԟ���Z��$�ARG_��D ?�	���;���  	�$Z�	[O�]�O��Z�p�.�SBN�_CONFIG S;��������CII_SAVE  Z�����.��TCELLSET�UP ;�%HOME_IOZ�~Z�%MOV_��
�REP�lU�(�UTOBACKܠ���FRwA:\z� \�,z�Ǡ'`�z���\ǡi�INI�0z����n�MESS�AG���ǡC���ODE_D������%��O�4�n�PAUS�X!�;� ((O>��ϞˈϾϬ� ���������*�`߀N߄�rߨ߶�g�l TSK  wͥ�_��q�UPDT+��d�!�A�WSM_C5F��;���'�>-�GRP 2:�?�+ N�BŰA��%��XSCRD1�1
N7� �ĥĢ�� ��������*����� ��r�����������7� ��[�&8J\n���*�t�GROU�N�UϩUP_N5A�:�	t���_ED�17�
� �%-BCKEDT-�2�'K&�`���-t��z�q�q�z����2t1������q�k�(/��ED3/��/�.a/�/;/M/ED4�/t/)?��/.?p?�/�/ED5`??�?<?.�?O�?�?ED6O�?qO��?.MO�O'O9OED7�O`O_�O.�O\_�O�OED8L_,�_�^-�_ oo_�_�ED9�_�_]o�_	`-9o�oo%oCR _ 9]�oF�o�k�� � NO_DEL���GE_UNU�SE��LAL_?OUT �����WD_ABOR�ﰨ~��pITR_�RTN��|NO�NSk���˥C�AM_PARAM� 1;�!�
 8�
SONY X�C-56 234�567890 �ਡ@���?}��( А\��
���{����^�H�R5q�̹��ŏR5y7ڏ�Aff���KOWA SC�310M
�x��>��d @<�
� ��e�^��П\�� ��*�<��`�r�g��CE_RIA_I��!�=�F���}�z� ��_LeIU�]������<��FB�GP 1.��Ǯ�M�x_�q�0�C*  ��V��C1��9��@��iG���CR�C]��Ud��l��s��R��T���[Դm��v���������� C����(�����=�{HE�`ONFIǰ��B�G_PRI 1�{V���ߖπ�Ϻ����������C�HKPAUS�� ;1K� ,!uD� V�@�z�dߞ߈ߚ��� �������.��R�<�hb���O���������_MOR��� �^Biq-<���� 	 ��� ��*��N�`����䡑��?��q?;�;�����K��9�P��|�ça�-:���	�

��M��@�pU�ð��<��,~���DB���튒)�
mc:cpmi�dbg�f�:�L0���+¥�p�|/�  �(��(��� �sV>��pY�pZU��?􌐨�bUg�/���p�Uf�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����o=L���*MC��1����?43���1��t�īCz�  BHH�CPU�eB�_B�y�;��>C����CnY
K�E�?{hD]^Dْ?r���1�D��^�=G	���F��F���Cm	fF�O��F�ΫY	��,�&w�1���s����.�pT����BDw�M@x8��1�2�����g@D�p@�0�EY�1X�E�Q�EJP F��E�F� G���=F^F �E�� FB� �H,- Ge���H3Y��:�  �>�33 ����~  n8�~@F��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMO�FS�p�.8��)T}1��DE ��fF 
Q��;�(PG  B_<_��R�����	op6C4P�Y
s@ ]AQ�2s@�C�0B3�MaC{@@�*cw��UT�pFP?ROG %�z�o�oigI�q���v��ld�KEY_TBL � �&S�#� �	
��� !"�#$%&'()*+,-./01i��:;<=>?@A�BC� GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������vq���͓���������������������������������耇����������������������p`LCK�l4�p`��`STAT ��S_AUTO_DO����5�INDT_'ENB!���R�Q?��1�T2}�^�STO�Pb���TRLr`L�ETE��Ċ_S�CREEN ~�Zkcsc���U��MMENU �1 �Y  <�l�oR�Y1�[��� v�m���̟�����ٟ �8��!�G���W�i� �������ïկ��4� ��j�A�S���w��� ��迿�ѿ����T� +�=�cϜ�sυ��ϩ� ��������P�'�9� ��]�o߼ߓߥ���� ����:��#�p�G�Y� ����������$� ���3�l�C�U���y� ���������� ��	�VY)�_MANU�AL��t�DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[/ , 
�odP�&/~&lMZ�IdP�x@P@#ONTImMه� d�`&�
�e�MOTN�END�o�REC�ORD 1(�[8g2�/{�O��!�/ ky"?4?F?X?�(`? �?�/�??�?�?�?�? �?)O�?MO�?qO�O�O �OBO�O:O�O^O_%_ 7_I_�Om_�O�_ _�_ �_�_�_Z_o~_3o�_ Woio{o�o�_�o o�o Do�o/�oS�o L�o����@� ��+�yV,�c�u� �������Ϗ>�P�� ���;�&���q���� ����P�ȟ�^���� ��I�[����� ����$�6�������jTOLERENCwsB���L�͖ �CS_CFG �)�/'dMC�:\U�L%04dO.CSV�� c���/#A ��CH��z� //.ɿ��(S��RC_OUT �*���SGN� +��"��#��17-FEB-�20 18:57~015-JANp��0:51+ P/Vt�ɞ�/.���f�pa�m���PJPѲ��V�ERSION �Y�V2.0�.84,EFLOG�IC 1,� 	:ޠ=�ޠL���PROG_ENqB��"p�ULSk'� ����_WRS�TJNK ��"fE�MO_OPT_S�L ?	�#
 	R575/# =�����0�B����TO  �ݵϗ��V_F EX�d��%��PATH ;AY�A\����\�5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAqU��z�^"MSWX��.��4,#�Y�/�
!J�6%Z�I~m��$SBL__FAUL(�0�^9'TDIA[�1<��� ���1�234567890
��P��HZ l~������ �/ /2/D/V/h/�Z� P� ѩ� yƽ/��6�/�/�/? ?/?A?S?e?w?�?�?��?�?�?�?�?�,/�U3MP���� �A�TR���1OC@PM�El�OOY_TEM=P?�È�3F���G�|DUNI��.�Y�N_BRK 2�_�/�EMGDI_�STA��]��ENC�2_SCR 3�K7(_:_L_^_l& _�_�_�_�_)��C�A14_�/oo/oAo�Ԣ�B�T5�K� ϋo~ol�{_�o�o�o '9K]o� �������� #�5��/V�h�z��л` ~�����ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T���x��������� ү�����,�>�P� b�t���������ο� ���(�f�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������:� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ���*<N` r������� &8J\n� ���������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?��?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O��O__NoETMO�DE 16�5��Q �d�X
�X_j_|Q�PRROR�_PROG %fGZ%�@��_  �U�TABLE  �G[�?oo)oRjR�RSEV_NUM�  �`WP��QQY`�Q_AUT�O_ENB  ��eOS�T_NOna �7G[�QXb W *��`��`��`	��`d`+�`�o�o�o�dHISUc�aOP�k_ALM 18G[� �A��l�P+�ok}����r�o_Nb�`  G[��a�R
�:PTCP_VER !GZ�!�_�$EXTL�OG_REQv9�i\�SIZe�W��TOL  �aD�zr�A W�_BWD�p��xf́t�w_DI�� 9�5��d�T�asRֆS�TEP��:P�O/P_DOv�f�P�FACTORY_�TUNwdM�EATURE :�5�̀rQHa�ndlingTo�ol �� \sf�mEngli�sh Dicti�onary��ro�duAA V�is�� Mast�er����
EN�̐nalog I�/O����g.fd�̐uto Sof�tware Up�date  F �OR�matic Backup���H596,�g�round Ed�itޒ  1 H�5Camer�a�F��OPLG�X�ell𜩐II�) X�ommՐs�hw���com��c9o���\tp����pane��  o�pl��tyle �select��a�l C��nJ�Ցo�nitor��RD�E��tr��ReOliab𠧒6U�Diagnos(��푥�5528�u���heck Sa�fety UIF���Enhance�d Rob Se�rv%�q ) "�S�r�User F�r[�����a��xt�. DIO �f�iG� sŢ��en]dx�Err�LF�� pȐĳr됮� ܻ���  !��FCTN Menu`��v-�ݡ���TP �Inېfac� � ER JG�C�pבk Exczt�g��H558��igh-Spex��Ski1�  2�
P��?���mmuwnic'�ons���&�l�ur�ې��S�T Ǡ��con�n��2��TXPL��ncr�str�u����"FAT�KAREL C�md. LE�ua�G�545\��Ru�n-Ti��Env��d
!���ؠu++�s)�S/W���[�Licen3seZ��� 4T�0��ogBook(S�yڐm)��H54�O�MACROs,~\�/Offse��7Loa�MH�������r, k�Mec�hStop Pr�ot���� lic�/�MiвShif8����ɒMixx���)���xStS�Mo�de Switc�h�� R5W�Mo��:�.�� 74 H���g��K�2h�?ulti-T=�M����LN (P{os�Regiڑ�������d�ݐt Fun�ǩ�.������Num~����� l�ne��ᝰ Ad�jup�����  �- W��tatu�w᧒T�RD�Mz�ot��sco+ve U�9����3Ѓ�uest 492�*�o������62;�SNPX yb ���8 J7`���Libr��J�48���ӗ� �Ԅ�
��6O�� Part�s in VCCMt�32���	�{�ޤ�J990��/I�� 2 P��TM/ILIB��H���P�AccD�L�7
TE$TX�ۨ�7ap1S�Te����pkey��wգ��d��Unex�ceptx�mot�nZ���������є�� O���� �90J�єSP CSXC<�f��Ҟ�� Py�We}���P3RI�>vr�t��men�� ��iPɰa�����v�Grid�pla�y��v��0�)�H1��M-10iA(_B201 �2\�� 0\k/�Ascii�l�Т�ɐ/��Col��ԑGuaMr� 
�� /P-��ޠ"K��st{P�at ��!S�Cyqc�҂�orie�v�IF8�ata- quҐ�� ƶ��moH574��RL���am���Pb�HM/I De3�(b����PCϺ�Pas�swo+!��"PE�? Sp$�[���tp\��� ven��Tw��N�p�YELLO�W BOE	k$Ar�c��vis��3�*�n0WeldW�cGial�7�V#tѓOp����1y� �2F�a�portN�(�p�T1�T� ��� ��xy]�&T5X��tw�igj�1�� b� ct\�J�PN ARCPS�U PR��oݲO�L� Sup�2fi�l� &PAɰאcr=o�� "PM(�����O$SS� eвtex�� r���=�=t�ssagT��	P��P@�Ȱ�锱�rtW��H'>r��dpn��n1
�t�!� z ��as�cbin4psy�n��+Aj�M H�EL�NCL V�IS PKGS �PLOA`�MB ��,�4VW�RI�PE GET_V�AR FIE 3�\t��FL[�OO�L: ADD R�729.FD \Kj8'�CsQ�QE���DVvQ�sQNO �WTWTE��}PD�  �^��biRFwOR ��ECTn��`��ALSE A�LAfPCPMO-�130  M" �#h�D: HAN?G FROMmP��AQfr��R709� DRAM AV�AILCHECK�SO!��sQVPCS� SU�@LIMC�HK Q +P~dFF� POS��F�Q �R5938-12 CHARY��0�PROGRA �W�SAVEN`A�ME�P.SV��7��$En*��p?FU��{�TRC|� SH�ADV0UPDAT� KCJўRSTA�TI�`�P MUC�H y�1��IMQ� MOTN-00�3��}�ROBOG�UIDE DAU�GH�a���*�toQu����I� Šhd��ATH�PepMOV�ET�ǔVMXP�ACK MAY ?ASSERT�D���YCLfqTA�rB�E COR vr�*Q3rAN�pRC OPTIONSJ1�vr̐PSH-1k71Z@x�tcǠSU1�1Hp^9R!�Q�`C_T�P��'�j��d{tby app wa 5I�~d�P�HI���p�aTEL��MXSPD TIB5bLu 1��UB6@��qENJ`CE2�6�1��p��s	�ma�y n�0� R6�{�R� �Rtraf�f)�� 40*�p���fr��sysv�ar scr Jq7��cj`DJU���bH V��Q/�PS?ET ERR`J`� 68��PNDA�NT SCREEN UNREA��4'�J`D�pPA���p=R`IO 1���P�FI�pB�pGROUN�PD��G��R�P|�QnRSVIP !p��a�PDIGIT �VERS�r}BLo��UEWϕ P06s  �!��MAGp0�abZV�DI�`� SSUE�ܰ��EPLAN JO�T` DEL�pݡ#�Z�@D͐CALLOb�Q ph��R�Q�IPND��IMGޏR719��MN�T/�PES �pV:L�c��Hol�0Cq����tPG:�`C�M��canΠ��pg�.v�S: 3D �mK�view d2�` �p��ea7У�b� of �Py����ANNOT AC?CESS M��Ɓ�*�t4s a��lyok��Flex/�:�Rw!mo?�P�A?�-�����`n�p�a SNBPJ AUTO-�06f����TB��PIABL�E1q 636��P�LN: RG$�pl�;pNWFMDB�V�I���tWIT 9tx�0@o��Qui#0|�ҺPN RRS?p�USB�� t &� remov�@ �)�_��&AxEPFT�_=� 7<`�pP:��OS-144 ���h s�g��@O�ST� � CRASH DU 9���$P�pW� .}$��LOGIN���8&�J��6b046� issue 6� Jg��: Sl�ow �st��c (Hos`�c��z�`IL`IMPRWtSPOT:Wh:0\�T�STYW ./ЏVMGR�h�T0C�AT��hos��EP�q��� �O�S�:+pRTU' k�-�S� ����E:��ppv@�2�� t\hߐr��m ��all���0�  $�H� WA�͐��3 CNT0s T�� WroU�alarm���0s�d � �0SE1���r: R{�OMEBp����K� 55��RE�àSEst��g  �   �KAN�JI�no���I�NISITALI1Z-p�dn1weρ<�6�dr�� lx`��SCII L�f�ails w�� <��`�YSTEa���8o��Pv� IIH����1W�Gro>Pm 7ol\wpSh@�P���Ϡn cflx�L@АWRI �OF� Lq��p?�F�u�p��de-rel}a�d "APo �SY�ch�Abet�we:0IND t0$gbDO���r�y `�GigE�#�operabilf  PAbHi�H`���c�lead�\e�tf�Ps�r�OS� 030�&: fig��GLA )P ���i��7Np tps�wx�B��If�g�������5aE�a EXCE#dU�_�tP�CLOS��"ro�b�NTdpFaU�c�!���PNIO_ V750�Q1�8�Qa��DB ��P� M�+P�QED�D�ET��-� \rk~��ONLINEhSBUGIQ ߔĠi`�Z�IB�S apA�BC JARKY�Fq� ���0MILT�`� R�pNД �p�0GAR��D*pR8��P�"! jK�0c�T�P�Hl#n�a�Z�E V�� TASK�$VP2(�4`
��!�$�P�`WIBP�K05�!FȐB/���BUSY RUNN�� "�򁐈�2�R-p�LO�N�wDIVY�CUL���fsfoaBW �p���30	V���ˠIT`�a505�.�@OF�UNE�X�P1b�af�@�E���SVEMG� N�MLq� D0pCC_SAFEX 0c�0u8"qD �PET�`9N@�#J87����RsP�A'�M�K��`K�H GUN�CHG۔MECH��pMc� T�  y�, g@�$ ORY LEAKA�;��ޢSPEm�Ja��V�tGRIܱ�@�oCTLN�TRk��FpepR�j50�E�N-`IN�����p `�`�Ǒk!��T3/d\qo�STO�0A�#
�L�p �0�@�Q��АY�&�;pb1TO8pP�s���FB�@YpL`�`DU��aO�sHupk�t4 � P�F� �Bnf�Q�PSVG�N-1��V�SRS	R)J�UP�a2�Qx�#D�q l O��~�QBRKCTR5� ��|"-�r�<pc�j!�INVP�D ZO�� ��T`h#�Q�cHs�et,|D��"DU�AL� w�2*BRV�O117 A]�T�Nѫt�+bTa247`3��q.?��sAUz��i�B�comple�te��604.�� -�`hancZ�U� F��e8�'�  ��npJtPd!�q��`��� 5h596p�!5d�� "p �P�P�Q�0�P2�p�A�� xP��R(}\xPeJ� aʰI���E���1��p� j  �� xSt��^t �A�ApxP�q 5 sig��a��"AC;a��p
�bCexPb_p���.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o�dxPX�b]o2�� �cb�c��ixP�jupfrmp�dxP�o�`exe�ax�oFdxPtped}o���u`�cptlibxzxP�lcr�xrxP�\�blsazEdxP_fm�}gcxP�x���o�|sp�o�mc(��ob_jzop�u6�wQf��t��wms�1q���sld�)��jmc�o\�n��nuhЕ��|cst�e��>�pl�q�p�iwck���uv�f0uߒ��lvisyn�CgaculwQ�
E F  ! �Fc.fd�Qv�� �qw���Data Acquisi���nF�|1�RR631�`��TR�QDMCM� �2�P75H�1��P583xP1��7�1��59`�5�P5�7<PxP�Q����(0���Q��o pxP!/daq\�oA���@�� ge/�etd�ms�"DMER"؟,�pgdD���.��m���-��qaq.<᡾xPmo��h����f{�u�`13��MA�CROs, Sk�saff�@z����03��SR�Q(��Q6��1"�Q9ӡ�R�ZSh��P^xPJ643�@7ؠ�6�P�@�PRS�@����e �Q�UС PI�K�Q52 PTLqC�W��xP3 (��p/O��!�Pn ��xP5��03\s�fmnmc "M�NMCq�<��Q��\$AcX�FM���ci ,Ҥ�X����cdpq+�6
�sk�SK�xP�SH560,P���,�y�refp "GREFp�d�A�jxP6	�of�OFc�<g6y�to�TO_���<�ٺ���+je|�u��caxis2��xPE�\�e�q"IS�DTc��]�prax ��MN��u�b�isde܃h�\��w�xP! isba�sic��B� P�]��QAxes�R�6������.�(Ba�Q�ess��xP����2�D�@�z�atis���(�{����h��~��m��FMc��u�{�
ѩ�MNIS ��ݝ����x����xٺ��x� j75���Devic�� Interfac�R<ȔQJ754��� xP�Ne`��xP��ϐ2�б����d=n� "DNE���~
tpdnui5cUI��ݝ	bd�b�P�q_rsof�Ob
dv_ar�o��u�����stchkc��z	 8�(}onl��G!ffL+H�J(��"l"/�n�b���z�hamp��T�C2�!i�a"�59��S�q��0 (�+P�o��u�!2��xpc_2p�cchm��CHMqP_�|8бpevwsp��2쳌pcsF���#C SenxPa�cro�U·�-�R6�Pd�xPk�����p���gT�L��1d M �2`��8�1c4ԡ�3v qem��GEM,�\i(��Dgesnd��5���H{�}Ha�@s1y���c�Isu�xD��Fmd��I��7�4����u���AccuC�al�P�4� ��ɢ7TޠB0��6+6f�6��99\aFF q�SA(�U��2�
X�p�!�Bd��cb_�SaU=L��  �� ?��ܖto��otplus\tsrnغ(�qb�Wp��t���1���Tool (N. A.)�[K�7�Z�(P�m����bdfcls� k94��"K4p��qtpa=p� "PS9H�>stpswo��p�L7��t\�q���� D�yt5�4�q��w�qк�� �M�uk��rkey����s��}tҾsfeatu6�E!A��� cf)t\Xq��0���d�h5����LRC0�md�!�587���aR�(����d2V��8c?u3l\�pa3}H�&r-�Xu�b��t,�� �q "�q �Ot��~,���{�/��1c�}����y�p�r� �5���S�XAg�-�y����Wj874�-? iRVis���Queu�� Ƒ� -�6�1���(����u���tӑ����
��tpvtsn "VTSN�3C�+�� v\pRDV����*�/prdq\�Q�&�vstk=P����Ƥ�nm&_�դ�cl�rqν���get@�TX��Bd���aoQ8Ͽ�0qstr�D[�� ��t�p'Z����nqpv��@�enlIP�0��D!x�'�|���s1c ߸��tvo/�� 2�q���vb��� �q���!���h]���(� Contr{ol�PRAX�P�5��556�A@5m9�P56.@56@�5A�J69$@9�82 J552 IDVR7�hqA����16�H���La��� ��Xe�frl�parm.f�FRL�am��C9�@(F�����w6{����A��QJ643�� 50�0LSE�
_pVAR $�SGSYSC��R�S_UNITS ��P�2�4tA�TX.�$VNUM_OLD 5�1�xP{��50+�"�` Funct���5tA� }�(�`#@�`3�a0�cڂb��9���@H5נ� �P���(�A���� �۶}����ֻ}���bPRb�߶~ppr4�TPSPI�3�}�r�10�#;A� t��
`���1���96 �����%C�� Aف��=J�bIncr�	�� ��\���1o5q{ni4�MNINp	�xP�`���!��Ho�ur  r� 2�21 �?AAVM����0 ��TUP� ��J545� ��6162��VCAM  (��CLIO ��R6�N2��MSC "P ~�STYL�Cv�28~ 13\��NRE "FHR�M SCH^��DCSU%ORSsR {b�04 ��EIOC�1 �j 542 � o�s| � egis�t�����7�1~�MASK��934"7 ��O�CO ��"3�8Ļ�2���� 0 �HB��� 4�"39�N� Re�� �L�CHK
%OPLG�%��3"%MHCR&.%MC  ; 4? ���6 dPI�54��s� DSW%MDr� pQ�K!637�0Ƚ0p"�1�Р"4 ��6<27 CTNY K � 5 ���"I7��<25�%/�T�%OFRDM� �Sg!<��930 FB( �NBA�P� ( HL�B  Men�S�M$@jB( PVC ���20v��2HT�C�CTMI�L��\@PAC 116U�hAJ`SAI \@�ELN��<29s�?UECK �b�@�FRM �b�OR\���IPL��Rk0�CSXC ���V�VFnaTg@HTTsP �!26 ���G�@obIG{UI"%IPGS�r>� H863 qb�!8�07r�!34 �r�84 \so`! QLx`CC3 Fb�21��!96 rb!51� ���!53R% 1�!s3!��~�.p"9�js VATFUJ7�75"��pLR6^RP�WSMjUCTO��@xT58 F!80����1XY ta3!7�70 ��885&�UOL  GTSo
�<{` LCM �r| gTSS�EfP6 W�>\@CPE `��0cVR� l�QNL"���@001 imrb�c3 =�b�0����0�`6 w�b-P-� R-�b8n@5EW�b9 �Ґa� ����b�`ׁ�b2 20�00��`3��`4*5�`5!�c�#$�`�7.%�`8 h60�5? U0�@B6E�"aRp7� !Pr8� t�a@�tr2 'iB/�1vp3�vp�5 Ȃtr9Σ�a4r@-p�r3 F�Ⴐr5&�re`u��r7� ��r8�U�p9 �\h738�a�R/2D7"�1f���2&�7� �3 7)iC��4>w5Ip�NOr60 C�L�1bE6N�4 I�pyL�uP0��@N�-PJ8�N�8NeN�9 H�r`��E�b7]�|���88�Вࠂ9 2��a�`0�qЂ5�%U0O97 0��@1�0����1 (�q�3 5R���0���@mpU��0�0�7*��H@(q�\P"RB6�q124�b;��@����@06� x�3 pB/x�u ��x��6 H606�a1x� ��7 6 ����p�b155 �����7jUU162� �3 g��4�*�65 2e "_��P�4U1`���B�1���`0'�174� �q��P�E186g R ��P�7 ��P�8&�3 (�9o0 B/�s191�����@202��6� 3���A�RU2x� d��2 b2h`��4�᪂2�4����19v Q�2��u2Jd�Tpt2� ��H�a�2hP�$�5���!U2�p�p
�2�p��@!5�0-@��8 @��9��TX@�� �e5N�`rb26Af�2^R��a�2Kp��1y�b5(Hp�`
�5�0@�gqGA���a52ѐ�Ḳ-6�60ہ5� ׁ�2��8�E��9�EU)5@ٰ\�q5hQ`S*�2ޖ5�p\w�۲��pJ �-P��5�p1i\t�H�4��PCH�7j��phiw�@��P��x��559 ldu� P�D���Q�@������� �`.��P>�:��8�581�"�q�58�!AM۲T�Aw iC�a589��0@�x����5 �a��12׀0.�1���,��2����,�!P\h8���Lp ��,�7��6��0840\� ANRS 0C}A��p���{��ran��FRA��Д�е�� �A%���ѹ�Ҍ��� ��(����Ќ���� ����������ь�����$�G��1��ը���������� sxS�`q�  ������`64��M��iC/50T-H��`����*��)p46���� C��N����m7;5s֐� Sp���b46��v����Г/M-71?�7�З����42������C�2��-�а�70�r�E��/h����`O$��rD���c7c7C�q��Ѕ����L��/��2\imm7c7�g������`���(��e� ����"�������a0 r��c�T,�Ѿ�"��,�� ��x�Ex�m77t����k����5�����)�iC��-HS-�  B
_�>���+�Т�7U�]���Mh7
�s��7�������-9?�/260L�_������Q��������]�9pA/ @���q�S�х����h621��c��92����8��.�)92c0�g $�@�����)$��5$���pylH"O"
��21���t?�350����p��$�0�
�� �350!����0��9�U/0\{m9��M9A3�P��4%� s��3M$���X%u���"him�98J3����� i d �"m4~�103p�� <����h794̂�&R���H�0����\� ��g�5AU��՜��0�� �*2��00��#0�6�АՃ�է!07{r ���������kЙ@����EP �#������?��#!��;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?�ҽCD25L����u0�"l�2BL
#��B��\20�2_�r �re���X��1��N����A@��z��`C��pU��`��04H��DyA�\�`fQ���sU���\�5  ��� p�g�^t��<$85��p�+P=�ab1l��G1LT��lA8�!puDnE(�20T��qJ�1 e�bH85��h�b�Ռ�5[�16B@s��������d2�8�x��m6t!`Q ����bˀ���b#�(�6iB;S�p�!��3 � ��b�s��-`Є_�W8�_����6�I	$�X5�1�U85��R�p6S����/ �/+q�!�q��`�6o���5m[o)�m6s�W��Q�?��setC06p ��3%H�5��10p$����g/��JrH��  9��A�856���d�F�� ���p/2��@h�܅�✐)�5���̑v��(��m6���Y�H�ѝ̑m�6(�Ҝ��a6�DM����#-S�+��H2��� ��Ҽ�� �r̑���✐��l���p1����F���2�\t6h T6H����� ��'Vl���ᜐ�V@7ᜐ/����;3A7��p~S��������4�`圐�V���!3��2�PM[��%�ܖO�chn��ve�l5����Vq���_a�rp#��̑�.���2l_hemq$�.�'�6415���5����?����F�����5 g�L�ј[���1���𙋹1����M7NU�М��eʾ����Euq$D;��-�4��3&H�f�c�Ĝ�h�� ����u���〜���ZS�!ܑ4���M	-����S�$̑�ք �� 0��<�����.07shJ�H�v�� ��sF��S*󜐳����̑���vl�3�A�T��#��QȚ�Te��q�p�r����T@75j�5 �dd�̑1�(UL�&�(� ,���0�\�?���̑�a��� xSt ���a�e�w�2��(�2	�2�C��A/����\�+p�����21 9(ܱ�CL S���� B̺��7F���?�<�lơ1L����c�� ���u9�0����e!/q��O���9�K��r9 (��,�Rs���ז�5�G�m20Ac��i��w�2��:�0`�$��2�2l�0�@k�X�S� ,�ι2��hO���1!41w����2T@� _std ��G�y� �ң�H� jdgm����w0\�  �1L���	�P�~� W*�b��t 5�������3�,���E {������L��5\L��3�L�|# ~���~!���4�#�� O����h�L6A�������2璥����44�����[6\j4s��·���#��ol�E"w�8Pk��� ��?0xj�H1�1Rr��>��]�2a�2AHw�P ��2��|41�8 ��ˡ��{� �%�A<��� +�?�l��0�&�"��|�`Am1�2������3�HqB�� K�R��ˑb�W���Fs ���)�ѐ�!���ah�1����5��16�16C��C����0\imBQ��d���(�b��\B5�-���DiL���O�_�<��PEtL�E�RH�ZǠP8gω�am1l��u� ��̑�b�<����<�$�T�̑�F����I ̑�Dpb��X"�ᒢް�p� ���^�t��9�0\� j9�71\kckrcfJ�F�s�����c��e "CTME�r������!�a�`mai�n.[��g�`run}�_vc�#0�w��1Oܕ_u����bctme��Ӧ�`ܑ��j735�- K�AREL Use% {�U���J��(1���p� Ȗ�9��B@��L�9��7j�[�atk208 C"K��Kя��\��9��a��̹����c�KRC�a�o ��kc�qJ�&s�����Gr ſ�fsD��:y��s���A1X\j|хrdtdB�, ��`.v�q��� �sǑIf�Wfj�52�TKQuto� Set��J� �H5K536(�9i32���91�58(�i9�BA�1(�74O�,A$�(TCP A@k���/�)Y� ��\tpqtool�.v��v���! �conre;a#�C�ontrol R�e�ble��CNRE(�T�<�4�2���pD�)���S�552��q(g�� (򭂯4X��cOux�\sfu;ts�UTS`�i�栜���t�棂���? 6�T�!�SA OO+D6������ ���,!��6c+� igt�t6i��I0�TW8 ���la��vo58�o�bFå����i�Xh��!Xk�|0Y!8\m6e�!G6EC���v��6��@�������<16�A���A�6s����U�`g�T|ώ���r1�qR��˔Z4�T��� ��,#�eZp)g����<ONO0���uJ��t�CR;��F�a� xS�t�f��prdsuGchk �1��2&&$?���t��*D%$�r (�✑�娟:r��'��s�qO��<scr�c�C�\At�trld J"o�\�V�����Paylo�nf�irm�l�!�87���7��A�3ad �! �?ވI�?plQ��3��3"�q��x pl�`���d7��l�calC�uDu�8��;��mov������initX�:s8�O��a�r4 ��r6�7A4|�e Generatiڲ���q7g2q$��g R�� (Sh��c ,D|�bE��$Ԓ\P�:�"��4��4�4,�. sg��5�F�$d6"e�!p "�SHAP�TQ n7gcr pGC�a(��&"� ��"GDAL¶��r6�"aW<�/�$dataX:s�"tpad��[q�%tput;a__O7;a��o8�1�yl+s�r �?�:�#�?�5x�?�:	c O�:y O�:�IO�s`O%g�qǒ�?��@0\��"o�j92�;!�Ppl.Col�lis�QSkip #��@5��@J��D��@@\ވ�C@X�7���7�|s2��ptcls�LS�DU�yk?�\_ ets�`�< \�Q��@��d�`dcKqQ�FC;�b�J,�n��` (�D�4eN����T�{ ���'j(�c�q���/�IӸaȁ��̠H������зa�e\�mcclmt "�CLM�/��� ma�te\��lmpA�LM�?>p7qmc?����2vm�q��%�3s��_sv90�_x�_msu�2L^v_0� K�o�{in�8(|3r<�c_log8r��rtrcW�E �v_3�~yc롘�d�<�te��d�er$cCe� F	iρ�R��Q�?|�l�enter߄�|��(Sd��1�T�X�+fK�r�a99�sQ9+�5�r\t�q\� "FNDR����STD~n$LANG�Pgui��D⠓�S������sp�!ğ֙uf�ҝ�s����$�����e+�=����������������w�H�r\fn_�ϣ��$`x��tcpma��- �TCP�����R638 R�Ҡ��+38��M7p,���� ��$Ӡ�8p0Р�VS,�6>�tk��99�a�� B3���PզԠ��D�2�����UI��t���hq B���8��������p����re�ȿ��exe@4φ�B���e38�ԡG�rmpWXφ�var@�φ�3N�����vx�!ҡ��qҿRBT $c�OPTN as�k E0��1�R �MAS0�H593>/�96 H50�i�+480�5�H0��Dm�Q�K��7�0�g��Pl�h0ԧ�2�OR�DP��@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`m��b��7Г.f��u�d��r>��splayD�E����1w�UPDT |Ub��887 (��Di{���v�Ӛ�� �⧔��#�B��㟳��o  ����a������60q��B���>��qscan��B���ad@�������q`�䗣�#���8��`2�� vlv�䀃Ù�$�>�b���!y S��Easy/���Util��룙�511 J�����9R7 ��Nor֠��inc),<6Q�� �`c��"4�[���G986FVRx S1o����q�nd6��� �P��4�a\ (��
  �������d��K�b9dZ���men7���o- Me`tyF���Fb�0�TUa�'577?i3R��\�5�u?��!� n���f������l\mh�Ц�űE|hmn�	��<!\O���e�1�� l!��y��Ù�\|p����B�����mh�@��:. aG!���/�t�55�`6�!X�l�.us��|Y/k)ensubL�
��eK�h�� �B \1;5g?y?�?�?D��?�*rm�p�?Ktbox O2K|?�G��C?A%ds���?1ӛ#� �TR��/��P� 4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ă�Q23t.�P׀al��Pr+OP517��#IN0a��Q(}g�N�PESTf3ua�P B�l�ig�h�6�aq���P � xS���`  n�0mb�umpP�Q969�g�69�Qq��P0�b�aAp�@Q� BOqX��,>vche�s�>vetu㒣=w/ffse�3����]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q<t�waǂ tp�Q҄T�aror Rec�ov�b�O�P�642����a�q��a�⁠QErǃ�Qry�з`�P'�T�`�aarൄ����	{'�pak7971��71��m0���>�pjot��P�Xc��C�1�adb -v�ail��nag��<�b�QR629�a�Q���b�P  �
�  �P��$�$CL[q �����������$�PS_DIGI�T��� "�!�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv��������*璬�1:PRODUC�T�Q0\PGST�K�bV,n�9�9�\���$�FEAT_IND�EX��~��� 搠ILECOMP ;���)��"��SETUP2 <����  N� !�_AP2B�CK 1=� � �)}6/E+%,/i/��W/�/~ +/�/O/�/s/�/?�/ >?�/b?t??�?'?�? �?]?�?�?O(O�?LO �?pO�?}O�O5O�OYO �O _�O$_�OH_Z_�O ~__�_�_C_�_g_�_ �_	o2o�_Vo�_zo�o o�o?o�o�ouo
�o .@�od�o�� �M�q���<� �`�r����%���̏ [�������!�J�ُ n�������3�ȟW�� ����"���F�X��|� ���/���֯e����� �0���T��x���� ��=�ҿ�s�ϗ�,Ϡ��9�b�� P/� 2) *.VRiϳ�!�*�����0�����PC�7�>!�FR6:"�c��χ��T��߽߀Lը��ܮx���G*.F��>� �	N��,�k��ߏ��STM �����Qа����!�iPend�ant Pane	l���H��F���4�p�����GIF��������u����JPG&P��<�����	PANELO1.DT���� �����2�Y@�G��
3w������//�
4 �a/�O///�/��
TPEINS.�XML�/���\��/�/�!Custo�m Toolba�r?�PASS�WORD/�F�RS:\R?? %�Passwor�d Config �?��?k?�?OH�6O �?ZOlO�?�OO�O�O UO�OyO_�O�OD_�O h_�Oa_�_-_�_Q_�_ �_�_o�_@oRo�_vo o�o)o;o�o_o�o�o �o*�oN�or� �7��m��&� ��\�����y��� E�ڏi������4�Ï X�j��������A�S� �w�����B�џf� ������+���O���� �����>�ͯ߯t�� ��'���ο]�򿁿� (Ϸ�L�ۿpς�Ϧ� 5���Y�k� ߏ�$߳� �Z���~�ߢߴ�C� ��g�����2���V� ���ߌ���?���� u�
���.�@���d��� ����)���M���q��� ��<��5r� %��[�& �J�n��3 �W���"/�F/ X/�|//�/�/A/�/ e/�/�/�/0?�/T?�/ M?�??�?=?�?�?s? O�?,O>O�?bO�?�O O'O�OKO�OoO�O_ �O:_�O^_p_�O�_#_ �_�_Y_�_}_o�_�_�Ho)f�$FILE�_DGBCK 1�=��5`��� ( ��)
SUMMAR�Y.DGRo�\M�D:�o�o
`D�iag Summ�ary�o�Z
CONSLOG�o�o�a�
J�aConsole logK��[�`MEMCH�ECK@'�o��^qMemory �Data��W��)�qHADO�W���P��sS�hadow Ch�angesS�-c-���)	FTP�=��9����w`qm�ment TBD�׏�W0<�)ETHERNET̏��^�q�Z��aEthernet bp�figurati�on[��P��DCSVRFˏ��Ïܟ�q�%�� verify allߟ�-c1PY���DI�FFԟ��̟a��p{%��diffc���q��1X�?�Q��� ����X��CHGD��¯ԯ�i��px��� ���2p`�G�Y�� ��� �GD��ʿܿq���p���Ϥ�FY3ph�O�a��� ��(�GD������y���p�ϡ�0�UP?DATES.�Ц�~�[FRS:\������aUpdates List����kPSRBWLD'.CM.��\��B���_pPS_ROBOWEL���_���� o��,o!�3���W��� {�
�t���@���d��� ��/��Se��� ��N�r�  =�a�r�& �J���/�9/ K/�o/��/"/�/�/ X/�/|/�/#?�/G?�/ k?}??�?0?�?�?f? �?�?O�?OUO�?yO O�O�O>O�ObO�O	_ �O-_�OQ_c_�O�__ �_:_�_�_p_o�_o ;o�__o�_�o�o$o�o Ho�o�o~o�o7�o 0m�o� ��V �z�!��E��i� {�
���.�ÏR����� �����.�S��w�� ����<�џ`������ +���O�ޟH�������8���߯n����$�FILE_��PR����������� �MDONLY 1=4�~� 
 ��� w�į��诨�ѿ���� ���+Ϻ�O�޿sυ� ϩ�8�����n�ߒ� '߶�4�]��ρ�ߥ� ��F���j�����5� ��Y�k��ߏ���B� ����x����1�C��� g������,���P��� ������?��Lu~�VISBCKR�|<�a�*.VD||�4 FR:\���4 Visi�on VD file� :Lbp Z�#��Y�} /$/�H/�l/�/ �/1/�/�/�/�/�/ ? �/1?V?�/z?	?�?�? ??�?c?�?�?�?.O�? ROdOO�OO�O;O�O �OqO_�O*_<_�O`_��O�__%_�_�MR_GRP 1>4��L�UC4  ;B�P	 ]�o�l`�*u����RHB ���2 ��� �?�� ���He�Y �Q`orkbIh�oJd�o�Sc�o�oLP��ELcPxJ�]ߘF�5U�aS�3��o�o E��]�F�nE�wB�.��99�ʓ>�E}�A%%Az�-�lq?�R4Az���xq0~�� F�@ �r�d�a}J���NJk�H9��Hu��F!���IP�s}?��`�.9�<9��896�C'6<,6\b�1�,.�g�0R���^x�PA����� |�ݏx���%��I� 4�F��j�����ǟ�� �֟��!��E�`rv�UBH�P �~М������W
6�P=?��PQ��˯�o��oB��P5���@'�33@���4�m�^,�@UUU��U�~�w�>u.�?!x�^��ֿ���3���=[z�=����=V6<�=��=�=$q���~��@8�i�7G��8�D��8@9!��7ϥ�@Ϣ���cD��@ D�� CYϫo��C��P��P'�6��_V� m�o�� To��xo�ߜo����� �A�,�e�P�b��� �����������=� (�a�L���p������� ��^�������*��N 9r]����� ���8#\n Y�}������ �/ԭ//A/�e/P/ �/p/�/�/�/�/�/? �/+??;?a?L?�?p? �?�?�?�?�?�?�?'O OKO6OoO�OHߢOl� �ߐߢ��O�� _��G_ bOk_V_�_z_�_�_�_ �_�_o�_1ooUo@o yodovo�o�o�o�o�o �oNu �������� �;�&�_�J���n��� ����ݏȏ��%�7� I�[�"/�描����� ٟ�������3��W� B�{�f�������կ�� �����A�,�e�P� b��������O�O�O ��O�OL�_p�:_�� ���Ϧ��������'� �7�]�H߁�lߥߐ� �ߴ�������#��G� 2�k�2��Vw���� �������1��U�@� R���v����������� ��-Q�u� ��r��6�� )M4q\n� �����/�#/ I/4/m/X/�/|/�/�/ �/�/�/?ֿ�B?� f?0�BϜ?f��?���/ �?�?�?/OOSO>OwO bO�O�O�O�O�O�O�O __=_(_a_L_^_�_ �_�_���_��o�_o 9o$o]oHo�olo�o�o �o�o�o�o�o#G 2kV{�h�� �����C�.�g� y�`����������Џ ���?�*�c�N��� r��������̟�� )��M�_�&?H?���? ���?�?�?����?@� I�4�m�X�j�����ǿ ���ֿ����E�0� i�Tύ�xϱϜ����� ����_,��_S���w� b߇߭ߘ��߼����� ��=�(�:�s�^�� ���������'� 9� �]�o����~��� ����������5  YDV�z��� ���1U@ yd��v����� /Я*/��
/�u/� �/�/�/�/�/�/�/? ?;?&?_?J?�?n?�? �?�?�?�?O�?%OO IO4O"�|OBO�O>O�O �O�O�O�O!__E_0_ i_T_�_x_�_�_�_�_ �_o�_/o��?oeowo �oP��oo�o�o�o �o+=$aL�p �������'� �K�6�o�Z������ ɏ��폴� ��D� / /z�D/��h/ş�� �ԟ���1��U�@� R���v�����ӯ���� ��-��Q�<�u�`� ��`O�O�O���޿� �;�&�_�J�oϕπ� �Ϥ��������%�� "�[�F��Fo�ߵ��� �ߠo��d�!���W� >�{�b�������� ������A�,�>�w� b����������������=��$FN�O ����\�
�F0l q  FL�AG>�(RRM�_CHKTYP � ] ��d ��] ��OM� _�MIN� 	����� �  XT S�SB_CFG �?\ ����O�TP_DEF_O/W  	��,�IRCOM� >��$GENOVRD7_DO��<�l�THR� d�d�q_ENB] �qRAVC_GR�P 1@�I X(/ %/7//[/ B//�/x/�/�/�/�/ �/?�/3??C?i?P? �?t?�?�?�?�?�?O OOAO(OeOLO^O�O.oROU�F\� �,�B,�8�?���O�O��O	__���  DaE_�Hy_�\@@m_B�=�vR/��I�O�WSMT�G�SU�oo&oRHOST�C�1H�I� Ĺ�zMSM��l[bo�	1�27.0�`1�o  e�o�o�o #z�oFXj|�l6�0s	anonymous�����F�ao�&�&��o�x��o������ ҏ�3��,�>�a� O����������Ο�U %�7�I��]����f� x��������ү��� �+�i�{�P�b�t��� ���������S� (�:�L�^ϭ�oϔϦ� �������=��$�6� H�Zߩ���Ϳs����� ������ �2���V� h�z��߰������� ��
��k�}ߏߡߣ� ���߬���������C� *<Nq�_�� ����-�?�Q�c� eJ��n���� ���/"/E� X/j/|/�/�/� %'/?[0?B?T?f? x?��?�?�?�?�?? E/W/,O>OPObO�KDa�ENT 1I�K� P!�?�O  �P�O�O�O�O�O#_ �OG_
_S_._|_�_d_ �_�_�_�_o�_1o�_ ogo*o�oNo�oro�o �o�o	�o-�oQ u8n����� ���#��L�q�4� ��X���|�ݏ���ď�֏7���[���B�?QUICC0��h�z�۟��1ܟ��ʟ+��2,���{�!?ROUTER|�X��j�˯!PCJO�G̯��!19�2.168.0.�10��}GNAME� !�J!RO�BOT�vNS_C�FG 1H�I ��Aut�o-starte�d�$FTP�/ ���/�?޿#?��&� 8�JϏ?nπϒϤ�ǿ ��[������"�4ߵ& ����������濜��� �������'�9�K�]� o����������� ��/�/�/G���k��� �������������� 1T���Py�� ���"�4�	H- |�Qcu�VD� ���/�;/M/ _/q/�/����/
/ �/>?%?7?I?[?*/ ?�?�?�?�/�?l?�? O!O3OEO�/�/�/�/ �?�O ?�O�O�O__ �?A_S_e_w_�O4_._ �_�_�_�_oVOhOzO �O�_so�O�o�o�o�o �o�_'9Kno �o�����o*o <oNoP5��oY�k�}� ����pŏ׏���� 0���C�U�g�y���_��T_ERR J�;�����PDUSI�Z  ��^P�����>ٕWRD �?z���  �guest ���+�=�O�a�s�*��SCDMNGRPw 2Kz�Ð���۠\��K��� 	P01.�14 8�q  � y��B    ;�����{ �����������������������~ �ǟI�4�m�X��|��  i�  �  
����� ����+��������
����l�.x��
��"�l�ڲ۰s��d�������_G�ROU��L�� e��	��۠07K�QUPD  ����PČ�TYg������TTP_A�UTH 1M��� <!iPen'dan���<�_��!KAREL�:*�����KC�%�5�G��VISION SETZ���|��Ҽߪ��� ������
�W�.�@����d�v���CTRL� N�������
� �.FFF9�E3���FRS�:DEFAULT��FANUC� Web Server�
���� ��q��������������WR_CONFI�G O�� ����IDL_CP�U_PC"��B���= �BH#M�IN.�BGNR_IO��� ���% �NPT_SIM_�DOs}TPM�ODNTOLs >�_PRTY�=�!OLNK 1P���'9K�]o�MASTE�r �����O_CFG��UO����CYCLE���_ASG 1Q���
 q2/D/V/ h/z/�/�/�/�/�/�/��/
??y"NUM����Q�IPC�H��£RTRY�_CN"�u���SGCRN������1 ���R�����?��$J23_�DSP_EN������0OBPROqC�3��JOGV��1S_�@��8G�?�';ZO'??0C�POSREO�KANJI_�ϠuH�A#��3T ���E<�O�ECL_LM B2�e?�@EYLOGG+IN��������LANGUAGE� _�=� ,}Q��LG�2U���+�� �x�����P�C � �'0������MC:\�RSCH\00\�˝LN_DISP V������f�TOC�4Dz\�A�SOGBOOK W+��o���o�o���Xi�o�o�o�o�o~}	x(y��	ne�i�ekEl�G_BUFF 1%X���}2�� ��Ӣ������ '�T�K�]��������� ��ɏۏ���#�P���ËqDCS Z>xm =���%|d�1h`���ʟܟ�g�I�O 1[+ �?'����'�7�I�[� o��������ǯٯ� ���!�3�G�W�i�{�@������ÿ׿�El /TM  ��d��#� 5�G�Y�k�}Ϗϡϳ� ����������1�C߀U�g�yߋߝ߈t�S�EV�0m�TYP�� ��$�}��ARS"�(_�s�2F�L 1\��0� ��������������5�TP<P���>DmNGNAM�4�U��f�UPS`GI�5�A�5s�_LO{AD@G %j{%@_MOV�u�����MAXUALRMB7�P8��y��D�3�0]&q��Ca]s�3�~�� 8@=@]^+ طv	��+V0+�P�A5dƋr���U ������E (iTy���� ���/ /A/,/Q/ w/b/�/~/�/�/�/�/ �/??)?O?:?s?V? �?�?�?�?�?�?�?O 'OOKO.OoOZOlO�O �O�O�O�O�O�O#__ G_2_D_}_`_�_�_�_ �_�_�_�_o
ooUo 8oyodo�o�o�o�o�o��o�o�o-��D_L?DXDISA^��� �MEMO_AP�X�E ?��
 �0y�����������ISCw 1_�� � O����W�i����� Ə�����}��ߏD� /�h�z�a�������� ������@���O� a�5������������ u��ׯ<�'�`�r�Y� �����y�޿�ۿ� ��8Ϲ�G�Y�-ϒ�}� �ϝ�����m�����4���X�j�#�_MST�R `��}�SC/D 1as}�R��� N��������8�#�5� n�Y��}������� �����4��X�C�|� g��������������� 	B-Rxc� ������ >)bM�q�� ���/�(//L/ 7/p/[/m/�/�/�/�/ �/�/?�/"?H?3?l?�W?�?{?�?�?�?n�MKCFG b����?��LTARMu_�2cRuB� �3WpTNBpM�ETPUOp�2�����NDSP_CMNTnE@F�E��' d���N�2A��O�D�EPOSCF��G�NPSTOL� 1e-�4@�<#�
;Q�1;UK_YW 7_Y_[_m_�_�_�_�_ �_�_o�_oQo3oEo��oio{o�o�a�ASI�NG_CHK  y�MAqODAQ2C�fO�7J�eDEV� 	Rz	MC}:'|HSIZEn@�����eTASK �%<z%$123456789 ���u�gTRIG 1]g�� l<u%����3���>svvY�Paq��kEM_I�NF 1h9G� `)AT&FV0E0(����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ ߏP��t�������]� ί�����(�۟� ^��#�5�����k�ܿ � ϻ�ů6��Z�A� ~ϐ�C���g�y����� ���2�i�C�h�ό� G߰��ߩ��ߙϫ�� ������d�v�)ߚ��� ��y��������<� N��r�%�7�I�[��� ���9�&��J�[�g��>ONIwTOR�@G ?;{�   	EX�EC1�3�2�3��4�5��p�7*�8�9�3�n� R�R�RR RR(R4R@�RLR2Y2e2�q2}2�2�2��2�2�2�3�Y3e3��aR_�GRP_SV 1�it��q(�a>��0��Z����h�1�ȇ$�1�'x~q_DCd~��1PL_NAME� !<u� �!�Default� Persona�lity (from FD) �4�RR2k! 1j)TEX)TH��!�AX d�?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O�O�Ox2-?�O�O�O __0_B_T_f_x_�b<�O�_�_�_�_�_�_�o o2oDoVoho&xR�j" 1o�)&0\��b, �9��b~�a @D�  �a?��c�a?�`�a�a�A'�6�ew;��	l�b	 �xJp��`�`	p ��< �(p� ��.r� K�K� ��K=*�J����J���J�V��kq`q�P�x�|5p@j��@T;f�r�f��q�acrs�I�o����p���p��r�ph}�3���o�  ��>���ph�`z��;꜖"�Jm�q� H�N��ac���d�w��  � W P� Q� �� |  а�m�Ə�i}	'� � ��I� � � ����:�����È=����(�ts�a	���I  �n @H� i~�ab�Ӌ�b�w���urN0��  '�Ж�q�p@2�@����r�q5��C�pC0C�@ �C����`
S�A1]w@B�V~�X�
nwB0h�A��p�ӊ�p@����aDz���֏���Я�	�pv�( �� -��I��0-�=��A�a�we_q��`�p �?�f�f ��m��� ����Ƽuq@tݿ�>1�  P�apv(�`ţ� �=�qxst��?���`�x`�5p<
6b<�߈;܍�<��ê<� <G�&P�ό�AO���c1��ƍ�?fff�?O�?&��qt@��.�J<?�`��wi4����dly �e߾g;ߪ�t��p� [ߔ�߸ߣ����� �`���6�wh�F0 %�r�!��߷�1ى�����E�� E�~O�G+� F�!� ��/���?�e�P���t�,��lyBL�cB��E nw4�������+��R ��s�����<����h�Ô�>��I�m0Xj���A�y��weC������Ƀ�#/*/c/N/wi�6����v/C�`� CCHs/`
=$�p�<!��!��ܼ�'�3A��A�AR1A�O�^?�$�?���5p±
=�ç>����3�W
=�#�]��;e��?������{����<��>(�B��u��=B0�������	�R��zH�F�G����G��H��U`E���C��+��}I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0w/O*OONO9O rO]O�O�O�O�O�O�O �O_�O8_#_\_G_�_ �_}_�_�_�_�_�_�_ "oooXoCo|ogo�o �o�o�o�o�o�o	 B-fQ�u�� �����,��P� b�M���q�����Ώ�� �ݏ�(��L�7�p� [������ʟ���ٟ ���6�!�Z�E�W���:#1($1��9�K����ĥ%��x��Ư!3�8��<�!4Mgs���,�IB+8�J��a?���{�d�d������ȿ���ڼ%P8�P�=:GϚ�`S�6�h�z���R��������������  %�� ��h�Vߌ�z� ��&�g�/9�$�������7����A�S�e�w�  ��������������2 wF�$�&Gb���������!C����@���8�����F�� DzN��� F�P D�������)#B�'9�K]o#?��ͫ@@v
��8��8��8�.
 v���!3 EWi{�����:� ��ۨ��1��$MSKCFMAP  ��� ����(.�ONREoL  �!�9��EXCFEN�BE'
#7%^!FN�Ce/W$JOGOV�LIME'dO S"d��KEYE'�%��RUN�,�%��SFSPDTY�0g&P%9#SIGN|E/W$T1MOT�/�T!�_CE_G�RP 1p��#\x��?p��?�? �?�?�?O�?OBO�? fOO[O�OSO�O�O�O �O�O_,_�OP__I_ �_=_�_�_�_�_�_o�o�_:o�TCO�M_CFG 1qB	-�vo�o�o
Va__ARC_b"��p)UAP_CPL��ot$NOCHEC�K ?	+ �x�%7I[ m���������!�.+NO_WAIT_L 7%S2�NT^ar	+��s�_ERR_12s	)9�� ,ȍޏ���x���&��dT�_MO��t��, �Q/�p�8�PAR�AM��u	+���a�ß'g{�� =�?�345678901��,��K�]� 9�i�������ɯۯ��&g�����C��c�UM_RSPAC�E/�|����$ODRDSP�c#6p(�OFFSET_C�ART�o��DIS�ƿ��PEN_FI�LE尨!�ai��`O�PTION_IO��/��PWORK kve7s# �� V�ؤ��p�4�p��	 ���p��<����RG_DSBL'  ��P#������RIENTTOD ?�C�� !l����UT_SIM_ED$�"���V��?LCT w}�h��iĜa[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ���� ��ڐH(���H3k7HS�M5G�22G�?��Gp
͜��'f�/-,ڐCR�>�D!�M#{Z/���3�����4y H "�c/u/�/�0B_����=jc��t�!�/ �/�"t32���~�/6  ��UP%�Q%��%�|T���S62�q?'e	'�� � �2I�� �  ��+==��ͳ?�;	��h	�0�I  �n @�2�.���Ov;��ٟ?&gN�]O  ''�uD@!:� C�C�@F#H!��/�O�O sb
�T��@�@��@$�e0@B�QA�0Y�v: �13Uwz $oV_�/z_e_�_�_	���( �� -�2�1�1ta�UDa�c���:A-���~.  �?�ff���[o"o�_U�`oXâ0A8���o�j>�1  Po�V(���eF0��f�Y���L�?˙���xb0@<
�6b<߈;����<�ê<�? <�&�,�/aA�;r�@Ov0P?offf?�0?&ipޘT@�.{r�J<?�`�u#	�B dqt�Yc�a�Mw �Bo��7�"�[�F� �j�������ُ� ���3����,���~(�E�� E��3?G+� F��a�� ҟ�����,��P�(;���B�pAZ�>� �B��6�<OίD���P� �t�=���a�s������6j�h��7o��>�S��O�����Fϑ�A�a�_���C3Ϙ�/�%?��?Ƀ��������#	���P �N||CH����Ŀ������@�I�_�'�3A��A�AR1A�O�^?�$�?������±
=�ç>����3�W
=�#� U���e���B��@���{����<����(�B��u��=B0�������	��b�H�F�G����G��H��U`E���C��+��I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻�������� � �9�$�]�H�Z��� ~�������������# 5 YD}h�� �����
C .gR����� ��	/�-//*/c/ N/�/r/�/�/�/�/�/ ?�/)??M?8?q?\? �?�?�?�?�?�?�?O �?7O"O[OmOXO�O|O �O�O�O�O�O�O�O3_:Q(������b���gUU��xW_i_2�3�8��_<�_2�4Mgs�_�_��RIB+�_�_�a?���{�mi�Go5okoYo�o}l��P'rP�nܡݯ�o=_`�o�_�[R?�Q�u���  �p���o��/�� S��z
uүܠ�������ڱ�����������  /�M�w��e��������l2 wF�$��Gb���t��a�`�p�S�C��y�@p�5�G�Y�۠F�� Dz��� F�P D��]����پ��ʯܯ�� ��~�?��ͫ@@�?�K��K���K���
 �|�������Ŀֿ �����0�B�T�f�ܽ�V� ���{���1��$PARA�M_MENU ?�3�� � DEF�PULSEr�	�WAITTMOU�T��RCV�� �SHELL_�WRK.$CUR�_STYL���	�OPT��PT�B4�.�C�R_DECSN���e��� �ߣ����������� !�3�\�W�i�{����USE_PROG %��%�����CCR���e�����_HOST !F��!��:���T�`�V��/�X����_TIME��^���  ��GDEB�UG\�˴�GINP_FLMSK�����Tfp����PGA�  ����)CH�����TYPE���������� � -?hcu �������/ /@/;/M/_/�/�/�/ �/�/�/�/�/??%?�7?`?��WORD �?	=	RS�fu	PNSU�Ԝ2JOK�DRT�Ey�]TRACE�CTL 1x3���� �` &�`�`�>�6_DT Qy3�%@��0D �  #T�2@�8BU%6D&6D'6D(6DE)6D*6D`8B,6DU-6D.6D/6D06Dy16A�c�aB8@U��BR��HI��8BF�8B6D6D	�6D
6D6D6D�6D6D6D^�8B�6D6D6D6D�6D�8B6D6D�6D6DV�8Bj�8B�6D6DҀ8B�8B!6D"6D5OGOYOkO}OT�O�O�D�D�C �PM �R�O�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o������� ��#�5�G�Y�k�}� ������ŏ׈.A�Ev� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p���E r�����, >Pbt���� ���//(/:/L/ ^/p/�/�/�/�/�/�/ �/ ??$?6?H?Z?l? ~?�?�?�?�?�?�?�? O O2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�o �o�&8J\ n������� ��"�4�F�X�j�|� ������ď֏���� �0�B�T�f�x����� ����ҟ�����,� >�P�b�t��������� ί����(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l� ~ϐϢϴ����������� �*��$PGT�RACELEN � )�  ���(��>�_�UP z��e�m�u�Y�n��>�_CFG {Fm�W�(�~����PЬ� ��DEFS_PD |���a�P��>�IN��T_RL }��(��8��IPE_CO�NFI��~m�'�mњ��ԚҮ>�LID����~=�GRP 1���W��)�A ����&ff(�A+�33D�� D]�� CÀ A@1��Ѭ(�d�Ԭ���0�0�� 	 p1��1��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P;t _��������  Dz (�
 H�X~i�� ����/�/D/�//h/S/�/��
V�7.10beta�1��  A��E�"ӻ�Ay (�� ?!G��!/>���"����!����!BQ��!A\� �!���!2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?OO :O%O7OpO[O�OO�O �O�O�O�O_�O6_!_ Z_E_~_i_�_�_�_�_ �_�_'o2o�_VoAo So�owo�o�o�o�o�o �o.R=v1�<�/�#F@ �y�} ��{m��y=��1� '�O�a��?�?�?���� ��ߏʏ��'��K� 6�H���l�����ɟ�� �؟�#��G�2�k� V���z��������o ��ίC�.�g�R�d� ���������п	��� -�?�*�cώ���� �������B�;� f�x�������DϹ��� ���������7�"�[� F�X��|������� ����!�3��W�B�{� f��������� ��� ��/S>wbt ������ =OzόϾψ��� �ϼ� /.�'/R�d� v߈߁/0�/�/�/�/ �/�/�/#??G?2?k? V?h?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O���O�O�O_ _?_*_c_N_�_r_�_ �_�_�_�_o�_)oT fx�to���/ �o/>/P/b/t/ mo�|���� ���3��W�B�{� f�x�����Տ����� ��A�S�>�w�b��� �O��џ������+� �O�:�s�^������� ͯ���ܯ�@oRodo �o`��o�o�o��ƿ�o ���*<N�Y�� }�hϡό��ϰ����� ���
�C�.�g�Rߋ� v߈��߬�����	��� -��Q�c�N�ﲟ�� ��l��������;� &�_�J���n������� ����,�>�P�:L ����������� �(�:�3��0iT �x�����/ �///S/>/w/b/�/ �/�/�/�/�/�/?? =?(?a?s?��?�?X? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O*\&_8_r���_�_��$PL�ID_KNOW_�M  ��� Q�TSV ����P��?o"o4o�O�XoCoUo�o R�SM_GRP 1��Z�'0{`�@�`uf�e�`
�5� �g pk'Pe ]o�����������SMR�c�b�mT�EyQ}? yR ����������폯��� ӏ�G�!��-����� ������韫���ϟ� C���)���������`��寧���QST�a�1 1��)��v�P0� A 4� �E2�D�V�h������� ߿¿Կ���9��.� o�R�d�vψ��ϬϾϔ���2�0� Q�<3��3�/�A�S��4l�~ߐߢ��A5���������6
��.�@��7Y�k�}����8���������MAD  �)��PARNU/M  !�}o+���SCHE� S�
���f���S��UPD�f�x��_C�MP_�`H�� �'��UER_CHK-���ZE*�<RSr��_�Q_M�OG���_�X�__RES_G��!� ��D�>1bU �y�����/ �	/����+/ �k�H/g/l/��Ї/ �/�/�	��/�/�/� X�?$?)?���D?c?�h?����?�?�?�V� 1��U�ax�@c�]�@t@(@c�\�@�@D@c�[�*@��THR_INRr�J�b�U�d2FMASS?O �ZSGMN>OqCMO�N_QUEUE ���U�V P~P *X�N$ UhN�FV��@END�A��IEcXE�O�E��BE�@|�O�COPTIO�G���@PROGRAoM %�J%�@��?���BTASK_�IG�6^OCFG ���Oz��_�PDA�TA�c��[@Ц2=�DoVohozo�j 2o�o�o�o�o�o�);M jINFO
[��m��D�� ������1�C� U�g�y���������ӏ����	�dwpt�l �)�QE DIT ���_i��^WER�FLX	C�RGA�DJ �tZAЄ����?נʕFA��I�ORITY�GW�>��MPDSPNQ�����U�GD��OT�OE@1�X� _(!AF:@E� �c�Ч!tcp|n���!ud��>��!icm���?n<�XY_�Q�X�{��Q)� *�1�5��P��]�@� L���p��������ʿ ��+�=�$�a�Hυ�z��*��PORT)Q�H��P�E��_CARTREPP|X��SKSTA�H^�
SSAV�@�tZ�	2500H8�63���_x�
�'��*X�@�swPtS��ߕߧ���URGE��@B��x	WF��DO�F"[W\��������WRUP_DE?LAY �X��ԟR_HOTqX	B%��c���R_NOR�MALq^R��v�S�EMI�����9�Q�SKIP'��tUr�x 	7�1�1� �X�j�|�?�tU���� ����������$ J\n4���� ����4FX |j����� ��/0/B//R/x/�f/�/�/�/tU�$R�CVTM$��D��� DCR'����Ў!Bz8aB����C	0>?D���<?�7�{l2:��x�Ŝ�����ӷG���:�o?�� <
6�b<߈;܍��>u.�?!<�&�?h?�? �?�@>��?O O2ODO VOhOzO�O�O�O�O�O �?�O�O__@_+_=_ v_Y_�_�_�?�_�_�_ oo*o<oNo`oro�o �o�o�_�o�o�o�o �o8J-n��_� ������"�4� F�X�j�U������ď ���ӏ���B�T� �x���������ҟ� ����,�>�)�b�M� �����������ïկ �Y�:�L�^�p����� ����ʿܿ� ���� 6�!�Z�E�~ϐ�{ϴ� ������-�� �2�D� V�h�zߌߞ߰����� ����
���.��R�=� v��k�������� ��*�<�N�`�r��� ������������� &J\?���� �����"4�FXj|��!GN_ATC 1�	;� AT&�FV0E0��ATDP/6/9�/2/9�AT�A�,AT�%G1%B960��+++�,��H/,�!IO_TYPE  �%��#t�REFP�OS1 1�V+O x�u/�n �/j�/
=�/�/�/Q? <?u??�?4?�?X?�?��?�+2 1�V+ �/�?�?\O�?�O�?�!3 1�O*O<OvO��O�O_�OS4 1��O�O�O_�_t_�_>+_S5 1�B_T_�f_�_o	oBo�_S6 1��_�_�_5o�o��o�oUoS7 1� lo~o�o�oH3l�oS8 1�%�_���SMA�SK 1�V/  q
?�M��XNOS/��r������!MO�TE  n��$��_?CFG ����q����"PL_RAN�G�����POWE/R ������SM_DRYPR/G %o�%�P���TART ���^�UME_PR�O-�?����$_EX�EC_ENB  y���GSPD��pՐݘ��TDB���
�RM�
�MT_�'�T����OB�OT_NAME �o����OB�_ORD_NUM� ?�b!�H863  ��կ���P�C_TIMEOU�T�� x�S23�2Ă1�� L�TEACH ?PENDAN��wƋ�-��M�aintenance Cons�䃌s�"���KC�L/Cm��

����t�ҿ No Use-��Ϝ�0��NPO�򁋁���.�CH_Lf������q	��~s�MAVAIL������糅��SPA�CE1 2��, j�߂�D��s��߂� �{S�8�?�k�v�k�Z߬� �ߤ��ߚ� �2�D� ��hߊ�|��`����� ������ �2�D� ��h��|���`�����P����y���2��� �0�B���f�����@{���3 );M_�������/� /4 4FXj|*/�� �/�/�/?(??=?5Q/c/u/�/�/G?�/ �/�?O�?$OEO,OZO6n?�?�?�?�?dO �?�?_,_�OA_b_I_w_7�O�O�O�O�O �_�O_(oIoo^oofo�o8�_�_�_�_ �_�oo6oEf){���G �No� ���
M� ���*�<�N� `�r�������w���o �収���d.�� %�S�e�w��������� ��Ǐَ���Θ8�+� =�k�}�������ůׯ ͟����%�'�X�K� ]���������ӿ�������#�E�W� `� @����� ��x�����\�e��� ��������R�d߂� 8�j߬߾߈ߒߤ��� �������0�r��� X������������8����
�ύ�_MODE  �{^��S ��{|�2�0�����3��	S|)CWOR�K_AD��:���+R  �{��`� �� _INT�VAL���d���R_OPTION�� ��H VAT_GRP 2��uwp(N�k|��_ �����/0/B/ ��h�u/T� }/�/�/ �/�/�/�/?!?�/E? W?i?{?�?�?5?�?�? �?�?�?O/OAOOeO wO�O�O�O�OUO�O�O __�O=_O_a_s_5_ �_�_�_�_�_�_�_o 'o9o�_Iooo�o�oUo �o�o�o�o�o�o5 GYk-���u �����1�C�� g�y���M�����ӏ� ��	��-�?�Q�c��� �������������ǟ�;�M�_����$�SCAN_TIM��_%}�R ��(�#((�<}04d %d 
!D�ʣ��u�/�����+U��25���@�d5�P�g��]	���������dd��x�  P���w� ��  8� �ҿ�!���D�� $�M�_�qσϕϧϹπ�������ƿv��F�X��/� �;�ob��p�m��t�_D�iQ̡  � l�|�̡ĥ������ �!�3�E�W�i�{�� ������������� /�A�S�e�]�Ӈ��� ����������) ;M_q���� ���r���j� Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�%�/  0��6��!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O*�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo�O�OJ�o �o�o�o�o�o�o  2DVhz��������
�7?  ;�>�P�b�t����� ����Ǐُ����!� 3�E�W�i�{�������ß �ş3�ܟ� �&�8�J�\�n������������ɯ���;�,� �+��	123456{78�� 	� =5���f�x�������������
�� .�@�R�d�vψϚ�� ����������*�<� N�`�r߄߳Ϩߺ��� ������&�8�J�\� n�ߒ��������� ���"�4�F�u�j�|� �������������� 0_�Tfx�� �����I >Pbt���� ���!/(/:/L/ ^/p/�/�/�/�/�/�/�2�/?�#/9?�K?]?�iCz  �Bp˚   ��h2��*�$SC�R_GRP 1��(�U8(�\x�d�@� � ��'�	 �3�1�2�4(1*� &�I3�F1OOXO}m7��D�@�0�ʛ)���HUK�L�M-10iA 890?�90;��F;�?M61C D�:��CP��1
\&V �1	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^� oOUO>oPo#G�/血��o'o�o�o�o�oB�0�rtA9A�0*  @�BuD&Xw?��ju�bH0�{UzAF@ F�`�r��o��� ��+��O�:�s��m�Bqrr����������B�͏b����7�"�[� F�X���|�����ٟğ ���N���AO�0�B��CU
L���E�jqBq>gm󵔯$G@�@pnϯ B���G��I
E�0EL_DE�FAULT  ~�T��E���MIPOWE?RFL  
E*���7�WFDO�� *��1ERVENT 1���`�(�� L!DU�M_EIP��>���j!AF_IN�E�¿C�!FT$������!o:�� ��a�!RPC_MAINb��DȺPϭ�t�VIS�}�Cɻ����!TMP��PU�ϫ�d���E�!
PMON_�PROXYF߮�e 4ߑ��_ߧ�f�����!RDM_SR�V�߫�g��)�!�R�Iﰴh�u�!%
v�M�ߨ�id����!RLSYNC���>�8���!gROS��4��4�� Y�(�}���J�\����� ��������7��[ "4F�j|�� ��!�Eio��ICE_KL ?�%� (%S?VCPRG1n>���3��3���4//�5./3/�6V/[/�7~/�/�H�D�/�9�/�+� @��/��#?��K? ��s?� /�?�H/ �?�p/�?��/O� �/;O��/cO�?�O �9?�O�a?�O��? _��?+_��?S_� O{_�)O�_�QO�_ �yO�_��Os�� ��>o�o}1�o�o�o �o�o�o�o;M 8q\����� ����7�"�[�F� �j�������ُď�� �!��E�0�W�{�f� ����ß���ҟ�� �A�,�e�P���t���������ί�y_D�EV ���MC:��_]!�OUT���2��REC 1��`e�j� �� 	 ������ȿ���׿��!�
 ��PJ�%6 (޷&�!�a�}����,��0�  VZ� 3��3��Ge3�c���V��˒���  ���$��H�6�l�~� `ߢߐ��ߴ�������  ���V�D�z�h�� ������������
� �R�@�v���j����� ��������*N <^�r���� ��&J8Z �b������ �"/4//X/F/|/j/ �/�/�/�/��2��/�/ �/?:?(?^?L?�?�? v?�?�?�?�?�?�? O 6OOFOlOZO�O~O�O �O�O�O�O_�O2_ _ B_h_V_�_n_�_�_�_ �_�_
o�_.o@o"odo Rotovo�o�o�o�o�o �o<*`Np �x������ �8�J�,�n�\����� ����Ə�Ώ������F�4�j�X���`�p�V� 1�}� P��m���ܺ)I�� y!��TYPE\���HELL_CF�G �.�F��� � 	�����RSR������ӯ���� ���?�*�<�u�`�������������_�  ��!%Ϡ3�E��Q�\����M�o�p�����2���d]�K�:�HK ;1�H� u��� ����A�<�N�`߉� �ߖߨ������������&�8��=�OMM� �H���9�FT?OV_ENB&��!�1�OW_REG_�UI��8�IMWA�IT��a���OU�T������TIM������VAL|����_UNIT���K�1�MON_AL�IAS ?ew� ( he������ ������і��); M��q����d ��%�I[ m�<���� ��!/3/E/W//{/ �/�/�/�/n/�/�/? ?/?�/S?e?w?�?�? F?�?�?�?�?�?O+O =OOOaOO�O�O�O�O �OxO�O__'_9_�O ]_o_�_�_>_�_�_�_ �_�_�_#o5oGoYoko o�o�o�o�o�o�o�o 1C�ogy� �H����	�� -�?�Q�c�u� ����� ��ϏᏌ���)�;� �L�q�������R�˟ ݟ�����7�I�[� m��*�����ǯٯ� ���!�3�E��i�{� ������\�տ���� �ȿA�S�e�wω�4� �Ͽ����ώ����+� =�O���s߅ߗߩ߻� f�������'���K� ]�o���>������ ����#�5�G�Y���}���������o��$�SMON_DEF�PRO ������ �*SYSTEM*  d=���RECALL ?�}�� ( �}�/xcopy f�r:\*.* v�irt:\tmp�back7=>i�nspiron:?11828 Yb�t�� }0.a 6HZ_���4/s:orde�rfil.dat��Mbt�� }=+/mdb:�M Z��/�-�Q b/t/�/�/�</�a/��/??�!
xyz�rate 61 ��/�/�/n?�?�?�%|.7M(3304 H? Z?�?�?O�(3.@@�=aOsO�O�O� *��IO�4YO�O�O_�). ./A?�8�On_�_�_%. �/G_YR__�_oo'O 9O�O]_no�o�o�O�_ �O[o�o�o#_5_�_ Y_j|��_�_D�_ ���o1o�oUof� x����o�oJ��o��� ���-�Qb�t��� ���<������� )?��͟ߟp������?N'6368�?Y�� ���!�3�����a�s� ������E���Y���� �!�3�F�£ݿnπ� �ϥ�6�H�Š^���� �&�8���ܿm�ߑ� ����ȿZ������"� 4���X�i�{��ϲ� C���������0�����e�w�������U 2112ǯY����� !�3������n������400GY� �!�3߼߽as ����E�Y�� /!�3�F���n/�/ �/��6/H/� ^/�/? ?&8��m??�? ���Z?�?�?O"7��$SNPX_A�SG 1�����9A� �P 0 '%�R[1]@1.Y1O9?�$3%dO �OsO�O�O�O�O�O�O  __D_'_9_z_]_�_ �_�_�_�_�_
o�_o @o#odoGoYo�o}o�o �o�o�o�o�o*4 `C�gy��� ����	�J�-�T� ��c�������ڏ��� ��4��)�j�M�t� ����ğ������ݟ� 0��T�7�I���m��� �����ǯٯ���$� P�3�t�W�i������� �ÿ����:��D� p�Sϔ�wω��ϭ���  ���$���Z�=�d� ��sߴߗߩ�������  ��D�'�9�z�]�� ��������
���� @�#�d�G�Y���}��� ����������*4 `C�gy��� ���	J-T �c������ /�4//)/j/M/t/ �/�/�/�/�/�/�/?�0?4,DPARAM� �9ECA ��	��:P�4��0$HOFT_K�B_CFG  �q3?E�4PIN_S_IM  9K�6��?�?�?�0,@RVQSTP_DSB�>��21On8J0SR ���;� & �MULTIROB?OTTASK=Oq3��6TOP_O�N_ERR  ��F�8�APTN ��5�@A��BRING_PR�M�O J0VDT_GRP 1�Y9�@  	�7n8_ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2Dk hz������ �
�1�.�@�R�d�v� ��������Џ���� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\����������� ȯگ����"�I�F� X�j�|�������Ŀֿ ����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�tߛ� �ߪ߼��������� (�:�a�^�p���� �������� �'�$�6� H�Z�l�~���������������3VPRG_�COUNT�6�8�A�5ENB�O�M=�4J_UPD� 1��;8  
q2����� � )$6Hql ~�����/� / /I/D/V/h/�/�/ �/�/�/�/�/�/!?? .?@?i?d?v?�?�?�? �?�?�?�?OOAO<O NO`O�O�O�O�O�O�O �O�O__&_8_a_\_�n_�_�_�_YSDOEBUG" � �P�dk	�PSP_PA�SS"B?�[L�OG ���m�P�X�_  ��g�Q
MC:�\d�_b_MPC m��o�o�Qa�o� �vfSAV žm:dUb�U�\gSV�\TEM_TIME 1��� (�`"�S ��o	T1SVGU�NS} #'k��spASK_OPT�ION" �go�spBCCFG ��| �b�{�}`����a&�� #�\�G���k�����ȏ ������"��F�1� j�U���y���ğ��� ӟ���0��T�f��UR���S���ƯA��� ��� ��D��nd��t 9�l���������ڿȿ �����"�X�F�|� jϠώ��ϲ������� ��B�0�f�T�v�x� ���ߦؑ������� (��L�:�\��p�� ���������� �6� $�F�H�Z���~����� ��������2 V Dzh����� ����4Fdv ������/ /*/�N/</r/`/�/ �/�/�/�/�/�/?? 8?&?\?J?l?�?�?�? �?�?�?�?�?OO"O XOFO|O2�O�O�O�O �OfO_�O_B_0_f_ x_�_X_�_�_�_�_�_ �_oooPo>otobo �o�o�o�o�o�o�o :(^Lnp� ����O��$�6� H��l�Z�|�����Ə ؏ꏸ����2� �V� D�f�h�z�����ԟ ����
�,�R�@�v� d���������ίЯ� ��<��T�f����� ��&�̿��ܿ��&� 8�J��n�\ϒπ϶� �����������4�"� X�F�|�jߌ߲ߠ��� ��������.�0�B� x�f��R��������� ���,��<�b�P��� ����x��������� &(:p^�� ����� 6 $ZH~l��� �����/&/D/V/ h/��/z/�/�/�/�/��&0�$TBCS�G_GRP 2���%� � �1 
 ?�  /?A?+?e?O? �?s?�?�?�?�?�;2�3�<d, ��$A?1	 HC{���6>��@E~�5CL  B�'2�^OjH4J��B�\)LFY  A��jO�MB��?�IBl��O�O�@�JG_�@�  D	�15_ __�$YC-P{_F_`_j\��_�]@0�>�X�Uo �_�_6oSoo0o~o�o��k�h�0	V�3.00'2	mw61c�c	*�`0�d2�o�e>�JC0(�a�i ,p�m-w  �0����o�mvu1JCFG [��% 1 #0vz��rBr�|�|����z� � %��I�4�m�X���|� �������֏���3� �W�B�g���x����� ՟��������S� >�w�b�����'2A �� ʯܯ������E�0� i�T���x���ÿտ� �����/��?�e�1 �/���/�ϜϮ����� ���,��P�>�`߆� tߪߘ��߼������ ��L�:�p�^��� ���������� �6� H�>/`�r�������� �������� 0V hz8����� �
.�R@v d������� //</*/L/r/`/�/ �/�/�/�/�/�/�/? 8?&?\?J?�?n?�?�? �?�?���?OO�?FO 4OVOXOjO�O�O�O�O �O�O__�OB_0_f_ T_v_�_�_�_z_�_�_ �_oo>o,oboPoro to�o�o�o�o�o�o (8^L�p� ������$�� H�6�l�~�(O����f� d��؏���2� �B� D�V�������n���� ԟ
���.�@�R�d�� ��v��������Я� ��*��N�<�^�`�r� ����̿���޿�� $�J�8�n�\ϒπ϶� ��������ߊ�(�:� L���|�jߌ߲ߠ��� �������0�B�T�� x�f���������� ����,��P�>�t�b� �������������� :(JL^�� ���� �6 $ZH~l��^� ��dߚ //D/2/ h/V/x/�/�/�/�/�/ �/�/?
?@?.?d?v? �?�?T?�?�?�?�?�? OO<O*O`ONO�OrO �O�O�O�O�O_�O&_ _6_8_J_�_n_�_�_ �_�_�_�_�_"ooFo ��po�o,oZo�o�o �o�o�o0Tf x�H����� ��,�>��b�P��� t���������Ώ�� (��L�:�p�^����� ��ʟ���ܟ� �"� $�6�l�Z���~����� دꯔo��&�ЯV� D�z�h�������Կ¿ ��
��.��R�@�v�8dϚτ�  ����� �������$�TBJOP_GR�P 2ǌ���  ?�������������xJ�BЌ��9� �<� �X����� @���	 ��C�� t�b  �C����>��1͘Րդ�>̚й���33=�C�Lj�fff?��?�ffBG��ь������t�ц�>��(�\)�ߖ�E����;��hCY�j��  @h��B�  A����f�~��C�  Dh�8��1��O�4�N�����
:���Bl^��j�i�l�l�����Aə�A��"��D��֊=qqH���нp�h���Q�;�A}�j�ٙ�@L��D	2�������$�6�>B�\��T���Q��tsx�@33@���C���y�x1����>��Dh�����������<{�h�@i�  ��t��	��� K&�j�n| ���p�/�/(:/k/�ԇ���!��	V3.00J��m61cI�*� IԿ��/�' �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I��!CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;��;Q�T,8�4` *�ϴ?�2���3\�X/O���ESTPARS c ��	���HR@ABLE 1���I�0��
H�7 8��9
G
H
H����*
G	
H

H
HYE���
H
H
HN6FRDIAO�XO@jO|O�O�O�ETO"_�4[>_P_b_t_�^:BS _� �JGoYoko}o �o�o�o�o�o�o�o 1CUgy�� ��`#oRL�y�_�_�_ �_�O�O�O�O�OX:B~�rNUM  �ū�P��� �V@P:B_CFG �˭�Z�h�@��IMEBF_TT%ApU��2@�VERS��q��R 1̞��
 (�/����b� ����J�\��� j�|���ǟ��ȟ֟� ����0�B�T���x��������2�_���@��
��MI_CH�AN�� � ��DOBGLV����������ETHERA�D ?��O��������h�����R�OUT�!��!�������SNMA�SKD��U�25�5.���#�����O�OLOFS_DI�%@�u.�ORQC?TRL ����� }ϛ3rϧϹ������� ��%�7�I�[�:����h�z߯�APE_D�ETAI"�G�PON_SVOFF=����P_MON ��֍�2��STRTCHK �^������VTCOM�PAT��O�����FPROG %^��%MULTIROBOTTݱ��֞9�PLAY&H��_�INST_Mް 2������US�q�΃�LCK���QUICKME�=���oSCREZ�G�tps� ���u�z����_��@@n��.�SR_GRP �1�^� �O����
��+O=sa�쀚�
 m������L/ C1gU�y� ����	/�-//�Q/?/a/�/	1234567�0�/�/�@Xt�1���
 ��}ipnl/�� gen.htm��? ?2?D?V?`�Panel s/etupZ<}P�?`�?�?�?�?�? �? ?,O>OPObOtO�O�? �O!O�O�O�O__(_ �O�O^_p_�_�_�_�_ /_]_S_ oo$o6oHo Zo�_~o�_�o�o�o�o �o�oso�o2DVh z�1'��� 
��.��R��v����������ЏG���UA�LRM��G ?9� �1�#�5�f� Y���}�������џן����,��P��SEoV  �����ECFG ���롽�A��  w BȽ�
 Q� ��^����	��-�?� Q�c�u������������� �����eI��?���(%D� 6� �$�]�Hρ�lϥ� ���ϴ�������#��G���� �߿U��I_Y�HIST �1��  (��� ��3/S�OFTPART/�GENLINK?�current=�editpage,��,1���!�3�ν�� ����me;nu��962�߆������K�]�o�36 u�
��.�@���W�i� {���������R����� /A��ew� ���N�� +=O�s��������f��f/ /'/9/K/]/`�/�/ �/�/�/�/j/�/?#? 5?G?Y?�/�/�?�?�? �?�?�?x?OO1OCO UOgO�?�O�O�O�O�O �OtO�O_-_?_Q_c_ u__�_�_�_�_�_�_ ��)o;oMo_oqo�o �_�o�o�o�o�o�o %7I[m�  �������3� E�W�i�{������Ï Տ�������A�S� e�w�����*���џ� ����ooO�a�s� ��������ͯ߯�� �'���K�]�o����� ����F�ۿ����#� 5�ĿY�k�}Ϗϡϳ� B���������1�C� ��g�yߋߝ߯���P� ����	��-�?�*�<� u����������� ��)�;�M������ ����������l� %7I[���� ���hz!3 EWi����� ��v////A/S/�e/P���$UI_�PANEDATA 1�����!�  	�}w/�/�/�/�/?? )?>?��/i? {?�?�?�?�?*?�?�? OOOAO(OeOLO�O �O�O�O�O�O�O�O_.&Y� b�>RQ? V_h_z_�_�_�__�_ G?�_
oo.o@oRodo �_�ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_ ��!�3�E�W��{� �_����ÏՏ���`� �/��S�:�w���p� ����џ������+� �O�a��������� ͯ߯�D����9�K� ]�o��������ɿ�� �Կ�#�
�G�.�k� }�dϡψ����Ͼ��� n���1�C�U�g�yߋ� �ϯ���4�����	�� -�?��c�J���� ������������;� M�4�q�X������� ����%7��[ �������@ ��3WiP �t�����/ �//A/����w/�/�/ �/�/�/$/�/h?+? =?O?a?s?�?�/�?�? �?�?�?O�?'OOKO ]ODO�OhO�O�O�O�O N/`/_#_5_G_Y_k_ �O�_�_?�_�_�_�_ oo�_Co*ogoyo`o �o�o�o�o�o�o�o�-Q8u�O�O}��������)�>��U-�j�|��� ����ď+��Ϗ�� �B�)�f�M������� �������ݟ�&�S��K�$UI_PA�NELINK 1��U  ��  ���}1234567890s��������� ͯդ�Rq����!�3� E�W��{�������ÿ�տm�m�&����Qo�  �0�B�T�f� x��v�&ϲ������� ��ߤ�0�B�T�f�x� ��"ߘ���������� �߲�>�P�b�t��� 0������������ $�L�^�p�����,�>�������� $�0,&�[gI�m� ������> P3t�i��� �� -n��'/9/K/ ]/o/�/t�/�/�/�/ �/�/?�/)?;?M?_? q?�?�UQ�=�2"� �?�?�?OO%O7O�� OOaOsO�O�O�O�OJO �O�O__'_9_�O]_ o_�_�_�_�_F_�_�_ �_o#o5oGo�_ko}o �o�o�o�oTo�o�o 1C�ogy�� ���B�	��-� �Q�c�F�����|��� ����֏�)��M� ��=�?��?/ȟڟ ����"�?F�X�j� |�����/�į֯��� ��0��?�?�?x��� ������ҿY���� ,�>�P�b��ϘϪ� ������o���(�:� L�^��ςߔߦ߸��� ����}��$�6�H�Z� l��ߐ��������� y�� �2�D�V�h�z� ���-���������
 ��.RdG�� }����c��� <��`r���� ����//&/8/J/ �n/�/�/�/�/�/7� I�[�	�"?4?F?X?j? |?��?�?�?�?�?�? �?O0OBOTOfOxO�O O�O�O�O�O�O_�O ,_>_P_b_t_�__�_ �_�_�_�_oo�_:o Lo^opo�o�o#o�o�o �o�o ��6H� l~a����� ���2��V�h�K� ������1�U
� �.�@�R�d�W/���� ����П������*� <�N�`�r��/�/?�� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��+������:� L�/�p���e������� ���� ��6����ۏ��$UI_�QUICKMEN�  ����}��REST�ORE 1٩��  �A
�8m3 \n���G�� ��/�4/F/X/j/ |/'�/�/�//�/�/ ??0?�/T?f?x?�? �?�?Q?�?�?�?OO �/'O9OKO�?�O�O�O �O�OqO�O__(_:_ �O^_p_�_�_�_QO[_ �_�_I_�_$o6oHoZo loo�o�o�o�o�o{o �o 2D�_Qc u�o������ �.�@�R�d�v����ଏ��Џ⏜SCR�E� ?��u1sc� u2��3�4�5�6��7�8��US#ER����T���Sks'���4��5���6��7��8��� N�DO_CFG mڱ  �  � PDATE h���None��SEUFRAM/E  ϖ���RTOL_ABRqT����ENB(�~�GRP 1��	��Cz  A� ~�|�%|�������įB֦��X�� UH��X�7�MSK  hK�S�7�N�%u�T�%�����VIS�CAND_MAX�I�I�3���FA?IL_IMGI�z ��% #S���IMR_EGNUMI�
����SIZI�� ��ϔ,�ONTM�OU'�K�Ε��&����a��a���s�FR�:\�� � �MC:\(�\L�OGh�B@Ԕ �!{��Ϡ�����z MCV�����UD1 �EX�	�z ��PO6�4_�Q��nm6��PO!�LI��Oڞ�e�V�N�fy@`�I�� =	_�wSZVmޘ��`��WAImߠ�STAOT �k�% @��4�F�T�$#�x ��2DWP  ���P G��=���͎���_J�MPERR 1��
  �p2345678901�� ��	�:�-�?�]�c� ��������������<��$�MLOW�ޘ������_TI/�˘'���MPHASE'  k�ԓ� ���SHIFT%�1 Ǚ��<z�� _����F /|Se���� ���0///?/x/ O/a/�/�/�/�/�/�����k�	VSF�T1\�	V��MN+3 �5�Ք p�����A�  B8*[0[0�Πpg3a1bY2�_3Y�7ME���K�͗	6e���&%���M���b���	��$��TDINGEND3�4��4OH�+�G1�OS2OIV �I���]LREL�EvI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�Y?BOX �ǝf_V\��b�2�TI�190.0.��P83p\�V2�54p^�Ԓ	 ��S�_�[b��?robot84q_   p�<9o\�pc�PZo Mh�]Hm�_Jk@1�o�ZABCd��k�, ���P\�Xo}�o0 );M�q���������>��aZ�b��_V