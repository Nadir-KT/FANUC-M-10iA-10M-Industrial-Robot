��   �A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���F�SAC_LST_�T   8 �$CLNT_NA�ME !$I�P_ADDRES}SB $ACCN �_LVL  �$APPP   � �$8 AO  O���z�����o VIRTUAqLw�'DEF\ �� � �����ENABL�E� �����L?IST 1 ��?  @!������
[. @�d����� /�3//W/*/</�/ `/�/�/�/�/�/�/�/ ??S?&?8?J?�?n? �?�?�?�?�?O�?�? OO"OsOFO�OjO|O�O �O�O�O_�O�O7__ \_B_�_f_x_�_�_�_ �W