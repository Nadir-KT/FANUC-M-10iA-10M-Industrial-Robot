��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ���(�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1��'|U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|  �ARG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"�SB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5�UTOB�ACKU0 $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�:�OFF_ N�3D;ELHLOGn25Aa2?i1@N�?�� -M��W�+0�$Y $DB\� 6COMW!2�MO� 21\D.	� \rVE�1$qF��A{$O���D�B�CTMP1_5F�E2�G1_�3�B��2	�XD�#�
 d $CA�RD_EXIST�4$FSSB_�TYPuAHKBgD_S�B�1AGN �Gn $SL?OT_NUMJQoPREV,DBU� �g1�;1_EDIT�1 � 1G�=� S�0%$�EP�$OP��AETE_�OKRUS�P_CRQ$;4�V� ^0LACIw1`�RAPk �1x@ME@$D�V�Q�P�v�A{oQL� OUzR ,mA�0��!� B� LM_O��^eR�"CAM_�;1 xr$ATTR4NP� �ANN�@5IMG?_HEIGHQ�c�WIDTH4VT�� �UU0F_ASwPECQ$M�0gEXP��@AX�f��CFT X O$GR� � S�!z�@B@NFLI�`<t� UIRE 3dT�uGITCHC�`N�� S�d_L�`�C��"�`EDlpE� J�4S�0� �zsa�!ip�;G0 � 
?$WARNM�0f�!,P� �s�pNST�� CORN�"a1F�LTR�uTRAT�� T�p H0AC�Ca1���{�OcRI
`"S={RT0�_S�BMO�CHuG,I1 [ �Tp�"3I9�TYP�D,P*2 �`w@�� �!R*HD�cJ�* C��2��3��4���5��6��7��8���94�qO�$ <� $6xK3 1�w`O_M�@�C �t � E#6NGP�ABA� �c��@ZQ���`���@nr��� ��P�0����x�p�PzPb26h����"J�_R���BC�J��3�JVP��tBS��}Aw���"�tP_*0OFS�zR @� RO_�K8���aIT�3��N'OM_�0�1ĥ384 ��T �� $�d��AxP��K}EX��� �0g0I01��p�
�$TFa��C$MDM3��TO�3�0U� ^�� �Hw2J�C1|�EΡg0wE�{vF�vF�40CPhp@�a2 
P$A`�PU�3N)#�dR*�AX�!sDEwTAI�3BUFV8��p@1 |�p۶��pPIdT� PP�[�MZ�Mg�Ͱj�F>[�SIMQSI�"�0��A.����kx 	Tp|zM��P�B��FACTrbHPE�W7�P1Ӡ��v��M]Cd� �$*1�JB�p<�*1DEC�Hښ�H��(�c� �� +PNS_E;MP��$GP���B,P_��3�p�@Pܤ��TC��|r��0�s ��b�0�� �B���!
����JR� ��SEGKFR��Iv �aR��TkpN&S,�PVF�4��� & k�Bv�u�cu��aE�� �!2��+�MQ��E�SI!Z�3����T��P������aRSINF �����kq���������LX�����F�C3RCMu�3CClpG� �p���O}���b�1��������2�V�DxIC��C���r����P��L{� EV �zF�_��F�pNB0��?������A�! �r�Rx����V�lp �2��aR�t�,�g��}RTx #� 5�5"2��uAR���`�CX�$LG�p��B@�1 `s�P�t�aA�0�{�У+0R���tM�E�`!BupCrRA 3tAZ�л�pc��OT�FC�b�`�`F�Np���1��ADI +�a%��b�{��p $�pSp�c�`S�P�L�a,QMP6�`Y�3z��M'�CU���aU  $>�TITO1�S�S�!���$�"0�DBPXW�O��!��$SiK��2�@DB��"�"@�PR8�� 
� ���# �>�q1$��$��+�L9$?(�V�R%@?R4C&_?�R4ENE��'�~?(�� RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@4a��C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!� C{S_)  `IS#� �� �s3S�AQ汯 4Rx�ZS W�AQ�p�@1UW��cT'NTV)�5RV
a�@��|c�éWƃ��JBx��x0��SAFEۥ��V_SV�bEXC�LUU�;��ON�L��cYg�~az�OyT�a{�HI_V? ���R, M�_ *Ȥ0� ��_z�2� ��QSGO  +�rƐm@�A�c~b����w@��V�i�b�fA�NNUNx0�$�dI%DY�UABc�@Sp��i�a+ �j�f�"�pO�GIx2,��$F��b�$ѐOT�@A� $DUMMY ��Ft��Ft±� 6�U- ` !�HE�|s��~bc�B@ �SUFFI��V4PCA�Gs5Cw�6dr�!MSWU.{ 8��KEYI��5�TM�1�s�qoA�v�INޱE��!, /{ D��HOST�P!4���<���<�°<��p<�EM'���Z�n� SBL� UL��0  �	�����DT�01 ϴ $��9USAMPLо�/����ĺ�$ I@갯 $SUBӄ��w0QS��8���#��SAV������c�S< 9�`�fP�$�0E!� YN_�B�#2 0��DI��d�pO|�m��#$�F�R_IC� �?ENC2_Sd�3  ��< 3�9����� cgp����4��"��2�A��ޖ5���`ǻ�@Q@�K&D-!�a�AVE�R�q����DSP
���PC_�q��"�x|�ܣ�VALU3��HE�(�M�IP\)���OPPm �CTH�*��S" $T�/�Fb�;�d�����d D�qЗ16� H(rLL_DU ǀ�a�@��k���֠OT�"U�/���@@�NOAUTO7�0�$}�x�~�@sT��|�C��C� �2v�L�� 8/H *��L� � ��Բ@sv��`� �� � ����Xq��cq���q��T�q��7��8��9���0���1�1 �1�-�1:�1G�1T�1*a�1n�2|�2��U2 �2-�2:�2G�U2T�2a�2n�3|ʥ3�3� �3-�3�:�3G�3T�3a�3zn�4|��'�����9 <���z�ΓKI����H硵Ba�FEq@{@: ,<��&a? P_P�?��>�����E@�@���!QQ��;fp�$TP�$V�ARI����,�UP�2Q`< W�߃TD ��g���`���������BAC�"= T2����$)�,+r³�p IFI��p�� q M�P"�l@``>t ;��6����ST����T ��M ����0	��i� ��F���������kRt �����FORCEUyP�b܂FLUS
p�H(N��� ��6bD_CM�@E�7N�� (�v�P��REM� Fa��@j����
K�	N���EcFF/���@IN�Q�OV��OVA��	TROV DyT)��DTMX: e �P:/��Pq�XvXpCLN _�p���@ ��	_|��_QT: �|�&PA�Q	DI���1���0�Y0RQm�_�+qH���M���CL�d#�RIV{�ϓN"�EAR/�IO�P�CP��BR��C�M�@N 1b 3GgCLF��!DY�(ء�a�#5T�DG����� �%iaFSS� )�? P(q1�1��`_1"811R�EC13D;5D6O�GRA���@��i���PW�ON2EBUG�S�2��C`gϐ_E A� ��o��TE�RM�5B�5���O�RIw�0C�5���GSM_-`���0D�5�L��TA�9E�IUP��F� -QϒA�P�3�@�B$SEGGJ� E�L�UUSEPNFI��pBx��1@��4�>DC$UF�P��C$���Q�@C��ĳG�0T�����SNSTj�PATۡg��AOPTHJq�A�E*� Z%qB\`F�{E��F�q��pARxPY�aSHF�T͢qA�AX_SH�OR$�>��6 @$�GqPE���OVRH���aZPI@P@$U?r= *aAYLO���j�I�"��Aؠ��ؠERV��Qi�[Y)� �G�@R��i�e��i��R�!P�uASYM���uqAWJ�G)��AE��Q7i�RD�U[d@�@i�U��C�%UP��X�P���WOR�@M��u�GRSMT��GƇ�GR��3�aPA�@��p5�'�H �� j�A�TOC�jA7pP]Pp$O�Pd�O��C�%�p��O!��RE.pRĈC�AO�?��Be�5pR�EruIx'QG�eo$PWR) IMdu��RR_$s��5��B �Iz2H8�=�_A�DDRH�H_LE�NG�B�q�q:�x�Rj��So�J.�SS��SK������ ��F-�SE*���rSN�[MN1K	�j�05�@r�֣OL��\��WpW�Q�>pACRO �p���@H ����Q�� ��OUPW3�b_">�I��!q�a1���� ����|���������-���:���iIO
X2S=�D�e��]���L $��p�!�_OFF[r_�PR�M_�v�HTT�P_�H��M (��pOBJ�"�pG�-$H�LE�C��ٰ�N � 9�*�AKB_�T��
�S�`l�S��LV��KRW"~duHITCOU?[BGi�LO�q�����d� Fpk�GpS9S� ���HWh�wA��O.��`INC�PUX2VISIO ��!��¢.�á<�á~-� �IOLN)�P 87�R'�[p�$SL�bd PU�T_��$dp�P�z �� F_AS:2Q/�$LD����D�aQT U�0]P�A0���0��PHYG灱�Z���5�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp���hx��ٶr�UJ���S����NE�WJO9G�G �DIS��r�1KĠ��3T |��AqV��`_�CTR!S�^�FLAGf2r�LG�dU �n�:��~�3LG_SIZ���ň��=���FD��I����Z �ǳ��0 �Ʋ�@s��-ֈ�-�=��-���-��0-�ISC#H_��Dq��N?���V��EE!2�C�D��n�U�����`L��n��DAU��EA��0Ġt����GHr��I�BOO)�WL3 ?`�� ITV����0\�REC�SCRf 0�a�D^�����MARG��`!P�)� T�/ty�?I�S�H��WW�I���T�JGM���MNCH��I�F�NKEY��K��PRG��UF��P��FWD��HL�STP��V��@�����RSS�H�` �Q�C�T1�ZbT�R ���U�����|R��t�i�2��G��8PPO��6��F�1�M��FOCU���RGEXP�TU%I��IЈ�c�� n��n����ePf����!p6�eP7�N���CA�NAI�jB��VAI�L��CLt!;eDCS_HI�4�.��O�|!�S �Sn�'��_�BUFF1XY��PT�$�� �vP��fĘ�1�A�rYY���P �����pOS1�2�3���>0Z �  ��apiE�*��IDX�d	P�RhrO�+��A&+ST��R��Yz�<!� Y$EK&C K+���Z&m&z��5�0[ L��o�0�� ]PL�6pwq�t^����w���7�_ \ �����瀰�7��#�0C��] ��CLD�P��;eTRQLI��jd.�094FLG z�0r1R3�DM�R7Ɩ�LDR5<4R5ORG.���e2(`���V�8�.��T<�4�d^ ��q�<4��-4R5S�`T�00m��0DFRCLMC!D�?�?3I@���MIC��d_ d����RQm�q�DgSTB	�  �Flg�HAX;b �H>�LEXCESZr��RrBMup�a`��B�;doE`��`a��F_A�J��$[�O�H:0K�db \��ӂnS�$MB��LIБ~}SREQUIR�R�>q�\Á�XDEBUT��oAL� MP�c�b�a��P؃ӂ!BoAND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@qt��o��UPST8�w e�rLOC��RI�p�EX�fA��p��AoAODAQnP�f X��ON��[rMF�����f)�"�I��%�e��T�$��FX�@IGG� g �q��"E�0�h�#���$R�a%;#�7y��Gx��VvCPi�D'ATAw�pE:�y���RFЭ�NVh t_ $MD�qIёA)�v+�tń�tH�`��P�u�|��sANSAW}��t�?�uD��)�b�	@Ði �@CU��V�T0�ewRR2�j Dɐ��Qނ�Bd$CALII�@F�G�s�2⠧RIN��v�<��NTE���kE���,�X�b����_Nl���ڂ��kDׄRm�DIViFDH�@ـn�$V��'c!;$��$Z������~�[��o�H �$BELT|b��!ACCEL+q��ҡ��IRC��t����T/!��$SPS�@#2L�@qЀƔ83������� ��P�ATH��������3̒Vp�A_�Q�.�4��B�Cᐈ�_MGh�$DDQ���G�$FWh��p��m�؝���b�DE��PP�ABNԗROTS�PEED����00J��Я8��@���@$OUSE_��P��Fs�SY��c�A kq�YNu@Ag��OF�F�q�MOUN�N�Gg�K�OL�H�INC*��a��q��Bj�<L@�BENCS��q`�Bđ���D��IN#"�I̒��4�\BݠVE�O�w�Ͳ23_UP�E�߳LOWL ���00����D���B wP��� �1RCʀƶ�MOSIV�JRMO����@GPERCH  �OV��^� �i�<!�ZD<!�c�� d@�P��V1�#P͑��L���EW��ĸ�UP������TR�Kr�"AYLOA 'a�� Q-�̒<�1Ӣ`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H����b��DUM2(�S_BCKLSH_C̒ ��>�=�q�#�U��ԑ����2�t�]ACLAL�vŲ�1n�P�CH�K00'%SD�RTY@4�k��y�1�q_6#N2�_UM$Pj�Cw��_�SCL��ƠLM?T_J1_LO��@���q��E�����p�๕�幘SPC��07������PCo���!H� �PU�m�C/@�"sXT_�c�CN_��1N��e���SFu���V�&#����9�̒��2=�C�u�SH6#�� c����1�Ѩ�o�0�͑�
��_�PAt�h�_	Ps�W�_10��4�R�P01D�VG�J� L�@�J�OGW���TO7RQU��ON*�M����sRHљ��_W��-�_=��C��I���I�I�II�F��`�JLA.�1[�VEC��0�D�BO1Up�@i�B\JRKU���	@DBL_S�Md�BM%`_DLC�BGRV��C��I��H_� ��*COS+\�(LN�7+X>$C�9)I�@9)u*c,)�Z2 �HƺMY@!�( "T�H&-�)THET0�NK23I��"=��A CB6CB=�C �A�B(261C�616�SBC�T25GTS QơC��aS$" ��4c#�7r#$DU D�EX�1s�t��B�6��r�AQ|r�f$NE�D�pIB U�\B5��$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2�&P�C�J�&!�VAHV6HT3�YLVhJVuKV�KUV�KV�KV�KV�IHAHZF`RXM��wXuKUH�KH�KH�KH�KUH�IO2LOAHO�Y�WNOhJOuKO�KO��KO�KO�KO�&F��2#1ic%�d4GSP�BALANCE_l�!�cLEk0H_�%SP��T&�bc&�br&PFULC�hr�g�rr%Ċ1ky�UT�O_?�jT1T2Cy��2N&�v�ϰct�w�g�p�0Ӓ~���T���O���� INSsEGv�!�REV�v�!���DIF��1�l�w�1m
�OB0�q
����MIϰ1�~�LCHWAR��波AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|���7ROBR�CR��zN���MSK_�`�f�p P Np_���R����΄ݡ�1 ��ҰТ΀ϳ��΀"��IN�q�MTC�OM_C@j�q � L��p��$ONORE³5����$�r 8� GRl�E�SD�0ABF��$XYZ_DAx5A���DEBU�qXI��Q�s �`$�wCOD�� ���k�F�f�$BU_FINDXР��MOR��t $-�U��)��r�B���������Gؒu �� $SIMU�LT ��~�� ���O�BJE�` �ADJ�US>�1�AY_I�k��D_����C�_[FIF�=�T�  ��Ұ��{��p� ������p�@��D�FRI4��ӥT��RO� ���E�����OPW�O�ŀv0��S�YSBU�@ʐ$SCOP����#�U"���pPRUN�I�P�A�DH�D����_�OU�=��qn��$}�IMAG��4ˀ�0P�qIM�����IN�q���RGO�VRDȡ:���|�P0~���Р�0L_6p���i��RB���02��M���EDѐF� ��N`M*��ඁ�˱SL�`ŀw x $OVSL�vwSDI��DEXm�@g�e�9w�����V� ~�N���w����Û�4�ȳ�M����q|<��� x Hˁ�E�F�ATUS����C�0àǒ��BT�M����If���4p����(�ŀy Dˀ!Ez�g���PE�r��p���
���EXE���V��E�Y�$Ժ ŀz3 @ˁ��UP{�h�3$�p��XN����9�H� �PG�"�{ h $S#UB��c�@_��01�\�MPWAI��PL����LO��-�F�p��$RCVFA�IL_C�-�BW�D"�F���DEFS}Pup | Lˀ�`�D�� U�UN!I��S���R`���_L�pP��̐���ā}��� B�~����|��`ҲN�`KET���y���P� $�~z���0SIZE��ଠ{���S<�OR~��FORMAT/p` � F���rEMR��y�UX����LI7�ā  �$�P_SWI|���AX_PL7�?AL_ �ސR�A��B�(0C��Dnf�$Eh�����C_=�U� �� � ���~�J�3�0����TIA4���5��6��MOM������� �B�AD��*��* PU70NRW���W R����� A$PI�6���	 ��)�4l�}6�9��Q���c�SPEED�PGq�7�D� >D����>tMpt[��SAM�`�痰>��MOV ���$��p�5��5�D�1�$2��������{�Hip�IN?,{�F(b+=$��H*�(_$�+�+GAM�M�f�1{�$GE�T��ĐH�D����
�^pLIBR�ѝI.��$HI��_��Ȑ$*B6E��*8A$>G086LW=e6\<G9�6�86��R��ٰV��$PDCK�DQ�H�_����;" ��z�.%�7�4*�9�� �$IM_SRO�D�s"���LH�"�LE�O�0\H��6@�R� �ŀ��P�qUR_S�CR�ӚAZ��S_?SAVE_D�E��NO��CgA�Ҷ� �@�$����I��	�I � %Z[� ��RX"  ��m���"�q�'" �8�Hӱt�W�U�pS�����U�M�� O㵐.'}q��Cg�� �@ʣ����S�M�AÂ�� � $PY���$WH`'�NGp���H`��Fb��Fb��Fb��PLM���	�P 0h�H�{�X��O���z�Z�eT�M���� pS��C��O_�_0_B_�a��_%�� |S����@	�v��v �@���w�v��E�M��%O�fr�B�ːt��ftP��PM���QU� �U�Q���A-�QTH=�H{OL��QHYS�3ES�,�UE��B���O#��  -�P�0�|�gAQ���ʠu���O��ŀ�ɂv�-�8�A;ӝROG��a2D�E�Âv�_�Ā^Z�INFO&��+�h���bȜ�OI��� ((@SLEQ /�#������o���S`c0O�0�051EZ0NUe�_��AUT�Ab�COPAY��Ѓ�{��@M���N�����1�P�
� ���RGI�����X_�Pl�$�����`
�W��P��j@�G����EXT_CY�Ctb���p�����h�_NA�!�$�\�<�RO�`]��� � m��P�OR�ㅣ���SReVt�)����DI �T_l���Ѥ{�ۧ�Шۧ �ۧ5٩6٩7�٩8��'�PS��B쐒��$�F6���PL�A�A^�TAR��@E `�Z�����<��d� ,�(@FLq`h��@YN�L���M�C���P�WRЍ�쐔e�D�ELAѰ�Y�pA�D#q�RQSKIPN�� ĕ�x�O�`�NT!� ��P_ x���ǚ@�b�p1� 1�1Ǹ�?� �?���>��>�&�>�3�>�9��J2R;쐖� 4��EX� TQ ����ށ�Q���[�K�Fд�8�RDCIf�S �U`�X}�R��#%M!*�0�)��$RGoEAR_0IO�T�JBFLG�igpE	Ra��TC݃�����ӟ2TH2N��� �1�b��Gq TN�0 ����M����`Ib��w�REuF�1�� l�h���ENAB��lcTPE?@���!(ᭀ ����Q�#�~�+2 (H�W���2�Қ���"�4�F�X�j�3�қ�{��������j�4�Ҝ��
��.�@�R�W ��5�ҝu�@����������j�6�����(:L��7�ҟo����(��P��8�Ҡ���"4Fj�SMS�K�����a��E��A��MOTE������@ "1��Q�IO�5"%I��P���Rd�Wi@쐣 � �����X�gpi�쐤���Y"$DSB_S�IGN4A�Qi�̰C|���tRS232%��Sb�iDEVIC�EUS#�R�RPA�RIT�!OPB�IT�Q��OWCONTR��Qⱓ֧RCU� M�SUX/TASK�3NB��0��$TATU�P%��S@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�UKPDl�ARB�#P%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG �G|�.2���F��1�!d�9Z�8+5K��+5��E�y�L0�4��X �0m�LN�T�3Hz��89��%�4�3%G��W�0�W�RdD�Z��Tܳ��K�a�3d��$cV 2!���1��I1H�0U2K2sk3K3J ci�aI�i�a�L��SLL��R$Vؠ�BV�E�Vk�]V*R��� � ,6Lc���9V2F{/P�:B��PS_�E���$rr�C�ѳ$A0��wPR���v�U�c�Sk�� {��8��� 0���VX`�!�tX`A��0P�Ё�
�5�SK!� �-qRH��!0���z�NJ SAX�!h�A�@LlA���A�THIC�1p�������1TFE��|�q>�IF_CH�3�A�I0�����G1@�x������9�Ɇ7_JF҇PR(����RVAT��� �-p��7@����D9O�E��COU(���AXIg��OFF{SE+�TRIG�S K��c���Ѽ�e�[�K��Hk���8�IGMA�o0�A-��ҙ�OR?G_UNEV���� �S�쐮d� �$������GgROU��ݓTO2���!ݓDSP��JO1G'��#	�_P'�2�OR���>P6KE�Pl�IR�0�PML�RQ�AP�Q��E�08q�e���SYSG��"v��PG��BRK*Rd�r�3�-��������ߒ<pAD�ݓJ�B�SOC� N�D?UMMY14�p\@�SV�PDE_OP�3SFSPD_O+VR��ٰCO��&"�OR-��N�0.��Fr�.��OV�S!Fc�2�f��F��!�4�S��RA�"LCH�DL�RECOV(��0�W�@M�յF�RO3��_��0� @�ҹ@VE}RE�$OFS�@3CV� 0BWDG�Ѵ`C��2j�
�TR�!���E_FDO>j�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�<#�8$CA�{�|����8$HBK|1,c��IO��.�:!aPPA"�N�3�^��F���:"�DVC_DB�C��d�w"���D�!��1���ç�3��^��ATIO� �q�0�UC�&CAB�BS�PⳍP��䖁�_0c�SUB'CPUq��S�Pa  aá�}0�Sb��c��r"~ơ$HW_C�����:c��IcA�A-�l_$UNIT��l���ATN�f����CY{CLųNECA���[�FLTR_2_�FI���(��}&��L�P&�����_SCT@SF_��F����G����FS|!�¹�CH�AA/����2��RSD�x"ѡb�r�: ;_T��PRO��OÖ� EM�_��8u�q u�q���DI�0e�RAIL�AC��}RMƐLOԠdC��:anq��wq�����PR��SLQ��pfC��30	��F�UNCŢ�rRIN�kP+a�0 ��!RA� >R 
Я��ίWAR�BLFQ��A������DA�����L�Dm0�aB9��nqBTIvrbؑ��μPRIAQ1�"AFS�P�!�����`(%b���M�I1UÇDF_j@��y1°L�ME�FA�@HRDiY�4��Pn@RS@Q��0"�MULSE�j@f�b�q �hX��ȑ���$.A[$�1$c1Ó~���� x~��EG�0ݓ�q!AR����09>B�%AXE��ROB���W�A4�_�-֣S�Y���!6��&S�'W�R���-1���ST�R��5�9�E��C 	5B��=QB90`�@6������OT�0�o 	$�ARY�8�w20���	%�F�I��;�$LINQK�H��1�a_63��5�q�2XY�Z"��;�q�3@��1��2�8{0B�{`D��� CFI���6G��
�{�_J���6��3aOP_dO4Y;5�QTBmAd"�BC
�z�DU"�z66CTURN3��vr�E�1�9�ҍGFL�`���~ �@�5<:y7�� 1�?0%K�Mc�68Cb�8vrb�4�ORQ��X �>8�#op������wq�Uf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W�� �Tυ� ;����QH� !`�ҽ��U�Q�WkeK#�kecXER��	BGE	0��S�dAWa Ǣ:D���7!�!AX�rB!{q��1 uy-!y�pz�@ z�@z6Pz\Pz�  z1v�y�y� +y�;y�Ky�[y��ky�{y��y�q�yD7EBU��$�����L�!º2WG`  A!B!�,��SV���� 
w���m���w� ���1���1���A���A ��6Q��\Q���!�m@���2CLAB3B��U�����S � ÐER���� �� $�@� Aؑ!p�PO��Z�q0�w�^�_MRAȑ�/ d  T�-��ERR��TYz�B�I�V3@�cΑ'TOQ�d:`L� �d�2�]�X�C[! /� p�`T}0i��_V1�r�a'�
4�2-�2<����@Pq�����F�$W���g��V_!�l�$��P����c��q"�	��SFZN_C;FG_!� 4��?� ��|�ų����@�ȲW� p ��\$� � n���Ѵ��9c�Q��(��FA�He�,�XE�DM�(�����!s��Q�g�P{RV HEL}Lĥ� 56��B_BAS!�RSQR��ԣo �#S��T[��1r�%��2ݺU3ݺ4ݺ5ݺ6ݺ�7ݺ8ݷ��ROO0I䰝0�0NLK!�C�AB� ��ACK��IN��T:�1�@p�@ z�m�_PU!�CO� ��OU��P�� Ҧ) ��޶��T�PFWD_KAR�ӑ�@��RE~��P8��(�QUE������P
��CSTOPI_AL�����0&p���㰑�0SEMl�db�|�M��d�TY|�3SOK�}�DI����p�(���_TM\�MANRQ�ֿ0E�+�|�$KEYSWITCH&	����HE
�BEAT4��cE� LEҒ��
�U��FO�����_O_HOM�O�7REF�PPRz�(�!&0��C+�OA��ECO��B�rI�OCM�D8׵�p]���8�` � D�1$����U��&�MH��<�P�CFORC���� ��OM�  �� @V��|�U�,3P� 1-�`� 3�-�4�]�NPXw_ASǢ� 0Ȱ�ADD����$S�IZ��$VAR\ݷ TIP]�\�
2�A򻡐���]�H_� �"S꣩!Cΐ���FRIF⢞�S0�"�c���NF��V ܻ�` � x�`SI��TES�R6SSG%L(T�2P&��AxU�� ) STMTQ2ZPm 6BW�P*�SHOWb��S�V�\$�� ���A00P�a�6���@�J�T�5��	6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	 f0u�	�0u�	�@uP[Pu%121?U1L1Y1f1sU2�	2�	2�	2�	U2�	2�	2�	2U22%222?U2L2Y2f2sU3P)3�	3�	3�	U3�	3�	3�	3U33%323?U3L3Y3f3sU4P)4�	4�	4�	U4�	4�	4�	4U44%424?U4L4Y4f4sU5P)5�	5�	5�	U5�	5�	5�	5U55%525?U5L5Y5f5sU6P)6�	6�	6�	U6�	6�	6�	6U66%626?U6L6Y6f6sU7P)7�	7�	7�	U7�	7�	7�	7U77%727?U7,i7Y7Fi7s۟'��VP�UP}D��  ��x|�԰��YSLOǢ� � z��и� ��o�E��`>�^t��А�ALUץ����CU����wFOqID_L��ӿuHI�zI�$FILE_���t�ĳ$`�JvSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_ �TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅�%L~�_Vj��+p�ޠ�� ` �GR�OU�pD��B�N�FLIC��RE�QUIREa�EB�UA��p����2��������c��{ \��APPR��iC���
�EN��CLOe��S_M� v�,ɣ�
���7� ��MC�&����g�_MG�q�C�� �{�9���|�BRKz�NOL��|ĉ R��_LI|��Ǫ�k�J����P
���ڣ������&���/���6��6��8������� ��8�%��W�2�e�PATH a�z�p�z�=�vӥ�ϰm�x�CN=�CA������p�IN�UCh��bq��CO�UM��!YZ������qE%����2������PAYL�OA��J2L3pR'_AN��<�L��F��B�6�R�{�R_F2�LSHR��|�LO�G��р��ӎ���ACRL_u�������.�r��H�p�$H{�^��FLEX
�s�}J�� :� /����6�2�����;�M�_�F16����n�@��������ȟ��Eҟ �����,�>�P�b� ��d�{�������������5�T��X ��v���EťmF ѯ�������&��/�A�S�e�D�Jx�� � ������j��4pAT����n�EL�  �%øJ���vʰJE��CTR�і��TN��F&��H�AND_VB[�
�pK�� $Fa2{�6� �rSWi��C�U��� $$	Mt�h�R��08��@<b 35��^6A�p3�kƈ�q{9t�A�̈p��A���A�ˆ0��U���D*��D��P��G��ICST��$A��$AN��DYˀ�{�g4�5D� ��v�6�v��5缧�^�@��P������#�,�5�>�(#�� &0�_�ER!V9�SQOASYM��] ��¤��x��ݑ���_SHl�������sT�(����(�:�JA���S�pcir��_VI�#�Oh9�``V_UN!I��td�~�J���b �E�b��d��d�f��n���������uN$���r��H����3��"CqEN� a�DI��>�ObtC�DpNx�� ��2IxQA����q��-��s �p� ����� ��/OMME��r4r�QTVpPT�P ���qe�i����P�x� ��yT�Pj� $DUMMY9��$PS_��RF�q�  ��:� p���!~q� X�����K�STs�ʰS�BR��M21_V�t�8$SV_ER�t�O��z���CLR�x�A  O�r?p? O�ր � D �$GLOB���#LO��Յ$�o��P�!SYSADR��!?p�pTCHM0 �� ,����W7_NA��/�e��$%SR��l (:]8:m�K6� ^2m�i7m�w9m��9�� �ǳ��ǳ���ŕߝ�9 ŕ���i�L����m��_�_�_�TD�XS�CRE�ƀ�� f��STF���}�pTТ6�B��] _v �AŁ� T����TYP�r�K��u�!�u���O�@ISb�!��tC�UE{tG� ����H�S����!RSM_�XuU?NEXCEPWv��CpS_��{ᦵ�ӕ�p��÷���COU ���� 1�O�U�ET�փr���PR�OGM� FLn!7$CU��PO*q���c�I_�pH;� �� 8��N�_HE�
p��Q��pRY ?���,�J�*���;�OUS�� �� @d���$B�UTT��R@���C�OLUM�íu�S�ERVc#=�PAN�Ev Ł� � N�PGEU�!�F��~9�)$HELP��^WRETER��)� ����Q�������@� P�P �IN��s�PNߠw v��1����� ����LN�� �䟀�_��k�$H��M TEX�#�����FLAn +REL�V��D4p�������M��?,��ӛ$�����P=�USR�VIEWŁ� <�d��pU�p0NFyIn i�FOCU��ni�PRILPm+��q��TRIP)��m�UNjp{t� �QP��XuWARN|Wud�SRTOLS��ݕ�����O|SO;RN��RAUư��9T��%��VI|�zu�� $�P�ATHg��CAC�HLOG6�O�LIMybM���'��"��HOST6�!��r1�R�OBOT,5���IMl� D�C� g!��E�L���i��VCPU_AVA�ILB�O�EX7�!BQNL�(���A�� Q���Q ��ƀ��  QpC���@_$TOOL6�$��_JMP� �<I�u$SS�!&�; SHIF��|s�P�p�6�s���R����OSURW�pRADIz��2�_�q�h�g! �q)��LUza$OUTPUT_BM��IML�oR6(`)��@TIL<SCO�@Ce�;��9�� F��T��a��o�@>�3�����w�2u1V�zu��%�D�JU��|#�WA�IT������%�ONE��YBO�ư �� �$@p%�C�SBn)T;PE��NEC��x"p�$t$���*B_T��R��%�qR� ���s	B�%�tM�+��t�.`�F�R!݀��OPm�wMAS�_DOG�OaT	�D����C3�S�	�O2DELAY���e2JO��n8E� �Ss4'#J�aP6%�����Y_��O2� �2����5��`? �-��ZABCS��  $�2��J��
B��$$CLA}S�����A�B�sp'@@VIRT8��O.@ABS�$��1 <E�� <  *AtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@��R�d�v�����M@[�A�XLր�&A�dC  ���IN��ā��GPRE������LARMRECOV <I䂥��NG�� \K	 A   J�\�M@�PPLIC�?�<E�E�H�andlingT�ool �� 
�V7.50P/2�8[�  �Pv��
�_SW��w UP*A� ��#F0ڑ����AG@��? 20��*A媗�:����[�FB 7D�A5�� '@�P@��Ngone������ ��Twk*A�4	Oxl�_���V����g�U�TOB�ค����HGAPON8@��LAz��U��D 1<EfA�����x����� Q 1שI Ԁ��Ԑ��:�i�n����#B=GB ���\��HE�Z�r�HTTHKY��$BI�[� m�����	�c�-�?� Q�o�uχϙϫϽ��� �����_�)�;�M�k� q߃ߕߧ߹������� �[�%�7�I�g�m�� ������������W� !�3�E�c�i�{����� ����������S/ A_ew���� ���O+=[ as������ �K//'/9/W/]/o/ �/�/�/�/�/�/�/G? ?#?5?S?Y?k?}?�? �?�?�?�?�?COOO 1OOOUOgOyO�O�O�O �O�O�O?_	__-_K_Q_��(�TO4�s����DO_CLEAN���e��SNM  9� �9oKo]o�oo�o�DSPDR3YR�_%�HI��m@&o�o�o#5G Yk}����"���p�Ն �ǣ�q�XՄ��ߢ��g�PL�UGGҠ�Wߣ��P�RC�`B`9���o�=�OB��oe�SEGF��K������ o%o����#�5�m���LAP�oݎ���� ������џ������+�=�O�a���TOT�AL�.���USE+NUʀ׫ �X����R(�RG_STR�ING 1��
_�M��Sc��
��_ITEM1 �  nc��.� @�R�d�v��������� п�����*�<�N��`�r�I/O �SIGNAL���Tryout �Mode�In�p��Simula�ted�Out���OVERR~�` = 100��In cycl����Prog OAbor����ĿStatus�	�Heartbea�t��MH Fa�ulB�K�Aler Uم�s߅ߗߩ߻���p������ �S ���Q��f�x��� ������������,� >�P�b�t�������,�WOR������V�� 
.@Rdv� ������p*<N`PO�� 6ц��o���� �//'/9/K/]/o/ �/�/�/�/�/�/�/�/�DEV�*0�? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O�qO�O�O�OPALTB��A���O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o�OGRI�p��ra�O Lo�o�o�o�o�o�o *<N`r��@����`o��RB� ��o�>�P�b�t��� ������Ώ������(�:�L�^�p����PREG�N��.���� ����*�<�N�`�r� ��������̯ޯ����&����$ARG�_��D ?	����i��  	$��W	[}�]}�������\�SBN_CONFIG i�������CII�_SAVE  ��۱Ҳ\�TCE�LLSETUP �i�%HOM�E_IO�͈�%�MOV_�2�8�R�EP���V�UTOoBACK
�ƽ�FRA:\��� �Ϩ���'�` ��������� ����$�6�c�pZ�lߙ��Ĉ���� ���������!凞�� M�_�q����2��� ������%�7���[� m��������@��������!3E$��� Jo�������WINI�@��ε���MESSAG�����q��ODEC_D$���O,0�.��PAUS�!��i� ((O l��������  /�//$/Z/H/~/�l/�/�'akTSK�  q�����UgPDT%�d0~;WSM_CF°�i�еU�'1G�RP 2h�93 �|�B��A�/S�XS�CRD+11
1; ����/�?�? �? OO$O��߳?lO ~O�O�O�O�O1O�OUO _ _2_D_V_h_�O	_|X���GROUN0|O�SUP_NAL��h�	�ĠV_E�D� 11;
 ��%-BCKED�T-�_`�!oEo$�A��a��o����Y�ߨ���e2no_˔o�o�b���ee�o8"�o�oED3�o��o ~[�5GED4�n#�� ~�8j���ED5Z���Ǐ6� ~���}���ED6����k�ڏ ~G�8��!�3�ED7��Z���~� ~�V�şןE�D8F�&o��Ů�}����i�{�ED9ꯢ�W�Ư
}3�����CRo����π3�տ@ϯ����P�PN�O_DEL�_�RGE_UNUSE�_��TLAL_OUT� q�c�QWD_ABOR� �΢Q���ITR_RTNz����NONSe����CAM_�PARAM 1��U3
 8
S�ONY XC-5�6 234567w890�H � @���?��ҟ( АV�|[�r؀~�X�HR5�k�|U�Q�߿�R57�����Aff���KOWA SC3W10M|[r�̀�d @6�|V ��_�Xϸ���V��� ����$�6��Z�l��CE_RIA_I8�57�F�1���R|]��_LI�O4W=� ��P<z~�F<�GP 1�,���_GY<k*C*  ���C1� 9� @� G�� �CLC]� d*� l� s�R� ���[�m� v� �� �� �� C��� �"�|W��7�H=EӰONFI� ���<G_PRI 1�+P�m®/���������'CH�KPAUS�  1E� ,�>/P/ :/t/^/�/�/�/�/�/ �/�/?(??L?6?\?4�?"O�����H^�1_MOR��� �0�5 	  �9 O�?$OOHO6K�2D	���=9"�Q?5�5��C�PK�D3P������a�A-4�O__|Z
�O G_�7�PO�� ��6_��Y,xV�ADB���=�'�)
mc:cpmidbg�_`��S�:�  ��P�ļ��Up�_)o�S  �  A����R�P�_mo8j��"��Koo�o9i�(�Փog�o�o�m���of�oGq:I�ZD�EF f8��)��R6pbuf.t�xtm�]n�@�����# 	`(Ж�A=�L���zMC�21��=��9���4��=�n׾�Cz  �BHBCCo�C�|��CqD���C���C��{iSZE@D����F.��F���E⚵F,�E�ٙ�E@F��N�IU��I?�O�I<#I6?�I�SY��)�vqG���Em�U(�.��(�(�1�<�q�G�x2��eҢ �� a�D�j�怀ES\E@EX��EQ�EJP� F�E�F�� G�ǎ^F� E�� FB�� H,- Ge�߀H3Y��� � >�33 9���xV  n2xQ�@��5Y��8B� A��AST<#�
� ��_'�%��wRSMOFS���~2�y�T1�0DE ��O@b 
�(�;��"�  <�6�z�Rb���?�j�C4�)�SZm� W��{�Jm�C��B-G�Cu��@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"�� , 
�^��P�o xvf`MT�I^��rl@�:sONTImM������Zv�i
õ�cMOTN�END���dREC�ORD 1(R�8a��ua�O��q� �sb�.�@�R��xZ� ������ɏۏ폄� ��#���G���k�}��� ��<�ş4��X��� 1�C���g�֟������ ��ӯ�T�	�x�-��� Q�c�u���������� >����)Ϙ�Mϼ� F�࿕ϧϹ���:��� ����%�s`Pn&�]�o� �ϓ�~ߌ���8�J��� ��5� ��k����� ���J�����X��|� ��C�U�����������0�����	��dbTOLERENCqdsBȺb`L�͐P�CS_CFG �)�k)wdMC�:\O L%04dO.CSV
�Pc��)sA �CH� z�P)~���hM�RC_OUT �*�[�`+P SG�N +�e�r���#�10-MAY�-20 09:0�7*V17-FEB�j1o9�k PQ�8��)~��`pa�m���PJPѬV�ERSION �SV2.0�.8.|EFLOG�IC 1,�[ 	DX�P7)�PF.�"PROG_ENqB�o�rj ULSew� �T�"_WRS�TJNEp�V�r`dE�MO_OPT_S�L ?	�es
 	R575)s 7)�/??*?<?'�$TO  �-��?�&V_@pEX�Wd��u�3PATH ;ASA\�?�?\O/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C���SqqF�PMAqU� t/XrMSWR�.�i6.|S/�Z!D_N�O0__T_�C_x_g_�_�tSBL__FAUL"0�[^3wTDIAU 16M�6p�A1�234567890gFP?BoTo foxo�o�o�o�o�o�o �o,>Pb�SZ�pP�_ ���_ s�� 0`���� �)�;�M�_�q����������ˏݏ��|)U3MP�!� �^��TR�B�#+�=�PM�EfEI�Y_TEM=P9 È�3@�3�A v�UNI�.(Y�N_BRK 2�Y)EMGDI_�STA�%W!bՐN�C2_SCR 3��1o"�4�F�X� fv���������#��ޑ14����)��;�����ݤ5�����x�f	u�ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/߭P�b�t��  ��xߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N���r������� ��������&8 J\n����� ���"`�FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/4 ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O?�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�O�O�o�o�o 
.@Rdv� �������� *�<�N�`�r����o�� ��̏ޏ����&�8� J�\�n���������ȟ�ڟ����H�ETM�ODE 16��]� ��ƨ�
R�d�v�נRRO�R_PROG �%A�%�:߽�  ���TABLE  A������#�L��RRSEV_NU�M  ��Q���K�S���_AU�TO_ENB  q��I�Ϥ_NOh�� 7A�{�R��  *������������^�+��Ŀֿ迄�HISO�͡I��}�_ALM 18.A� �;�����+�e�wωϛϭ����_H���  �A���|��4�TC�P_VER !�A�!����$EXTLOG_REQ�s�{�V�SIZ_�~Q�TOL  ͡{Dz��A Q�_BWD����r����n�_DI�� 9��}�z�͡m���STEP����4��_OP_DO����ѠFACTORY�_TUN�dG�E�ATURE :�����l�H�andlingT�ool ��  -� CEngl�ish Dict�ionary��O�RDEAA �Vis�� Mas�ter���96 �H��nalog �I/O���H55�1��uto So�ftware Update  ���J��matic �Backup��P�art&�gr�ound Edi�t��  8\ap�Cameraz��F��t\j6R��ell���LOA�DR�omm��sh�q��TI" ��cyo��
! o����pane�� �
!��tyle select��H59��nD���o�nitor��48�����tr��Rel�iab���adi�nDiagn�os"����2�2 u�al Check� Safety �UIF lg\a���hanced �Rob Serv> q ct\��lUser FrU���DIF��Ext�. DIO ��f�iA d��en]dr Err L@���IF�r��  �П�90��FCT�N MenuZ v�'��74� TP �In��fac � SU (G�=�p��k Exc�n g�3��Hig�h-Sper Sk]i+�  sO�H9 ~� mmunic!��onsg�teurh� ����V����^conn��2��{EN��Incr�stru���5.�fdKARE�L Cmd. L�?uaA� O�R�un-Ti� EnIv����K� ��+%��s#�S/W��74���License|T�  (Au* �ogBook(S�y��m)��"
�MACROs�,V/Offse6��ap��MH� �����pfa5�Mec�hStop Pr3ot��� d�b =i�Shif���/j545�!xr ��#��,^b o�de Switc]h��m\e�!oz4.�& pro��4��g��Mul�ti-T7G��n�et.Pos Regi��z�}P��t Fun����3 Rz1��Nu!mx �����9m�1>�  Adjuj��O1 J7�7�* ��<���6tatuq1EIKRDMt�ot��scove�� ��@By- }Ouest1�$Go� �� U5\SNPX b"���YA�"Libr����#b�� �$~@h�pd]0��Jts in VCCM�����0�q  �u!��2 R�0��/I�08��T�MILIB�M J�92�@P�Acc�>�F�97�TPT�X�+�BRSQelZ0�M8 Rm��q%��692��Une�xceptr mo�tnT  CVV�P���KC����+�-��~K  II)��VSP CSXC��&.c�� e�"�� =t�@Wew�gAD Q�8bvr �nmen�@�iP�� a0y�0�pfG�ridAplay !� nh�@*�3R�1�M-10iA(B�201 �`2V" y F���scii��load��83 �M��l����Gua=r�d J85�0�maP'�L`���stua�Pat�&]$Cyc8���|0ori_ x%oData'Pqu���ch�1��g`� mj� RLJam�5����IMI De�-B(\A�cP" #�^0C  etk}c^0asswo%q.�)650�ApU��Xnt��Pven��CTqH�5�0�YELLOW BqO?Y��� Arc�0�vis��Ch�W�eldQcial44Izt�Op� ��gs�` 2@�a��p�oG yRjT1� NE�#HT� xyWb��! �p�`!gd`���p\� =P���JPN ARCP�*PR�A�� �OL�pSup̂f�il�p��J�� ��cro�670�1C~E��d��SS�pe�t�ex�$ �P� Soz7 t� ssagN5� <Q�BP:� �9 �"0�QrtQC��P�l0dpn�笔�r�pf�q�e�ppm�ascbin4p�syn�' ptx�]08�HELNC�L VIS PK�GS �Z@MB �&��B J8@I�PE GET_V�AR FI?S (�Uni� LU�OO�L: ADD�@2/9.FD�TCm���E�@DVp���`A��ТNO WTWTOEST �� &�!���c�FOR ��E�CT �a!� AL�SE ALA`�CPMO-130���� b D: HAN?G FROMg���2��R709 D�RAM AVAI�LCHECKS �549��m�VPC�S SU֐LIM�CHK��P�0x�F_F POS� F��� q8-12� CHARS�ER>6�OGRA ��Z@wAVEH�AME��G.SV��Вאn$���9�m "y�TR}Cv� SHADP��UPDAT k�0>��STATI���? MUCH ����TIMQ MOTN-003��@�OBOGUIDE? DAUGH���b8��@$tou� �@�C� �0��PATH|�_�MOVET��� R64��VMX�PACK MAY ASSERTjS޴�CYCL`�TA���BE COR �71�1-�AN��R�C OPTION�S  �`��APSwH-1�`fix��2�SO��B��XO򝡆��_T��	�i��0j���du�byz p cwa��y�٠HI������U�pb XSP�D TB/�F� \�hchΤB0���EmND�CE�06\Q��p{ smay In@�pk��L ���traff#�	� ���~1from �sysvar s�cr�0R� ��d�DJU���H�!A���/��SET ER�R�D�P7����N�DANT SCR�EEN UNRE�A VM �PD�D���PA���R�I�O JNN�0�F�I��B��GROUNנD Y�Т٠��h�SVIP 5�3 QS��DIGI?T VERS��k���NEW�� P0�6�@C�1IMAG��ͱ���8� DIx`���pSSUE�5���EPLAN J=ON� DEL���1�57QאD��CALLI���Q��m����IPND}�IMG� N9 PZ�19޴�MNT/��ES� ���`LocR HCol߀=��2�Pn� �PG:��=�M��c�an����С: �3D mE2vie�w d X��e�a1 �0b�pof �Ǡ"HCɰ�AN�NOT ACCE�SS M cpite$Et.Qs a� {loMdFlex)a�:��w$qmo G
�sA9�-'p~0��h0�pa��eJ AU�TO-�0��!ip�u@Т<ᡠIABL�E+� 7�a FPL�N: L�pl lm� MD<�VI�����WIT HOCv�Jo~1Qui�t�"��N��USB�@��Pt & rem�ov���D�vAxi�s FT_7�PG�ɰCP:�OS-�144 � h s� 268QՐOST��p  CRASH� DU��$P��W�ORD.$�LOgGIN�P��P:	��0�046 iss�ueE�H�: Solow st��c�`6����໰I�F�IMPR��SPOT:Wh4���N1�STY��0VMGqR�b�N�CAT��-4oRRE�� � 58�1��:%�R�TU!Pe -M a�SE:�@pp���AGp�L��m@al�l��*0a�OCB �WA���"3 CN�T0 T9DWro>O0alarm�ˀm0d t�M�"0�2�|� o�Z@OME�<�� ��E%  #1�-�SRE��M�st�}0g     �5KANJI5n�o MNS@�I�NISITALI�Z'� E�f�we���6@� dr�@ f�p "��SCII� L�afails� w��SYSTaE[�i��  � tMq�1QGro8�m n�@vA����&���n�0q��RWR=I OF Lk���� \ref"�
�u�p� de-rel}a�Qd 03.�0�SSchőbet�we4�IND e�x ɰTPa�DOȬ l� �ɰGi�gE�soperawbil`p l,��aHcB��@]�le�Q0cflxz�Ð���OS {����v4pwfigi GLA�$��c2�7H� la�p�0ASB� Ifz��g�2 l\c�0��/�E�� EX'CE 㰁�P���$i�� o0��Gd`]���fq�l lxt��EFal��#0��i�O�Y�n�CLOSn��SRNq1NT^��F�U��FqKP�AN�IO V7/ॠ1p�{����DB �0ء�ᴥ�ED��DE�T|�'� �bF�N�LINEb�BUG�T���C"RLIB���A��ABC J�ARKY@��� r7key�`IL���P�R��N��ITGAR
� D$�R �Er�� *�T��a�U�0��h�[�ZE V� �TASK p.vr�P2" .�XfJ��srn�S谥dIB�P	c���B/��B�US��UNN�  j0-�{��cR'���LOE�DIVS�C�ULs$cb����BW!��R~�W`P���&��IT(঱tʠ�{OF��UNEXڠ�+���p�FtE��S�VEMG3`NML� 505� D*�C?C_SAFE�P*�p �ꐺ� PET��8'P�`�F  !���IR����c i S�>� K��K�H �GUNCHG��S^�MECH��M��T*�%p6u��tP�ORY LEAKr�J���SPEg�D��2V 74\G�RI��Q�g��CTLN��TRe @�_��p ���EN'�IN�������$���r��T�3)�i�STO�A$�s�L��͐X	����q��Y� ��TO2�J m��0F<�K�����DU�S��O��3$ 9�J F�&�����SSVGN-18#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRKC�TR/"� �q\j5���_�Q�S�qINVJ0D ZO�Pݲ�� �s��г�Ui ɰ̒�a��DUAL� J�50e�x�RVO1/17 AW�TH!�Hr%�N�247%�5q2��|�&aol ���R���at�Sd�cU8���P,�LER��i�x�Q0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�cб���{�U��RO�P 2�b�pB��ITP4M��b !�AUt c0< � pl�ete�N@� �z1^qR635 (�AccuCal2zkA���I) "�(ǰ�1a\�Ps��ǐ � bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etaca2��AT���PC�`��슰�_p�.pc�!Ɗ��:�circB���5�tl��Bɵ��:�fm+�Ί�V�b��ɦ�r�upfrma.����ⴊ�xed�8�Ί�~�pedA�D ��}b�ptlib0B�� �_�rt�߄	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆�D����c�Ӳ�5�j>ʌ����tcȐ��	�r(����mm 1��T�#sl^0��T�mѡ�&#�rm3��ub Y��q�std}��pl�;�&�ckv�=�r�vaf�䊰��9�vi������ul�`�0fp�q� �.f��� d�aq; i Data� Acquisi
��n�
��T`���1�89��22� DMCM RR[S2Z�75��9 ?3 R710�o�59p5\?��T{ "��1 (D�T� nk@���������E Ƒȵ��Ӹ�et3dmm ��ER����gE��1�q\mo?۳�=(G����[(

�2�` ! ��@JMACRO���Skip/Of�fse:�a��V�4�o9� &qR662����s�H�
 6�Bq8����9Z�4_3 J77� 6�J783�o ���n�"v�R5IK�CBq2 PTLC�Zg R�3 (�s, ��������03�	зJԷ\�sfmnmc "MNMC����ҹ�%wmnf�FMC"�Ѻ0ª etmcr�� �8����� ,^D&^�   874�\prdq>,jxF0���axisH�Process �Axes e�rol^PRA
�Dp� �56 J81j�5-9� 56o6� ��l�0w�690 98� �[!IDV�1��2(8x2��2ont�0�
 ����m2���?C���etis "I�SD��9�� FpraxRAM�P� D��defB�,�G�isbasicH�B�@޲{6�� 70U8�6��(�Acw: ������D
�/,��AMOX�� ��DvE��?�;T��>Pi� RAFM';�]�!PAM�V�W��Ee�U�Q'
bU�7y5�.�ceNe� �nterfaceh^�1' 5&!54�K<��b(Devam±��/�#���/<�Tane`"DNEWE���btpdnui �A�I�_s2�d_rsCono���bAsfj|N��bdv_arFv�f�xhpz�}w��hkH9xstc��gAp�onlGzv{�ff ��r���z�3{�q'Td>pcha�mpr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�!��pcchmp]aM�P&B�� �mpe�v�����pcs���YeS�� MacKro�OD��16Q! )*�:$�2U"_,��Y�(PC ��$_;�������o��J�geg{emQ@GEMSW�|~ZG�gesndy�<�OD�ndda��Sƕ�syT�Kɓ�su^Ҋ���n�m���L��O  ���9:p'�ѳ޲��spotplusp���`-�W�l�J�s��t[�׷p�key�ɰ�$��s��-Ѩ�m���\fea;tu 0FEAWD�oolo�srn '!2 p���a�As3���tT.� (N. A.)��!e!(�J# (j�,��o�BIB�oD -�.�n6��k9�"K��u[�-�_���p� "P�SEqW����wop "sEЅ�&�:� J������y�|��O8� �5��Rɺ���ɰ[� �X�������%�(
 ҭ�q HL�0k� 
�z�a!�B�Q�"(g�Q�����]�'� .�����&���<�!ҝ_�#��tpJ�H�~Z�� j�����y������2 ��e������Z����V� �!%���=�]�͂���^2�@iRV� on��QYq͋JF0� 8�ހ�`�	(^�dQueue���X\1����`�+F1tpvtsen��N&��ftpJ0v �RDV�	f���J1 Q���v�eyn��kvstk���mp��btkcl�rq���get�����r��`k�ack�XZ�st1rŬ�%�stl��~Z�np:!�`�� �q/�ڡ6!l�/Yr$�mc�N+v3�_`� ����.v�/{\jF��� �`�Q�΋ܒ�N50 (�FRA��+��͢f?raparm��Ҁ��} 6�J643�p:V�ELSE
�#�VAR $SG�SYSCFG.$��`_UNITS �2�DG~°@�4Jgfqr��4A�@FRL-� �0ͅ�3ې���L�0 NE�:�=�?@�8�v�9~Qx304��;�B�PRSM~QA�5T�X.$VNUM_�OL��5��DJ50�7��l� Functʂ"qwAP��琉�G3 H�ƞ�kP9jQ��Q5ձ� ��@jLJ zBJ[�6N�kAP�����S��"TPPRp���QA�prna�SV�ZS��AS8Dj5k10U�-�`cr�`8 ��ʇ�DJR`jYȑH  �Qm �PJ6�a21���48AAVM3 5�Q�b0 lB�`�TUP xbJ�545 `b�`61�6���0VCA�M 9�CLI�O b1�5 ����`MSC8�
rP� R`\sSTYL MNIN�`oJ628Q  �`�NREd�;@�`SC�H ��9pDCSU� Mete�`OR�SR Ԃ�a04 �kREIOC ��a5�`542�b9 vpP<�nP�a�`�R�`�7�`�MAS�K Ho�.r7 <�2�`OCO :��r�3��p�b�p���r0�X��a�`13\mn��a39 HRM"��q�q��LCH}K�uOPLG B��a03 �q.�pH�CR Ob�pCpP�osi�`fP6 i=s[rJ554�òp'DSW�bM�D�pqR��a37 }Rjr0 L�1�s4 �R6�7���52�r5 �2�r7� 1� P6���Re�gi�@T�uF�RDM�uSaq%�4�`930�uSNB�A�uSHLB̀\�sf"pM�NPI��SPVC�J5�20��TC�`"M�NрTMIL�I=FV�PAC W�poTPTXp6.%��TELN N M�e�09m3U�ECK�b�`UFR��`��VCOR��V�IPLpq89qSX9C�S�`VVF�J��TP �q��R62]6l�u S�`Gސ~�2IGUI�C���PGSt�\ŀH863�S�q�����q�34sŁ684`���a�@b>�3 :B抂1 T��96 :.�+E�51 y�q353�3�b1 ���b31 n�jr9 ���`�VAT ߲�q75� s�F��`�sAWSyM��`TOP u��ŀR52p���a809 
�ށXY q���s0 ,b�`885�QXрOLp}�"pE�v��tp�`LCMDў�ETSS���6� �V�CPE o�Z1�VRCd3
�NuLH�h��001m2�Ep��3 f��p��4� /165C��6�l���7PR��00�8 tB��9 -2[00�`U0�pF�1&޲1 ��޲2L"����p��޲4��5 �\hmp޲6 RB�CF�`ళ�fs�8� �Ҋ��~�J�7 OrbcfA�L�8\P0C����"�32m0u��n�K�Rٰn�5 5oEW
n�9 zΊ�40 kB��3 ��6ݲ�`00iB%/��6�u��7�u���8 µ������sU0��`�t �1 05\;rb��2 E��K���j���5˰��6A0��a�HУ`:�63�`jAF�_���F�7 ڱ�݀H�8�eHЋ��cUI0��7�p��1u��8u��9 73�������D7� ��5\t�97 ��8U�Q1��2��1�1:����h��1np�"��8�(�U1��\pyl���,࿱v ��B�85E4��1V���D�4��im��1�<���$>br�3pr�4@pGPr�6 B���цp���1����1�`͵15=5ض157 �2�у62�S����1�b��2����1Π"�2L���B6`�1<cf�4 7B�5 DR���8_�B/��18�7 uJ�8 06��90 rBn�1 �(��202 0E�W,ѱ2^��2��9�0�U2�p�2��2 �b��4��2�a"RiB����9\�U2�`xw�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`ڰR,:7 �2��V�2��5���2^��a^9���qr�����n�5����5᥁"�8Ha�Ɂ}�5B���5������`UA���� ��8�6 �6 S�0��5��p�2�#�529 ��2^�b1P�5�~�2`���&P5���8��5��u�!�5\��ٵ544��5��	R�ąP nB^z�c (�4�����SU5J�V�5��1�1@^��%�����5 �b21��gA��5m8W82� rb��95N�E�5890r�: 1�95 �"�� ����c8"a��|�L (���!J"5|6��^!"�6��B�"8�`#���+�8%�6B�AM�E�"1 iC��622�Bu�6V��d� �4��84�`ANR�SP�e/S� �C�5� �6� ��� \@� �6� �V� 3t��?� T20CA�R���8� Hf� 1DH��� AOE� ��w ,|�� �0X\�� �!64K��ԓ�rA� �1 (M-7�!/50T�[PM��P�Th:1�C�#P�e� �3�0� 5`M�75T"� �D8p�! �0Gc� u�4��i1�-710i�1� S�kd�7j�?6�:-HS,� �RN�@�UB��f�X�=m75sA*A6an���!/CB�B2.6A �0;A�C�IB�A�2�QF1�UB2:�21� /70�S� �4����Aj1�3p����r#0 B2\m*A@C��;bi"i1K��u"A~AAU� imm7c7��ZA@I�@�Df�A�D5*A�E� #0TkdR1�35Q1�" *�@�Q�1�QC)P�1 *A�5*A�EA�5B�4>\77
B7=Q�D�2H�Q$B�E7�C�D/qA	HEE�W7�_|`jz@@� 2�0�Ejc7(�`�E"l7�@7�A
1��E�V~`�W2%Q�R9\ї@0L_�#��� �"A���b��H3s=rA/2�R5nR4�7�4rNUQ1ZU�A�s\m9
1M92L2�!F!t^Y�ps� 2ci��-?�qhimQ�t  w0 43�C�p2�mQ�r�H_ �H20�Evr�QHsXBFSt62�q`s����� ��Pxq350_�*A3I)�2�d�u0X�@� '4TX�0�pa3i1A3sQ25L�c��st�r�VR1%e�q0
��j1��O 2 �A�UEiy�.�‐� �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ�� qA!Pvs� 5	15aU ���?PŅ���ဝQG9A6�zS*�7�q�b5�1����Q��00	P(��V7]u�aitE1 ���ïp?7� !?�z���rbUQRB1P�M=�Qa9��H��QQ�25L�������Q���@L��8ܰ��y0�0\ry�"R2B�L�tN  ��w� �1D&^�2�qeR�5���_bx�3�X]1m1lcqP!1�a�E�Q� 5F����!5���@M-16 Q�� f���r��Q�e�� ��� PN�LT_`�1��i1��9453�p�@�e�|�b1l>�F1u*AY2�
��R8`�Q����RJ�J3�D}T� 85
Qg�/0�� *A!P�*A�Ð𫿽�Y2ǿپ6t�6=Q����Pȓ��� AQ� g�*ASt]1^u�a jrI�B����~�|I��b��yI�\m�Qb�I �uz�A�c3Apa9q� B6S��S��m����}�85`N�N�  �(M���f1����6����161��5�s`�SC��U��A�����5\set036c����10�y�#h8��a6��6��9r�2HS ���Er���W@}�a��I�lB� ��Y�ٖ�m�u�C������5�B��B��h `�F���X0���A:���C�M��AZ��@��4��6i����� e�O�- 	���f1��F ������1F�Y	���T6HL3��U66~`���Ur�dU�9D20Lf0 ��Qv� ��fjq��N� �����0v
� ��i	��	��72lqQ2�������� \chngmove.V���d���@2l_arf	�f~�� 6������9C�Z��0�~���kr41 S���0��V��t����8��U�p7nuqQ%��A]��V�1\�Qn�BJ�2W�E�M!5���)�#:�648��F�e50S�\� �0�=�PV���e�� ����E������m7shqQSH" U��)��9�!A��(����� ,s^�ॲTR1!�L��,�60e=�4F�d����2��	 R-�� ���������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2��"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D�� �5V��@2cVE��Ȗ�T��pt갖�1L ~E�#�F�Q��9E�#Dce/��RT��59�� �	�A�EiR�������9\m20�20 ��+�-u�19r4�`� E1�=`O9`�1"ae��O�2��_$W}am41�4�3�/d?1c_std��1�)�!�`_T��r�_ 4\jdg�a�q�P J%!~`-�r�+bg8B��#c300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W �"PsA��e��� �t�i�P�W.�� c�FX.�e�kE1�4�44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�A Pf��coWo!\�[2a��2A;_2��QW2�bF�(�V11ă23�`��X5�Ra2�1�J*9�a:88�J9X�l5�m1a`첚��*���(85�& �������P6����R,52&A����,8fA9IfI50\u�z��OV
�v��}E֖J0���Y>� 16r�C �Y��;��1��L���A q�&ŦP1��vB)e��m�����1p� .�1D&^�27�F��KAREL Us�e S��FCTN<��� J97�FA+�� (�Q޵�p%�L)?�Vj9F?(�j�R�tk208 "Km�6Q�y�j��iæP�r�9�s#��v�kr;cfp�RCFt3����Q��kcctme��!ME�g����6�mWain�dV�� ��Cru��kDº�c��0�o����J�dt�F9 �»�.vrT�f�����E%�!��5�FR�j73B�K���UtER�HJ�O  J��# (ڳF���F�q� Y�&T��p�F�z��19�tkvBr���V�h�9p�E�y�<�k������p��;�v���"CT�� f����)�
І��)� V	�6���!��qFF ��1q���=�����O�@?�$"���$��je����TCP Aut��r�<520 H5n�J53E193��9��96�!8��9���	 �B574��5�2�Je�(�� Se%!Y�����u��ma>�Pqtool�ԕ������conr�el�Ftrol �Reliable��RmvCU!��H51������ a55�1e"�CNRE ¹I�c�&��it��l\sfutst "UTա��"X�\u��g@�i�6Q]V�0�B,Eѝ6A�  �Q�)C���X��Yf�hI�1|6s@6i��T6IU��vR�d�
$ae%1��2�C58�E6��8�Pv�iV4OFH�58SOeJ� mvBM6E~O58�I�0�E �#+@�&�F�0���F �P6a���)/++�</>N)0\tr1������P ,^ɶ�rmwaski�msk�a$A���ky'd�h	A	��P�sDispla�yIm�`v����J887 ("A��+Hyeůצprds�ҨI�:���h�0pl�2"�R2��:�Gt�@��PRD�TɈ�r�C�@�Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@��^Sp��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@�P�firmQ����P@p�2�=bk�6�r�3��6��tppl��PAL���O�p<b�ac�q 	��g1J�U�d�J��gait_9e��Y��&��Q���	�Sha�p��eratio�n�0��R674�51j9(`sGen@�ms�42-f��r�p`�5����2�rsgl��E��p�G���qF�20�5p�5S���Ձ�re�tsap�BP�O�\}s� "GCR��z�? �qngda�AG��V��st2ax�U��Aa]��bad��_�btputl�/�&�e���tpli1bB_��=�2.����5���cird�v�sqlp��x�hex���v�re?�Ɵx�key�v�pm��x�sus$�6�gcr���F������[�q27j9�2�v�ollis�mqSk�9O�ݝ� �(pl.���t��p!o��29$Fo8��cg�7no@�tptcls` CLS�o�b�F\�km�ai_
�s>�v�o	�t�b���ӿ�E�H��6�1e_nu501�[m���utia|$cal�maUR��CalMwateT;R51%�i=1]@-��/V� ���Z�� �fq1�9 "�K9E�L����2m�CLMTq�S#��3et �LM3!}t �F�c�nspQ�<c���c_moq��� ��c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 �̆�N�ve��C�cl�m�&Ao# �|$fi�nde�0S�TD ter FiLANG���R��
��n3���z0Cen���r, ������J����� � ��K��Ú�=���_�����r� "FNCDR�� 3��f��tguid�䙃N�."��J�tq�� ��� ����������J����_������c��	m��Z��\fndrA.��n#>
B2p��>Z�CP Ma������38A��� c��6� (���N�B���@���� 2�$�81�B�m_���"ex� z5�.Ӛ��c��0bSа�efQ���	��RBT;�OPTN �+#Q� *$�r*$��*$r*$%/ s#C�d/.,P�/0*ʲDPN��$����$*�Gr�$k E�xc�'IF�$MA�SK�%93 H5��%H558�$548 H�$4-1�$�d�#1(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9j0�"M�49�4  ���4�4tpsh���4�P�4- DQ�� �3�Q�4�R�4�pR@%0�2�r�4.b
E\���5�A�4��3adq}\�5K979":E��ajO l "DQ ^E^�3i�Dq ��4�ҲO ?R�? ��q@�5��T��3rAq�OF�Lst�5~��7p�5`��REJ#�2�@av^E�ͱ�F���4��.�5y� N� �2il(iqn�4��31 JH1��2Q4�251ݠ�4r'mal� �3)�RE o�Z_�æOx����4��8^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4$�REM���4yݱ"u<@�RER5932fO��47Z��5lity�,�U��e"Dil�\�5��o ��79�87�?�25 �3hk910�3��FE�0�=0P_�Hl\mhm �5��qe�=$�^��
E��u�IAympt�m�U��BU��vst e�y\�3��me�b�Dv I�[�Qu�:F�Ub�*_0�
E,�su��_	 Er��ox���4huse�E-�?�sn�������FE��,�Gbox�����c݌ ,"�������z���M��g��pdspw )�	��9���b���(��1���c�� Y�R�� �>�P���W�@�������'�0ɵ��[��͂��� � � ,@�� �A�bu�mpšf��B*�BCox%��7Aǰ60�pBBw���MC� (6��,f�t I�s� ST��*��}B������w��"BBF�
�>�`���)��\�bbk968 "��4�ω�bb�9�va69����etb�Š��X�����ed�	�F��u�f� �s�ea"������'�\���,���b�ѽ�oH6�H�
�x�$�f����!y���Q[�! toperr�fd� �TPl0o� Rec�ov,��3D��R/642 � 0��C@�}s� N@��(U�rro���yu2r���  �
 � ����$$CL~e� ������������$z�_�DIGIT��������.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�o$j��+c:PR�ODUCTM�0\�PGSTKD��V�&ohozf99��D����$FEAT_INDEX���xd�� � 
�`ILEC�OMP ;����#��`�cSET�UP2 <�e��b�  N ��a�c_AP2BC�K 1=�i G �)wh0?{%&c����Q�xe% �I�m���8� �\�n����!���ȏ W��{��"���F�Տ j���w���/�ğS�� �������B�T��x� �����=�үa����� �,���P�߯t���� ��9�ο�o�ϓ�(� :�ɿ^���Ϗϸ� G���k� �ߡ�6��� Z�l��ϐ�ߴ���U� ��y����D���h� �ߌ��-���Q����� �����@�R���v�� ��)�����_����� *��N��r�� 7��m�&��3\�i
pP }2#p*.VRc�*��� /��PC/1/�FR6:/].��/+T�`�/�/F%��/�,�`r/?�*#.F�8?	H#&?�e<�/�?;STM� �2�?�.K �?�=�iPenda�nt Panel�?;H�?@O�7.O�?8y?�O:GIF�O�O��5�OoO�O_:JPG _J_�56_�O_�_��	PANEL1'.DT�_�0�_�_�?O�_2�_So�W Ao�_o�o�Z3qo�o@�W�o�o�o)�Z4�o�[�WI��
�TPEINS.XSML��0\����qCustom� Toolbar�	��PASSW�ORDyFR�S:\L�� %�Password Config�� �֏e�Ϗ�B0��� T�f����������O� �s������>�͟b� �[���'���K��� �����:�L�ۯp��� ��#�5�ʿY��}�� $ϳ�H�׿l�~�Ϣ� 1�����g��ϋ� ߯� ��V���z�	�s߰�?� ��c���
��.��R� d��߈���;�M��� q������<���`��� ����%���I������ ��8����n��� !��W�{" �F�j|�/ �Se��/�/ T/�x//�/�/=/�/ a/�/?�/,?�/P?�/ �/�??�?9?�?�?o? O�?(O:O�?^O�?�O �O#O�OGO�OkO}O_ �O6_�O/_l_�O�__ �_�_U_�_y_o o�_ Do�_ho�_	o�o-o�o Qo�o�o�o�o@R �ov��;�_ ���*��N��G� �����7�̏ޏm�� ��&�8�Ǐ\�돀�� !���E�ڟi�ӟ��� 4�ßX�j�������� įS��w������B��#��$FILE_�DGBCK 1=���/���� ( �)�
SUMMARY�.DGL���MD�:�����Di�ag Summa�ry��Ϊ
CONSLOG��������D�ӱConso?le logE�ͫ���MEMCHECCK:�!ϯ���X��Memory D�ata��ѧ�{�)��HADOW�ϣϵ�J���Sh�adow Cha�ngesM�'�-��)	FTP7�Ф�3ߨ���Z�mment TBD���ѧ0=4)ET?HERNET��������T�ӱEth�ernet \�f�iguratio�nU�ؠ��DCSV�RF�߽߫������%�� veri?fy all��'��1PY���DIF�F�����[���%=��diff]�������1R�9�K���c ���X��CHGD������cB��r����2Z8AS� ��GD���k��qz��FY3b8I[� �/"GD���s/�����/*&UPDATES.� �/��?FRS:\�/�-�ԱUpdate?s List�/���PSRBWLD.CM(?���"<?�/�Y�PS_ROBOWEL��̯�?�?� �?&�O-O�?QO�?uO OnO�O:O�O^O�O_ �O)_�OM___�O�__ �_�_H_�_l_o�_�_ 7o�_[o�_lo�o o�o Do�o�ozo�o3E �oi�o���R �v���A��e� w����*���я`��� ������O�ޏs�� ����8�͟\����� '���K�]�쟁���� 4���ۯj������5� įY��}������B� ׿�x�Ϝ�1���*� g�����Ϝ���P��� t�	�ߪ�?���c�u� ߙ�(߽�L߶��߂� ��(�M���q� �� ��6���Z������%� ��I���B�����2�����h����$FoILE_� PR� ���������MDO?NLY 1=.��? 
 ���q ����������~ %�I�m �2��h��!/ �./W/�{/
/�/�/ @/�/d/�/?�//?�/ S?e?�/�??�?<?�? �?r?O�?+O=O�?aO �?�O�O&O�OJO�O�O �O_�O9_�OF_o_
?VISBCKL6>[*.VDv_�_>.PFR:\�_�^�.PVisio�n VD file�_�O4oFo\_joT_ �oo�o�oSo�owo �oB�of�o� +������� +�P��t������9� Ώ]�򏁏��(���L� ^�������5���ܟ k� ���$�6�şZ���~�����
MR_�GRP 1>.�L��C4  B���	 W������*u����RHB ���2 ��� ��� ���B����� Z�l���C���D��������Ŀ��K�wn�J���I�#�T��F�5U�P�Y䲿�ֿ �E�M.G��E$��;n���:G��@O����@���@��[�f @@��_�@�=Y*λ?� F@ ��������J��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<,6\b�π+�&�(�a�L߅�p�A��A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�PS@�P��I'��ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C��������0.��P/ ����/N��/r��/�� �/�??;?&?_?J? \?�?�?�?�?�?�?O �?O7O"O[OFOOjO �O�O�O�O�гߵ��O $_�OH_3_l_W_�_{_ �_�_�_�_�_o�_2o oVohoSo�owo�o�i ��o�o�o��); �o_J�j��� ����%��5�[� F��j�����Ǐ��� ֏�!��E�0�i�{� B/��f/�/�/�/���/ ��/A�\�e�P���t� �������ί��+� �O�:�s�^�p����� Ϳ���ܿ� ��OH� �o�
ϓ�~ϷϢ��� �������5� �Y�D� }�hߍ߳ߞ������� �o�1�C�U�y��� ������������� -��Q�<�u�`����� ����������; &_J\����� �����ڟ�F� j4������� ��!//1/W/B/{/ f/�/�/�/�/�/�/�/ ??A?,?e?,φ?P� q?�?�?�?�?O�?+O OOO:OLO�OpO�O�O �O�O�O�O_'__K_ �o_�_�_�_l��_0_ �_�_�_#o
oGo.oko Voho�o�o�o�o�o�o �oC.gR� v�����	�� �<�`�*<��` �����ޏ��)�� M�8�q�\�������˟ ���ڟ���7�"�[� F�X���|���|?֯�? �����3��W�B�{� f�����ÿ������� ��A�,�e�P�uϛ� b_�����Ϫ_��߀� =�(�a�s�Zߗ�~߻� ��������� �9�$� ]�H��l������ ������#��G�Y� � B�������z������� 
ԏ:�C.gRd ������	� ?*cN�r� ����/̯&/� M/�q/\/�/�/�/�/ �/�/�/?�/7?"?4? m?X?�?|?�?�?�?�? ��O!O3O��WOiO�? �OxO�O�O�O�O�O_ �O/__S_>_P_�_t_ �_�_�_�_�_�_o+o oOo:oso^o�o�op� �o�� ��$�� o�o�~��� ����5� �Y�D� }�h�������׏�� ��
�C�.�/v�<� ��8������П��� �?�*�c�N���r��� �����̯��)��? 9�_�q���JO����� ݿȿ��%�7��[� F��jϣώ��ϲ��� ����!��E�0�i�T� yߟߊ��߮��߮o�o ��o>�t�>�� b�����������+� �O�:�L���p����� ��������'K 6oZ�Z�|�~�� ���5 YD i�z����� �/
//U/@/y/@� �/�/�/�/���/^/? ??Q?8?u?\?�?�? �?�?�?�?�?OO;O &O8OqO\O�O�O�O�O��O�O�O_�O7_���$FNO ����VQ_�
F0fQ kP� FLAG8�(�LRRM_CHKT_YP  WP��^P�WP�{QO=M�P_MIN�P�����P�  �XNPSSB_CF�G ?VU ��_���S� ooIUTP_DEF_OW  ���R&hIRCOM��P8o�$GENO�VRD_DO�V��6�flTHR�V �d�edkd_ENB�Wo k`RAVC_GRP 1@�WCa X"_�o_ 1U<y�r� ����	��-�� =�c�J���n������� �ȏ����;�"�_�pF�X���ibROU�`�FVX�P��&�<b&�8�?���埘�������  D?�јs���@@g�B�7�p�)�ԙ���`SMT�cG��mM���� �LQHoOSTC�R1H����P��at�S5M��f�\���	127.0��=1��  e��ٿ �����ǿ@�R�d��vϙ�0�*�	ano?nymous����0�������/�[��
 � �����r��� �ߨߺ�����-��� &�8�[�I�π��� ����1�C��W� y���`�r������ߺ� ������%�c�u�J \n�������� �M�"4FX�� i������7 //0/B/T/��� m/��/�/�/?? ,?�/P?b?t?�?�/�? ��?�?�?OOe/w/ �/�/�?�O�/�O�O�O �O�O=?_$_6_H_kO Y_�?�_�_�_�_�_'O 9OKO]O__Do�Ohozo �o�o�o�O�o�o�o
 ?o}_Rdv�� �_�_oo!�Uo*� <�N�`�r��o������ ̏ޏ�?Q&�8�J��\���>�ENT 1=I�� P!􏪟  ����՟ğ �������A��M�(� v���^�����㯦�� ʯ+�� �a�$���H� ��l�Ϳ�����ƿ'� �K��o�2�hϥϔ� �ό��ϰ������� F�k�.ߏ�R߳�v��� ���߾���1���U���y�<�QUICCA0��b�t����1������%���2&����u�!ROUTE�Rv�R�d���!P�CJOG����!�192.168�.0.10��w�N�AME !��!?ROBOTp��S_CFG 1H��� ��Auto-sta�rted�tFTP������ � 2D��hz ����U��
/ /./�v���/� ��/�/�/�/�/�!? 3?E?W?i?�/?�?�? �?�?�?�?���AO �?eO�/�O�O�O�O�? �O�O__+_NO�OJ_ s_�_�_�_�_
OO.O oB_'ovOKo]ooo�o P_>o�o�o�o�oo �o5GYk}�_�_ �_��8o��1� C�U�$y�������� ӏf���	��-�?�� ���Ə���ϟ� ����;�M�_�q� ��.�(���˯ݯ�� P�b�t�����m����� ����ǿٿ�����!� 3�E�h��{ύϟϱ� ���$�6�H�J�/�~� S�e�w߉ߛ�jϿ��� �����*߬�=�O�a��s��YT_ERR� J5
���PDUSIZ  ��^J����>��W�RD ?t���  guest}��%�7�I��[�m�$SCDMN�GRP 2Kt;�������V$�K�� 	P01.14 8���   y�����B    �;����� ��������
 �������������~����C�.gR|��� � i  � � 
��������� +��������
���l .Vr���"�l��� m
d�������_GROU��L.�� �	�����07EQUPD � 	պ�J�T�Ya ����TT�P_AUTH 1�M�� <!i?Pendany���6�Y!KAREL:*��
-�KC///A/ �VISION SCETT�/v/�" �/�/�/#�/�/
??�Q?(?:?�?^?p>�C?TRL N�����5�
�FF�F9E3�?�F�RS:DEFAU�LT�<FAN�UC Web S_erver�:
� ����<kO}O�O�O�O��O��WR_CON�FIG O�� ��?��IDL_�CPU_PC@��B��7P�BH�UMIN(\��<TGNR_IO��������PNPT_SI�M_DOmVw[T�PMODNTOL�mV �]_PRTY��X7RTOLNK 1P����_o!o�3oEoWoio�RMAS�TElP��R�O_gCFG�o�iUO�|�o�bCYCLE�o��d@_ASG 19Q����
 ko, >Pbt����������sk�bN�UM����K@�`I�PCH�o��`RTRY_CN@oR���bSCRN����Q���� �b�`�bR���Տ��$J2�3_DSP_EN�	����OBP�ROC�U�iJO�GP1SY@��8�?�!�T�!�}?*�POSRE�~zVKANJI_�` ��o_�� ��T�L�6�͕����CL_L�GP<�_���EYLO�GGIN�`����LANGUA�GE YF7R�D w���LG��U��?⧈�x� ������=P��'0���$ NMC�:\RSCH\0�0\��LN_DISP V��
�ј������OC�R.RD�zVTA{�OGBOOK W
{��i0��ii��X���@��ǿٿ�����"��6	h������e�?�G_BUFF� 1X�]��2 	աϸ��������� ��!�N�E�W߄�{� �ߺ߱�����������J���DCS �Zr� =��� �^�+�ZE��������a�IO 1[
{# ُ!� �!�1� C�U�i�y��������� ������	-AQ cu�������EfPTM  �d �2/ASew� ������// +/=/O/a/s/�/�/��NSEV����TYP�/??y͒�RS@"���>��FL 1\
������?�?�?�?�?��?�?/?TP6���">�NGNAMp�ե�U`�UPS���GI}�𑪅mA_�LOAD�G �%�%DF_M�OTN���O�@MA?XUALRM<��@J��@sA�Q����WS ��@C �]m�-_����MP2�7�^
{ �ر�	�!P�+bʠ�;_/��Rr�W�_�WU�W�_��R 	o�_o?o"ocoNoso �o�o�o�o�o�o�o �o;&Kq\�x �������#� I�4�m�P���|���Ǐ ���֏��!��E�(� i�T�f�����ß��ӟ ���� �A�,�>�w� Z�������ѯ����د ���O�2�s�^��� ����Ϳ���ܿ�'���BD_LDXDI�SAX@	��MEM�O_APR@E ?=�+
 � *� ~ϐϢϴ���������~�@ISC 1_�+ ��IߨT��Q� c�Ϝ߇��ߧ����� w����>�)�b�t�[� ����{�������� ��:���I�[�/���� ��������o�����6 !ZlS��s ����2�A S'�w���� g��.//R/d/��_MSTR `��-w%SCD 1am͠L/�/H/�/�/? �/2??/?h?S?�?w? �?�?�?�?�?
O�?.O ORO=OvOaO�O�O�O �O�O�O�O__<_'_ L_r_]_�_�_�_�_�_ �_o�_�_8o#o\oGo �oko�o�o�o�o�o�o �o"F1jUg �������� �B�-�f�Q���u������ҏh/MKCFG� b�-㏕"L_TARM_��cL�w� σ�Q�N�<�METPU�I�ǂ���)NDSP_CMNTh�p��|�  d�.���ς�ҟܔ|�P�OSCF����PSTOL 1e'�{4@�<#�
5� ́5�E�S�1�S�U�g� ������߯��ӯ��� 	�K�-�?���c�u������|�SING_C�HK  ��;�ODAQ,�f��Ç�~�DEV 	L��	MC:!�HS�IZEh��-��T�ASK %6�%�$1234567�89 �Ϡ��TR�IG 1g�+ l6�%���ǃ�����8�p�YP[� ���EM_INF 1�h3� �`)AT&FVg0E0"ߙ�)���E0V1&A3&�B1&D2&S0�&C1S0=��)�ATZ������H@�����A���AI�@q�,��|���� � ��ߵ�����J���n� �����W��������� ��"����X��/� ���e������ 0�T;x�=� as��/�,/c =/b/�/A/�/�/�/ �/��?���^? p?#/�?�/�?s?}/�? �?O�?6OHO�/lO? 1?C?U?�Oy?�O�O3O  _�?D_�OU_z_a_�_~�ONITOR���G ?5�   	EXEC1Ƀ��R2�X3�X4�X5��X���V7�X8�X9Ƀ�RhBLd�RLd�R Ld�RLd
bLdbLd"b�Ld.bLd:bLdFbLc2�Sh2_h2kh2wh2��h2�h2�h2�h2��h2�h3Sh3_h3��R�R_GRP_�SV 1in���(�����C?BP�P�A4�>%���gY�>r���x�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f���ұ]�l��I��7�������������b��3��´7  ��`�>�����bϸ�z���=�����Jm��
� B�H�˱]����q�	� p� W P�pQ�p��p|  Ъ�g����c�	'� � ���I� � � ����:����
�È=����"�nÿ�	�ВI  �n @B� cΤ�\��ۤ��q��y�o�N���  '������@2�@�����/��C��C�C�@ �C������
��A��* # W @<�P�R�%
h�B�b�A��j������������Dz ۩��߹�����j���( �� -��C���'�7L������Y������ �?�ff ���gy ����o�:a��
�>+�  PƱj�( ����7	���^|�?����xZ��p<
6b<���;܍�<����<� <�&Jσ�AI�ɳ+�|���?fff?I��?&�k�@�.���J<?�` �q�.�˴fɺ�/ ��5/����j/U/�/ y/�/�/�/�/�/?�/0?q��F�?l? ?�?/�?+)�?�?ؿE�� E�I�G+� F��?)O �?9O_OJO�OnO�Of�BL޳B�?_h�.� �O�O��%_�OL_�?m_ �?�__�_�_�_�_�
��h�Îg>���_Co�_goRodo��o�GA�ds�q�C��o�o�o|���ؠ$]Hq���D���pC���pCHmZZ7t���6q�q���ܶN'�3A�A��AR1AO��^?�$�?��K/�±
=ç�>����3�W�
=�#�W��eۣצ�@�����{����<�����(�B�u���=B0������	L���H�F�G����G��H�U�`E���C�+����I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3�l� W���{��������՟ ���2��V�A�z��� w�����ԯ������ ��R�=�v�a����� �������߿��<� '�`�Kτ�oρϺϥ� �������&��J�\� G߀�kߤߏ��߳��� ����"��F�1�j�U� ��y���������� ��0��T�?�Q�����(���3/E�y���u����<��M3�8�����M4Mgs&�IB+2D�a���{�^^	�@�����uP2	P7Q4_A��M00bt��R��`����/   �/�b/P/�/t/�/  *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?��?�?O 2 F;�$�vGb�/�Aa��@�a�`�qC��C�@�o�Ot���KF�� DzH@�� F�P D���O�O�ys<O!_3_E_�W_i_s?���@U@pZ�422�!2~
  p_�_�_�_	oo-o?o Qocouo�o�o�o�o��Q ��+��1���$MSKCF�MAP  �5?� �6�Q��Q"~�cONREL7  
q3��bEXCFENB�?w
s1uXqFNC�_QtJOGOVLKIM?wdIpMrd�bWKEY?w�u�bWRUN�|�u�bSFSPDTY�xavJu3sSIGN?>QtT1MOT�Nq��b_CE_GRoP 1p�5s\r���j�����T�� ⏙������<��`� �U���M���̟��� ���&�ݟJ��C��� 7�������گ��������4�V�`TCOM_CFG 1q}��Vp�����
P�_/ARC_\r
jyUAP_CPL���ntNOCHECK� ?{  	r��1�C�U�g� yϋϝϯ����������	��({NO_WA�IT_L�	uM�NMTX�r{�[m�o_ERRY�2sy3� &��������r�c� ��T_�MO��t��, �~�$�k�3�PAR�AM��u{��	�[���u?�� =�9@345678901��&���E�W� 3�c�����{������������=��UM_RSPAC�E �Vv��$ODRDSP���jx�OFFSET_C�ARTܿ�DIS���PEN_FI�LE� �q��c֮�O�PTION_IO���PWORK kv_�ms �(P(�R�@�6$j.j	 ��Hj(�6$�p=�_DSBL'  �5Js�\���RIENTTO>p9!C��PqfA�� UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?p]a]�D�WcUa쪋l;�	�lmb�`�x7J�`�p����a�< ���`�m�a��H(���H3k7HSM�5G�22G���Gp
��
��c�'|��CR�	>�>q�GsuaT��3���  �4 spBpyr  ]o�*S�B_����j�]��t�q� ��rna �,����6  ��P�Q�|N��M�,k���	'� �� ��I� �  ��%�=��ͭ���ba�	���I  �n @��~���Dp�������N	 W�  '!o�:q�pC	 C�@@sBq�t|��� m�
�!*�h@ߐ�n����*�B	 �A���p�G �-�qbz��P��t�_�������( �� -��恊�n�ڥ[A"]Ѻ�b4�'!5�(p? �?�ff� ��
����OZ�R*��85�z���>΁  	Pia��(5���@����ک�a�c�dF#?��5�x��*�<
6�b<߈;܍��<�ê<� <�&�o&�)��A�lcΐI�*�?f7ff?�?&c����@�.uJ<?�`��Yђ^� nd��]e��[g��Gǡd <����1��U�@�y� dߝ߯ߚ����߼�	� ��-������&��"�E�� E��G+� Fþ����� �������&��J�5��bB��AT�8�ђ ��0�6���>���J� n�7��[m�0���h��1��>��M�I
��@��A�[��C�-�)��?�A��� /�YĒ�a�Jp��vav`CH/�������}!@I��Y�'�3A��A�AR1AO��^?�$�?�����±
=���>����3�?W
=�#����+�e��ܒ������{����<�����.(�B�u���=B0������	��*H�F�G����G��H�U�`E���C�+��-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�?O �?3OOWOBOTO�OxO �O�O�O�O�O�O_/_ _S_>_w_b_�_�_�_ �_�_�_�_oo=o(o aoLo�o�o�o�o�o�o �o�o'$]H �l������ �#��G�2�k�V��� z���ŏ���ԏ��� 1��U�g�R���v��� ��ӟ�������-���(�������y�a����Q�<c�,!3�8�}���,!4Mgs����ɢ�IB+կ篴a���{���A�@/�e�S���w��P!�	P�������7��0ӯ�ϑ�R9�K�`��oχϓϥ�  ���χ����)��M� �����z���{߉ߛ���ߒߤ�������  )�G�q�_����2 F;�$�&Gb���n�a�[ZjM!C�s��@j/�A�S�=�F�� Dz��� F�P D��W����)������������x?���@U@
9�=�=���=��
  v������ �*<N`�*�P ���˨�1���$PARAM�_MENU ?�-�� � DEFP�ULSEl	W�AITTMOUT��RCV� �SHELL_W�RK.$CUR_oSTYL�,�OPT�/PTB�./("C�R_DECSN���,y/�/ �/�/�/�/�/?	??�-?V?Q?c?u?�?�U�SE_PROG �%�%�?�?�3C�CR�����7_HOST !�#!�44O�:T̰�?�PCO)ARC�O�;_�TIME�XB� � �GDEBU�GV@��3GINP?_FLMSK�O�IqT`��O�EPGAPe �L��#[CH�O^�HTYPE����?�?�_�_�_�_�_ oo'o9obo]ooo�o �o�o�o�o�o�o�o :5GY�}�� �������1��Z��EWORD ?}	7]	RS`�_	PNS�$斂JOE!>�TE�s@WVTRACEC�TL 1x-�� �� ������ɆD/T Qy-��䀿D � ��7�4�P  :�L :�GP:�D :�@ :�8�,�>�P�b��� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� V�(�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_d��_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�_���*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p�������� //$)�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �#|"DEF�SPD |�,l!!J �8 IN �TRL }�-�" 8�%�!PE_C�ONFI� ~g%O�g!�$�%��$LID�#�-~74GRP 1�7�Q!�#!A ����&ff"!A+�33D�� D]�� CÀ A@+6�!�" d�$�9�9�*1*0� 	 �+9�(�&�"�? ´	C�?�;B@3AO�?�OIO3OmO"!>�T?�
5�O�O�N��O =��=#�
�O_�O_J_5_ n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_Roxoco�o �o�o�o�o�o�o�>)bM��;
�V7.10bet�a1�$  �A�E�rӻ��A " �p?!G�^�q>���r��0��q�ͻqBQ��qA\�p�q�4�q*�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏� ��4��1�j�U���y� ����֟������0� �T�?�x�c������� ү����!o�,�ۯP� ;�M���q�����ο�� �ݿ�(��L�7�p�x+9��sF@ �� �ͷϥ�g%������ +�!6I�[߆������� �ߠ���������!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ���=(aL ^������ �'9$]�Ϛ��� ��������/<� 5/`�r߄ߖߏ/>�/ �/�/�/�/?�/1?? U?@?R?�?v?�?�?�? �?�?�?O-OOQO<O uO`O�O�O�O�O���O _�O)__M_8_q_\_ n_�_�_�_�_�_�_o �_7oIot���o�o ���o�o�o(/!L/ ^/p/�/{*o��� ������A�,� e�P�b���������� Ώ��+�=�(�a�L� ��p������Oߟ񟠟 � �9�$�]�H���l� ~�����ۯƯ���#� No`oro�on��o�o�o �oԿ���8J\ ng����vϯϚ��� ����	���-��Q�<� u�`�r߫ߖ��ߺ��� ����;�M�8�q�\� ��������z������ %��I�4�m�X���|� ����������:�L� ^���Z�������� ���$�6�H�S wb����� ��//=/(/a/L/ �/p/�/�/�/�/�/? �/'??K?]?H?�?�� �?�?f?�?�?�?O�? 5O OYODO}OhO�O�O �O�O�O�O&8J4_ F_����_�_��_ �_"4-o�O*oco No�oro�o�o�o�o�o �o)M8q\ �������� �7�"�[�m��?���� R�Ǐ���֏�!�� E�0�i�T���x����� ���_$_V_ �2�l_�~_�_�����R�$P�LID_KNOW�_M  �T������SV� ��U͠�U��
��.� ǟR�=�O�����mӣ�M_GRP 1�T�!`0u��T@ٰ)o�ҵ�
���P зj��`���!�J� _�W�i�{ύϟϱ���`������߱�MR��Ņ��T��s�w�  s��ߠ޴߯߅��ߩ� ������A���'�� ����������� ��=���#����������}������S��ST^��1 1��U# ����0�_ A  .��,>Pb�� ������3 (iL^p���(��2*��'�<-/3/)/;/M/4f/x/�/�/�5�/�/�/�/6 ??(?:?7S?e?w?�?8�?�?�?�?~MAD  d�#`PARN_UM  w�\%OSCH?J ME�
�G`A�Iͣ�EUP�D`OrE
a�OT_CMP_��B@�P@�'˥TER_C;HK'U��˪?R�$_6[RSl�¯��_#MOA@�_�U_�_RE�_RES_G � �>�oo8o+o\o Oo�oso�o�o�o�o�o@�o�o�W �\�_ %�Ue Baf�S�  ����S0��� �SR0��#��S�0>� ]�b��S�0}������R�V 1�����rB@�c]��t�(@�c\����D@�c[�$���RTHR_INRl�DA��z˥d,�MASS9�� ZM�MN8�k�M�ON_QUEUE� ���˦��x� URDNPUbQN{�P[��END���_ڙ�EXE�ڕ�@BE��ʟ��OPTIO�Ǘ�[��PROGR�AM %��%�ۏ�O��TASK�_IAD0�OCFG� ���tO��ŠD�ATA���Ϋ@��27�>�P�b�t� ��,�����ɿۿ������#�5�G���INFOUӌ�������� �Ͽ���������+� =�O�a�s߅ߗߩ߻�@�������^�jč�� yġ?PDIT� �ίc���WE�RFL
��
RG�ADJ �n�A	����?����@���?IORITY{�QV}���MPDSPH������Uz����O�TOEy�1�R�� (!AF4�E��P]���!tc�ph���!ud|��!icm���ݏ6�XY_ȡ��R��ۡ)� *0+/ ۠�W :F�j���� ��%7[B��*��PORTT#�BC۠�����_CARTREP�
�R� SKSTA�z��ZSSAV����n�	2500H863���r�$!�U�R����q��n�}/�/�'� URGeE�B��rYWF� #DO{�rUVWV��$��A�WRUP_DELAY �R�>�$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?3A_QSKIP!�n�;l#x 	1/+O + OROdOvO9Hn��O �G�O�O�O�O�O_�O _D_V_h_._�_z_�_ �_�_�_�_
o�_.o@o Roovodo�o�o�o�o �o�o�o*<L�r`���n��$�RCVTM���]��pDCR!�L�ЈqB��C�*J�C$�>��$ >5?-;���04M¹�O���ǃ�������~��9On�Y��<
6b<߈�;܍�>u.��?!<�& {�b�ˏݏ��8���� �,�>�P�b�t����� ����Ο���ݟ�� :�%�7�p�S������ ʯܯ� ��$�6�H� Z�l�~�������ƿ�� �տ���2�D�'�h� zϽ��ϰ��������� 
��.�@�R�d�Oψ� �߅߾ߩ������� ��<�N��r���� ����������&�8� #�\�G�����}����� ������S�4FX j|������ ���0T?x �u����'/ /,/>/P/b/t/�/�/ �/�/�/�/�?�/(? ?L?7?p?�?e?�?�? ��?�? OO$O6OHO ZOlO~O�O�O�?�?�O �O�O�O __D_V_9_ z_�_�?�_�_�_�_�_ 
oo.o@oRodovo�X��qGN_ATC �1�� AT&FV0E/�� ATDP/6/9/2/9�h�ATA�n,�AT%G1%B�960/�++U+�o,�aH,�q�IO_TYPE � �u�sn_�oR�EFPOS1 1}�P{ x�o�Xh_�d_��� ��K�6�o�
���.�ාR����{{2 1�P{���؏V�ԏxz����q3 1���$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����<�>��S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB��-�f��S8 1� ����Y�������y��SMASK 1��P  
9�G��XNOM���a~߈�~�qMOTE  h��~t��_CFG ᢥ����рrPL_�RANG�ћQ��POWER ��e���SM_DRYPRG %i��%��J��TART� �
�X�UME_PRO'�9��~t�_EXEC_EN�B  �e��GS�PD������c��T3DB���RM���MT_!�T����`OBOT_NA_ME i�����iOB_ORD_�NUM ?
��\qH863�  �T���������bPC_TIMoEOUT�� x�`oS232��1��k� LTEA�CH PENDA1N �ǅ�}����`Mainte�nance Co#ns�R}�m
"{�d?KCL/Cg��Z� ��n� ?No Use}�8	��*NPO��Ѯ����(C7H_L��������	�mMAVA#IL��{��ՙ��SPACE1 2��| d��(>��&���p��M,?8�?�ep/ eT/�/�/�/�/�W/ /,/>/�/b/�/v?�? Z?�/�?�9�e�a�=? ?,?>?�?b?�?vO�O�ZO�?�O�O�Os�2�/O*O<O�O`O �O�_�_u_�_�_�_�_[3_#_5_G_Y_o }_�_�o�o�o�o�o[4.o@oRodovo $�o�o����"�	�7�[5K]o� �A����	�̏�?�&�T�[6h�z��� ����^�ԏ���&�� ;�\�C�q�[7���� ����͟{���"�C�@�X�y�`���[8�� ��Ưدꯘ��0�?π`�#�uϖ�}ϫ�[Gw �i� ��:�
G� ���� $�6�H�Z�l�~ߐ��8  ǳ�����߈��d(���M�_�q�� ����������?� ��2�%�7�e�w����� ��������������� !�RE�W����� �����?�Q `�� @ 0��ߖrz	�V_�����
/ L/^/|/2/d/�/�/�/ �/�/�/?�/�/�/*? l?~?�?R?�?�?�?�?@�?�?�?2O�?
���O[_MODE � �˝IS �"��vO,*ϲ��O-_��	M_v_#dCWORK_AD�M���%aR  ���ϰ�P{_�P_?INTVAL�@�����JR_OPTI[ON�V �EBp�VAT_GRP �2����#(y_Ho �e_vo �o�oYo�o�o�o�o�o *<�bOoNDp w������	� ��?�Q�c�u����� /���ϏᏣ����)� ;���_�q��������� O�ɟ���՟7�I� [�m�/�������ǯٯ 믁��!�3���C�i� {���O���ÿտ��� ϡ�/�A�S�e�'ω� �ϭ�oρ������� +�=���a�s߅�Gߕ� �����ߡ���'�9� K�]��߁����y� ���������5�G�Y���E�$SCAN_GTIM�AYuew��R �(�#(�(�<0.a+aPaP
TqA>��Q��oX�����OO�2/��:	d/JaR��WY��^��p�^R^	r  P���� � � 8�P�	�D��GYk} ��������Qp/@/R/x/)P;�o\T���Qpg-�t�_DiKT��[  � lv%��� ���/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OWW �#�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o lO~Od+No`oro�o�o �o�o�o�o�o& 8J\n����8��u�  0�"0g �/�-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q�����$o ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E��� ��Do��������ҿ� ����,�>�P�b�t� �ϘϪϼ���������w
�  58�J�\� n߀ߒߜկ������� ��	��-�?�Q�c�u�p����� �� -����� �2�D�V�@h�z�������������������& ���%	123�45678�" +	��/� ` r������� �(:L^p ������� / /$/6/H/Z/l/~/� �/�/�/�/�/�/? ? 2?D?V?h?�/�?�?�? �?�?�?�?
OO.O@O o?dOvO�O�O�O�O�O �O�O__*_YON_`_ r_�_�_�_�_�_�_�_ ooC_8oJo\ono�o �o�o�o�o�o�oo "4FXj|���������	���s3�E�W�{�C�z  Bp��  � ��2���z��$SCR_GRP� 1�(�U8(�\x^ �@  �	!�	 ׃�� �"�$� ��-��+���R�w����D!~�����#����O����M-10i�A 890990�5 Ŗ5 M61CA >4��Jׁ
� ���0�����#�1�	"�z���О���¯Ҭ � ��c���O�8�J� ������!�����\ֿ��B�y����������A��$�  !@��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ �϶�������%��I� 4�m��<�l߃ߕ��߹�B���\���� 1��U�@�R��v�� ����������;���*<=�
F���?�<d�<�>7�����s@�:��� B����ЗЙ���EL�_DEFAULT�  �����B�MIP�OWERFL  ��$1 WFD�O $��ER�VENT 1������"�pL!�DUM_EIP���8��j!AF�_INE �=�!'FT���9!��4 ��[�!RPC_MAIN\>�J�n'VISw=���o!TP�PU��	d�?/!
PM�ON_PROXY@/�e./�/"Y/��fz/�/!RDMO_SRV�/�	g�/�#?!R C?�h,?o?!
pM�/��i^?�?!RLSgYNC�?8�8�?>O!ROS�.L�4�?SO"wO�#DO VO�O�O�O�O�O_�O 1_�OU__._@_�_d_ v_�_�_�_�_o�_?o�ocoiICE_K�L ?%y (�%SVCPRG�1ho8��e���o�m3��o�o�`4 �`5�(-�`6PU�`7@x}�`���l9��{�d:?��a�o� �a�oE��a�om��a ���aB���aj叟a ���a�5��a�]� �a����a3����a[� ՟�a�����a��%��a ӏM��a��u��a#��� �aK�ů�as���a�� mob�`�o�`8�}�w� ������ɿ���ؿ� ��5�G�2�k�VϏ�z� �Ϟ����������1� �U�@�y�dߝ߯ߚ� �߾�������?�*� Q�u�`������� �����;�&�_�J� ��n������������sj_DEV ~y	�MC:���_OUT�",REC� 1�Z� d �   	�    ��@�� ����A�����
 �PS?D#6 r��UO� �� �� `��� �Z�{� �r� *�  +X�- � I- �- !
- � �X�YZ��PSJ;4 ��?  (� E � ��R ���� E- �� �/e/�l!4�/��� X� (,/>/P/�/�/*�""4� =�!� � ؀  ?"S1h��'!�/���("- ��\?�?$=�= �?�?�?"OOFO4OjO |O^O�O�O�O�O�O�O �O_ __T_B_x_f_ �_�_�_�_�_�_�_o ooPo>oto�oho�o �o�o�o�o�o(
 L:\�p���w,����4� "�X�F�|���p����� ֏ď����0��@� f�T���x�����ҟ� Ɵ���,��<�b�P� ��h�z������ί� �(�:��^�L�n�p� ������ܿ�п� � 6�$�Z�H�jϐ�rϴ� �����������2�D� &�h�Vߌ�z߰ߞ��� ��������
�@�.�d��R��ZjV 1��w P����j� 
�� ��<��
TYPEV�FZN_CFG ;��5d��4�GRP 1��A�c ,B� A�� D;� B����  B4�RB21HE�LL:�(
��?x���<%RS'! ��H3lW� {������`2Vh������%w�����#!�1�����7�2�0d�����HK 1��� �k/f/x/�/�/�/ �/�/�/�/??C?>?�P?b?�?�?�?�?��OMM ����?���FTOV_ENB� ���+�HOW_R�EG_UIO��I_MWAITB�.JKOUT;F��LIwTIM;E���O�VAL[OMC_UN�ITC�F+�MON�_ALIAS ?�e�9 ( he ��_&_8_J_\_B_ �_�_�_�_j_�_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]n��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� ���������ӟ~��� 	��-�?��c�u��� ����V�ϯ����� �;�M�_�q������ ��˿ݿ����%�7� I���m�ϑϣϵ�`� ������ߺ�3�E�W� i�{�&ߟ߱������� ����/�A�S���w� ����X������� ���=�O�a�s���0� ������������' 9K]���� b���#�G Yk}�:��� ���/1/C/U/ / f/�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_O
O�O�O�O �O�OvO�O__%_7_��C�$SMON_�DEFPRO ����`Q� *SY�STEM*  d�=OURECAL�L ?}`Y (� �}xyzr�ate 61=>�inspiron�:4060 ck�\*.*�X507�6 �Q�_�_�_	o � }3copy �frs:orde�rfil.dat� virt:\tmpba�P�]Soeo�wo�o`* bmdb:�P5o�ZKo�o�o i.x d:�Q�l�[@�R�o`r�e/ ua(:�PP��� o*o�o�o_�q����o��o�oL�ݏ���6� �2�empC�192.168.4E�?46:795�_f�px���p �*.d4�@F�O������
�W ����ϟ`�r�����Y;�6 @�R�������tpdisc 0������ѯ�b�t����tpc?onn 0 )�;� M�޿���'���˿ \�nπ�̢���9�K������ ߓ���N�6244����b�t߆�� +�=�O�������)�792����a�s���9 �2�*�<��������0����3���b��t����4 �|=�4� U�����
 }5 �������gy�� +=O���)�6580 ��c u����5�6�� ��"��5�b/t/��/��5�O�1652 W/�/�/�/���/ �)�/`?r?�?�)�;? M?�?�?O'�4�? �?cOuO�O��5/�' �O�O�O/"/�O�(�O b_t_�_����KTV_ �_�_o�_�_>@�_ hozoo�O�O:_�_�o �o
_�oA_�odv ��_.o;�_��� o��Oo`�r����o �o2�oޏ���'�K\�n������$�SNPX_ASG 1�������� P �0 '%R[1]@1.1����?���%֟�� &�	��\�?�f���u� �������ϯ��"�� F�)�;�|�_������� ֿ��˿���B�%� f�I�[Ϝ�Ϧ��ϵ� ������,��6�b�E� ��i�{߼ߟ������� ����L�/�V��e� ������������ 6��+�l�O�v����� ����������2 V9K�o��� ����&R5 vYk����� /��<//F/r/U/ �/y/�/�/�/�/?�/ &?	??\???f?�?u? �?�?�?�?�?�?"OO FO)O;O|O_O�O�O�O �O�O�O_�O_B_%_ f_I_[_�__�_�_�_ �_�_�_,oo6oboEo �oio{o�o�o�o�o�o �oL/V�e �������� 6��+�l�O�v��������PARAM ���� ��	��P�����OFT_KB_?CFG  ⃱����PIN_SIM  ���C�U��g�����RVQST_P_DSB,���������SR ��/�� & CA�R�����TOP_ON_ERސ����PTN� /�@��A	�RING_�PRM� ��V�DT_GRP 1y�ˉ�  	�� ����������Я��� ��*�Q�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߣߠ߲��� ��������0�B�i� f�x���������� ���/�,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZ�~��� ����/ /G/D/ V/h/z/�/�/�/�/�/ �/?
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8___\_��VPRG_COUNT���@���RENB�U��UM�S��__U�PD 1�/�8  
s_�oo*o SoNo`oro�o�o�o�o �o�o�o+&8J sn������ ���"�K�F�X�j� ��������ۏ֏��� #��0�B�k�f�x��� ������ҟ������ C�>�P�b����������ӯί�����UY?SDEBUG�P�P��)�d�YH�SP_�PASS�UB?~Z�LOG ��U+�S)�#�0��  ��Q)�
M�C:\��6���_M�PC���U���Q�ñ8� �Q�SAV �����ǲ%��ηSV;�TE�M_TIME 1]��[ (�P�T�y�ؿT1SVGgUNS�P�U'�U����ASK_OPTION�P�U�Q�Q���BCCFG 3��[u� n�X�G�`a�gZo��߃� ���߹�������:� %�^�p�[����� ���� �����6�!�Z� E�~�i���������%�������&8�� nY�}�?��� � ��(L: p^������ �/ /6/$/F/l/Z/ �/~/�/�/�/�/�/�/ �/2?8 F?X?v?�? �??�?�?�?�?�?O *O<O
O`ONO�OrO�O �O�O�O�O_�O&__ J_8_n_\_~_�_�_�_ �_�_�_o�_ o"o4o joXo�oD?�o�o�o�o �oxo.TBx ��j����� ���,�b�P���t� ����Ώ��ޏ��(� �L�:�p�^������� ʟ��o��6�H� Z�؟~�l�������د ���ʯ ��D�2�h� V�x�z���¿���Կ 
���.��>�d�Rψ� vϬϚ��Ͼ������� *��N��f�xߖߨ� ��8���������8� J�\�*��n����� ��������"��F�4� j�X���|��������� ����0@BT �x�d���� �>,Ntb� �����/�(/ /8/:/L/�/p/�/�/ �/�/�/�/�/$??H? 6?l?Z?�?~?�?�?�? �?�?O�&O8OVOhO zO�?�O�O�O�O�O�O 
__�O@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<o^o�oro�o �o�o�o�o�o  J8n$O���� �X���4�"�X��B�v��$TBCS�G_GRP 2��B�� � �v� 
 ?�  ������׏�� �����1��U�g�z����ƈ�d, ����?v�	 HC{��d�>����~e�CL  B����Пܘ������\)��Y  A��ܟ$�B�g�B�Bl��i�X�ɼ���X��  D	J���r������C����үܬ���D�@v�=�W�j�}� H�Z���ſ���������v�	V�3.00��	mw61c�	*X�0P�u�g�p�>���v�(:�� ��p͟�w  O����p������z�JCFG [�B��� ���������=��=�c�q�K�q� �߂߻ߦ�������� '��$�]�H��l�� �����������#�� G�2�k�V���z����� ���������p* <N���l��� ����#5GY }h����v� b��>�// /V/D/ z/h/�/�/�/�/�/�/ �/?
?@?.?d?R?t? v?�?�?�?�?�?O�? *OO:O`ONO�OrO�O �O��O�O�O_&__ J_8_n_\_�_�_�_�_ �_�_�_�_�_oFo4o jo|o�o�oZo�o�o�o �o�o�oB0fT �x������ �,��P�>�`�b�t� ����Ώ������� &�L��Od�v���2��� ��ȟʟܟ� �6�$� Z�l�~���N�����د Ư�� �2��B�h� V���z�����Կ¿� ���.��R�@�v�d� �ψϪ��Ͼ������ �<�*�L�N�`ߖ߄� �ߨ����ߚ����� ��\�J��n���� �������"���2�X� F�|�j����������� ����.TBx f������� >,bP�t �����/�(/ /8/:/L/�/�ߚ/�/ �/h/�/�/�/$??H? 6?l?Z?�?�?�?�?�? �?�?O�?ODOVOhO "O4O�O�O�O�O�O�O 
_�O_@_._d_R_�_ v_�_�_�_�_�_o�_ *ooNo<oro`o�o�o �o�o�o�o�o&�/ >P�/���� �����4�F�X� �(���|�����֏� ���Ə0��@�B�T� ��x�����ҟ����� �,��P�>�t�b��� ������������ :�(�^�L�n������� 2d�����̿�$� Z�H�~�lϢϐ����� ���Ϻ� ��0�2�D� zߌߞ߰�j������� ���
�,�.�@�v�d� ������������ �<�*�`�N���r��� ����������& J\�t��B� �����F4 j|��^���8�/�  2 6#� 6&J/6"�$�TBJOP_GR�P 2����  ?��X,i#�p,� ��xJ� �6$�  �<� �� �6$� @2 �"	 ��C�� �&b  �Cق'�!�!>��1�
559>�0+1��33=�C�L� fff?+0?�ffB� J1�%Y?�d7�.��/>���2\)?0�5����;��hCY�� �  @� �!B�  A�P?�?�3~EC�  D�!8�,�0*BOߦ?�3�JB��
:���Bl�0��0�$�1�?�O6!Aə�A�̔C�1D�G6�=qq�E6O0�p��B��Q�;�A}�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH�1�ts�A@33@?1� C�� �@�_x�_&_8_>��D�U�V_0�LP�Q30<{�zR� @�0�V�P !o3o�_<oRifoPo^o �o�o�oRo�o�o�o�o M(�ol�p~(��p4�6&�q5	V3.00�#�m61c�$*�(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�Na�F���F�^l�F���F�:
�F�)F��3�G�G���G��G,I�R�CH`�C�d�TDU�?D���D��DE(!�/E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[�
F���F��{M;S@;Q��|8�`rz@/&�8�6&<��1�w�^$�ESTPARS c *({ _#HR��ABLE 1�p+IZ�6#|�Q� � 1�|�|�|�5'=!*|�	|�
|�|�˕�6!|�|�|�N��RDI��z!ʟ@ܟ� ��$���O�������¯ԯ�����S��x# V���˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� U-����ĜP�9�K�]� o��-�?�Q�c�u���~6�NUM  ��z!� >  �Ȑ����_CFG ������!@b IMEBF_TT��p��x#��a�VER���b�w�a�R 1Ξp+
 (3�6"1 ��  6!������ ���� �9�$�:�H�Z� l�~����������������^$��_��@�x�
b MI_CH�ANm� x� kDOBGLV;0o�x��a!n ETHERA�D ?�� ��y�$"�\&n R�OUT��!p*!�*�SNMA�SK�x#�25�5.h�fx^$O�OLOFS_DI�[ՠ	ORQC?TRL �p+;/ ���/+/=/O/a/ s/�/�/�/�/�/��/��/�/!?��PE_D�ETAI��PON_SVOFF��33P_MON ��H�v�2-9STRTCHK ����42VTCOM�PATa8�24:0FPROG %��%CA)&O�3I�SPLAY��L:_�INST_MP 2GL7YDUS���?��2LCK�LPKQUICKMEt �O�2oSCRE�@�
tps��2�A�@�I��@_Y���9��	SR_GRP �1�� ���\�l_zZg_�_�_�_�_�_�^�^�oj �Q'ODo/ohoSe��o o�o�o�o�o�o�o !WE{i�������	1234567��!�ڎ�X�E1�V[
 ��}ipnl/�a�gen.htm�no��������ȏ~��Panel s/etup̌}�?�`�0�B�T�f� �� 񏞟��ԟ���o� ���@�R�d�v����� �#�Я�����*� ��ϯůr��������� ̿C��g��&�8�J� \�n�����϶����� ����uϣϙ�F�X�j� |ߎߠ����;��������0�B��*NUA�LRMb@G ?�� [������ ������ ��%�C�I��z�m�������v�SEoV  �����t�ECFG �Ё=]/BaA$  w B�/D
 �� /C�Wi{��� ���� PRց; �To\o�eI�6?K0(%�� ��0�����/ /;/&/L/q/\/�/�/�/l�D �Q�/�I_�@HIST �1ׁ9  (�  ��(/S�OFTPART/�GENLINK?�current=�menupage?,153,1?v?8�?�?�?�� >?P=962c?�?
OO.O�?�?�136�?|O�O �O�OAOSOeO�O__ 0_�HM___q_�_�_�_ �_H_�_�_oo%o7o �_[omoo�o�o�oDo �o�o�o!3E ��a81�ou��� ���o���)�;� M��q���������ˏ Z�l���%�7�I�[� ��������ǟٟh� ���!�3�E�W���� ������ïկ�v�� �/�A�S�e�Pb�� ����ѿ������+� =�O�a�s�ϗϩϻ� ������ߒ�'�9�K� ]�o߁�ߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y��� v�����������	 �?Qcu��( ����)� M_q���6� ��//%/�I/[/ m//�/�/�/D/�/�/ �/?!?3?�/W?i?{? �?�?�?�����?�?O O/OAOD?eOwO�O�O �O�ONO`O�O__+_ =_O_�Os_�_�_�_�_ �_\_�_oo'o9oKo �_�_�o�o�o�o�o�o jo�o#5GY�o�}������?���$UI_PAN�EDATA 1������  	�}��0�B�T�f�x��� ) ����mt�ۏ���� #�5���Y�@�}���v� ����ן�������1���U�g�N������ �1��Ïȯگ� ���"�u�F���X�|� ������Ŀֿ=���� ��0�T�;�x�_Ϝ� �ϕ��Ϲ������,���M��j�o߁ߓ� �߷������`��#� 5�G�Y�k��ߏ��� �����������C� *�g�y�`��������� F�X�	-?Qc ����߫���� ~;"_F� �|�����/ �7/I/0/m/�����/ �/�/�/�/�/P/!?3? �W?i?{?�?�?�?? �?�?�?O�?/OOSO eOLO�OpO�O�O�O�O �O_z/�/J?O_a_s_ �_�_�_�O�_@?�_o o'o9oKo�_oo�oho �o�o�o�o�o�o�o# 
GY@}d�� &_8_����1�C� �g��_��������ӏ ���^���?�&�c� u�\�������ϟ��� ڟ�)��M����� ������˯ݯ0��� ��7�I�[�m������ ����ٿ�ҿ���3� E�,�i�Pύϟφ���0����Z�l�}���1� C�U�g�yߋ�)߰� #������� ��$�6� ��Z�A�~�e�w��� ��������2��V��h�O�����v�p��$�UI_PANEL�INK 1�v��  ��  ��}12�34567890 ����	-?G � ��o�����a ��#5G�	�����p&���   R�����Z� �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?.O@O ROdOvO�O O�O�O�O �O�O_�O�O<_N_`_0r_�_�_�0,���_ �X�_�_�_ o2ooVo hoKo�ooo�o�o�o�o �o�o��,>r} ��������� ���/�A�S�e�w� �������я���t v�z����=�O�a� s�������0S��ӟ� ��	��-���Q�c�u� ������:�ϯ��� �)���M�_�q����� ����H�ݿ���%� 7�ƿ[�m�ϑϣϵ� D��������!�3�E� �_i�{�
�߂����� �������/��S�e� H���~��R~'�'� a��:�L�^�p��� ������������  ��6HZl~�� �#�5��� 2 D��hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?�/ �?�?�?�?�?�?m?O O&O8OJO\O�?�O�O �O�O�O�O�O[�_�� 4_F_)_j_|___�_�_ �_�_�_�_o�_0oo Tofo��o��o��o �o�o,>1b t����K�� ��(�:����{O ������ʏ܏�uO� $�6�H�Z�l������� ��Ɵ؟����� �2� D�V�h�z�	�����¯ ԯ������.�@�R� d�v��������п� ��ϕ�*�<�N�`�r� ���O�Ϻ�Io������ ���8�J�-�n߀�c� �߇����߽����o 1�oX��o|���� ���������0�B� T�f������������ ��S�e�w�,>Pb t��'���� �:L^p� �#���� // $/�H/Z/l/~/�/�/ 1/�/�/�/�/? ?�/ D?V?h?z?�?�?�??? �?�?�?
OO.O��RO dO�߈OkO�O�O�O�O �O�O_�O<_N_1_r_ �_g_�_7OM�m��$UI_QUI�CKMEN  >��_Ao�bRESTORE� 1�?  �|��Rto�o�im�o�o�o�o �o:L^p� %������o� ���Z�l�~����� E�Ə؏���� �Ï D�V�h�z���7����� ��/���
��.�@�� d�v�������O�Я� ����ßͯ7�I��� m�������̿޿��� �&�8�J��nπϒ� �϶�a�������Y�"� 4�F�X�j�ߎߠ߲� �����ߋ���0�B�T�gSCRE`?�#mu1s]co`u2��3��U4��5��6��7��y8��bUSERq�dv��Tp���ks����4��5��6��7���8��`NDO_�CFG �#k � n` `PDA�TE ����NonebSE�UFRAME  ��TA�n�RTO?L_ABRTy�l�Α�ENB����GR�P 1�ci/aCz  A�����Q@�� $6HR�d��`U�����MSK  �����MNv�%�U�%����bVISCAN�D_MAX�I���FAIL_�IMG� �PݗP#���IMREGN�UM�
,[SI�Z�n`�A�,~VONTMOU��@���2���a��a��~��FR:\� � MC{:\�\LOG�7B@F� !�'/�!+/O/�Uz �MCV�8#U�D1r&EX{+�S|�PPO64_���0'fn6PO��LIb�*�#9V���,f@�'�/�� =	�(SZV��.����'WAI��/STAT 	����P@/�?�?�:�$�?�?��2DW�P  ��P yG@+b=��� H��O_JMPE�RR 1�#k
 � �2345678901dF�ψO{O �O�O�O�O�O_�O*_�_N_A_S_�_
� M�LOWc>
 �_�TI�=�'M�PHASE  ���F��PSHI[FT�1 9�]@<�\�Do�U#oIo �oYoko�o�o�o�o�o �o�o6lCU �y����� �@�	�V�-�e2����	VSFT1�2�	VM�� ��5�1G� ���%A_�  B8̀̀E�@ pكӁ˂�у���z�ME@�?��{��!c>&%�aM�1��k�0�{ �$�`0TDINEND��\�O� �z���S��w��P��=�ϜRELE�Q���Y���\�_ACT�IV��:�R�A ���e���e�:�R�D� ���YBOX� �9�د�6���02���1�90.0.�83v��254�:�QF�	 �X��j��1�ro�bot���  � p�૿�5pc��̿������7�����-�f�ZABC�����,]@U��2 ʿ�eϢωϛϭϿ� ���� ���V�=�zߐa�s߰�E�Z��1� Ѧ