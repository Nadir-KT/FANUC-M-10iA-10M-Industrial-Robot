��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ����ALRM_�RECOV1   $ALMO�ENB��]ON�i�APCOUPwLED1 $[�PP_PROCE�S0  �1��FPCUREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYO12 � u3|�4|GRG_ST�R1 � $�TITP$I��1�{���T��5�6�7�8�9�0��z������1�1��1 '1
'2"(��ASBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�H UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2F�G1_�3�B�2G�XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�Al{G BL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa4 hq;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S~�BSS�CHG,]I1 [ Tp4�"3I9�TY�D,P*2 �`w@� �!,R*HD�cJ* C���2��3��4��5���6��7��8��9�4!� CO�$ <� $6xK3 1w`�O_M�@�C t� � E#6NGP�ABA� �c��ZQ ���`���@nr��� ��P�0���p� �v�p�PzPb26h����"J�_R���BC�J��3�JVP��tBS��}Aw���"�tP_*0OFS�zR @� RO_�K8���aIT�3��N'OM_�0�1ĥ3q���T �� �$���AxP��K}EX �� �0g0I01��p��
$TFa��C$M�D3��TO�3�0U�� �� �H�w2�C1|�EΡg0�wE{vF�vF�40C�Pp@�a2 
P$�A`PU�3N1)#�dR*�AX�!sD�ETAI�3BUFpV��p@1 |�p�۶�pPIdT� PP[�MZ�Mg�Ͱj�}F[�SIMQSI �"0��A.���F��lw' Tp|zM��P��B�FACTrbHPEW7�P1Ӡ��vv��MCd� ��$*1JB�p<�*1D#ECHښ�H���b�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF���� &k�Bv�u�cu��a E�� !2��+�MQ��EчSIZ�3����T��P�����aRSINF�����kq��������LX������F�CRCMu�3CC lpG��p���O}���b��1�������2�V�D
xIC��C���r����0P��{� EV �zUF_��F�pNB
0�?������A�! �r�Rx���� V�lp�2��aR�t�,��gp�RTx �#�5�5"2��uARt���`CX�$LG�p��B�1 `s�P�t�a!A�0{�У+0R���tME�`!BupCr3RA 3tAZ�л4�pc�OT�FC�b�`��`FNp���1��ADI+�a%��b��{��p$�pSp�c�`S0�P��a,QMP6�`IY�3��M'�pU���aU  $m@TITO1�S�S�!���$�"0�DBPXW�O��!��$S1K��2��DB��"�"@�PR8� �
� ���# lm@q1$��$��
+�L9$?(�V�)%@?R4C&_?�A����PE��'�~?(�� RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@4a��C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!��DCS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�o CdSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc �@Sp�i�a+ �j�f�"��pOGIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�� 6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6dr�!MSW�U. 8��KEYI��5�TM�1�s�qoA�vINޱE��!, �/ D��HOST�P!4���<���`<�°<��p<�EM'����Z�R��pL� U}L��0  �	8����DT�0?1 � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0�QS�����#��SAV �����c�S< 9�`��fP$�0E!� YwN_B�#2 0��DI�d�pO|�m��#�$F�R_IC�� �ENC2_Sd3  ��< 3����� cgp����B4�"��2�A��ޖ5���`ǻ��@Q@K&D-!�a�A�VER�q����D3SP
���PC_�q���"�|�ܣ�VALMU3�HE�(�M�sIP)���OPPm �TH�*���S" T�/�Fb�;�dp����d D�(��{ET6 H(rLL_DUǀ�a�@`��k���֠OT�"�U�/��o�@@NOA�UTO70�$�}�x�~�@s��|�CJ� ��C� �ia�z�L�� 8H *��L� ���Բ @sv��`� �� ÿ��� Xq��cq���q���q��U7��8��9��0����1�1 �1-�1�:�1G�1T�1a�1Jn�2|�2��2 �U2-�2:�2G�2T�U2a�2n�3|�3ʩ3� �3-�3:�3�G�3T�3a�3n�4�|�2w�����9 A<���z�ΓKI��0��H硵BaFEq@{@�: ,��&a?3 P_P?��>�
����E�@��iaQQ���;fp$TP~�$VARI��ܮ�,�UP2Q`< W�߃TD��g���`�������!��BAC��"= T2����$)�,+r³�p IFI@��p�� q M�P"��l@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� FW�@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(��a�#5T�DG���� �%��FSS� )�?C P(q1�1�`Q_1"811�EC�13D;5D6�GR)A���@�����P�W�ON2EBUG�S�2�C`gϐ_E A ���?����TERuM�5B�9ORIw�0C�5r��SM_h-`���0D�9TA�9�E�7 �UP��F�� -QϒA��P�3�@B$SEG�GJ� EL�UUSE.PNFI��pBx���1@��4>DC$UF�P��$���Q�@"C���G�0T������SNSTj�PATxۡg��APTHJ�A�E*�Z%qB\`F�{E��F�q�pARxPY�aSHFT͢qA�AX_SHOR$�>��6% @$GqPE���GOVR���aZPI@P�@$U?r *aAYLO���j�I�"d��A8ؠ��ؠERV��Q i�[Y)��G�@R��i�e��i�R�!P�uA�SYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C��%UP���P���WORڒ@M��k0SM5T��G��GR��3�aPA�@��p5�'�_H � j�A�'TOCjA7pP]Pp$OPd�O��C��%�p�O!��R%E.pR�C�AO�?��Be5pR�EruIx|'QG�e$PWR) 3IMdu�RR_$s��\5��B Iz2H8��=�_ADDRH�H_LENG�B�q�qT:�x�R��So�J.�SS��SK�����0� ��-�SE*��m@HSN�MN1K	�j�5�@r�֣OL��\�WpW�Q�>pACRO�p���@�H ����Q� ��OSUPW3�b_>�I��!q�a1�������� |��������-���X:���iIOX2S=��D�e��]���L� $��p�!_OFyF��_�PRM_�{�aTTP_��H��M (�pOB�J�"�pG�$H�L�E�C��ٰN �s 9�*�AB_��T��
�S�`�S��L�V��KRW"duHIoTCOU?BGi�LO�q����d�0 Fpk�GpSS� ��G�HWh�wA��O.�}�`INCPUX2VISIO��!���¢.�á<�á-� ��IOLN)�P 8�7�R'���$SLz�bd PUT_��$dp�Pz ��^� F_AS2Q/�$LD���D�aQT U�0]P�A������PHYG灱Z�̱5�sUO� 3R `F� ��H�Yq�Yx�ɱvpP�Sdp���x��ٶ�%�UJ��S����N�E�WJOG�G �DIS��&�KĠ��3T |��AV��`_��CTR1S^�FLA�Gf2@LG�dU ��n�:��3LG_SIZ��ň��,=���FD��I���� Z �ǳ��0�Ʋ�@s�� -ֈ�-�=�-���-��0<-�ISCH_��DqR��N?���V��EAE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�BOO>)�WL ?`�� �ITV���0\�REC�SCRf 0�a��D^�����MARG ��`!P�)�T�/ty�?I�S�H�WW�I����T�JGM��MNC�H��I�FNKEY���K��PRG��UqF��P��FWD��HL�STP��V`��@�����RSS�H�` �Q�C�T1�ZbT�R ���U����� |R��t�i���G��8PCPO��6�F�1�M���FOCU��RGE]XP�TUI��I���c��n��n�� ��ePf���!p6�eP7�9N���CANAI�jB޾�VAIL��CL�t!;eDCS_HI�4�.��O�|!�S Sn瘱^I�BUFF1XY�5�PT�$�� ��v��f�L6q1Y�Y��P �����pO+S1�2�3����_�0Z � � ��aiE�*��ID%X�dP�RhrO�+��A&ST��R��Y�z�<! Y$EK&CK+���Z&m&KF�1[ L��o�0 ��]PL�6pwq�t^�����w��7�_ \ �`��瀰�7��#�0�C��] ��CL�DP��;eTRQL�I�jd.�094FLAGz�0r1R3�DM��R7��LDR5<4R5ORG.���e2(`���V��8.��T<�4�d^ A�q�<4��-4R5S�`�T00m��0DFRCLMC!D�?�?3I�@��MIC��d_ Yd���RQm�q��DSTB	�  ؏Fg�HAX;b |�H�LEXCESZr��rBMup�a`�p@�B;d��rB`��`a��F_A�J��$[�Ot�H0K�db \���ӂS�$MB��LI�Б}SREQUIR��R>q�\Á�XDEB�U��oAL� MP�c@�ba��P؃ӂ!BoA#ND���`�`d�҆��c�cDC1��IN@�����`@�(h?Nz��@q��o�PT�SP�ST8� e�rL�OC�RI�p�E�X�fA�p��AoAOwDAQP�f X��3ON��(2MF���� �f)�"I��%�e��T�v��FX�@IGG� g �q��"E��0��#���$R�a% ;#7y��Gx��VvCPi�ODATAw�pE:��y��RFЭ�NVh �t $MD�qI�ё)�v+�tń�tH��`�P�u�|��sAN�SW}��t�?�uD��)�b�	@Ði -�@CU��V�T0�eRR2�j D�ɐ�Qނ�Bd$CA�LI�@F�G�s�2��RIN��v�<?$�INTE����kE���,��b����_Nl��ڂ��kDׄ�Rm�DIViFD�H�@ـn�$�V��'c!$���$Z�����~��[��oH �$�BELTb��!ACCEL+��ҡ���IRC�t����T</!��$PS�@#2L  �Ė83����x��� ��PATH���������3̒Vp�A_@�Q�.�4�B�C�_MGh�$D�DQ���G�$FW�h��p��m�����b�D}E��PPABNԗROTSPEED����00J�Я8��@���̐$USE_d��P��s�SY���c�A kqYNu@A�g��OFF�q�M�OUN�NGg�K�O9L�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I̒��4��\BݠVEO�w�Ͳ2�3_UPE�߳LOWL���00����D���BwP��� ��1RCʀƶMOSI�V�JRMO���@GP�ERCH  �OV��^��i�<!� ZD<!�c��d@�P��BV1�#P͑��L�0��EW��ĸUP��Ŝ���TRKr�"AYLOA'a�� Q-��̒<�1Ӣ`0 ��RT1I$Qx�0 MO���Ѐ�B R�0J��D��s��H����b�DUM2�(�S_BCKLSH_C̒��>�=�q� #�U��ԑ���2�t�]ACLALvŲ�1nМP�CHK00'%SD�RTY4�k��y�1�q_6#2�_UM�$Pj�Cw�_�SCL���ƠLMT_J1_LO��@���q��E�����๕�幘SPC��7������PCo���H� �PU�2m�C/@�"XT_�c�CN_��N��e���SFu���V�&#�� ��9�̒��=�C�u�SH6#��c����1�р��o�0�͑
��_�P�At�h�_Ps�W�_ 10��4�R�01D�VG��J� L�@J�OG|W���TORQU��ON*�Mٙ�sRH�L���_W��-�_=���C��I��I�IJ�II�F�`�JLAX.�1[�VC��0�D�BO1U�@i�B\�JRKU��	@D�BL_SMd�BM�%`_DLC�BGR�V��C��I��H�_� �*COS+\�(LN�7+X >$C�9)I�9)u*c,�)�Z2 HƺMY�@!�( "TH&-�)T�HET0�NK2a3I��"=�A CB6CB=�C�A�B(2061C�616SBC�T2N5GTS QơC� �aS$" �4c#�7r#$DUD�EX�1s� t��B�6���AQ|r�f'$NE�DpIB U�H\B5��$!��!A�%�E(G%(!LPH$U�2׵�2SXpCc% pCr%�2�&�C�J�&!�EVAHV6H3�YLVhJUVuKV�KV�KV�KV�KV�IHAHZF`RPXM��wXuKH�KH�KUH�KH�KH�IO2L�OAHO�YWNOhJO�uKO�KO�KO�KO
�KO�&F�2#1ic%��d4GSPBALA�NCE_�!�cLE6k0H_�%SP��T&��bc&�br&PFUL�C�hr�grr%Ċ1=ky�UTO_?�j�T1T2Cy��2N &�v�ϰctw�g�p�0(Ӓ~���T��O���>� INSEGv�!��REV�v!���DI�F��1l�w�1m
�OB�q
�����MIϰ1��LCHgWAR��
�AB&~u�$MECH,1�� :�@�U�AX:�P���Y�G$�8pn 
pZ��|���ROBR��CR̒��N�(��MSK_�`f�p� P Np_��R ����΄ݡ�1��Ұ�Т΀ϳ��΀"�IN��q�MTCOM�_C@j�q  �L��p��$NO�RE³5���$�7r 8� GR�E��SD�0ABF�$?XYZ_DA5A���DEBU�qI���Q�s �`$�COD�� ��k�F��f�$BUFIwNDXР  ���MOR��t $-�U��)��r�B������Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��E����E3 �OPsWO�ŀv0���SYSBU�@ʐ$�SOP����#�U<"��pPRUN�I�PA�DH�D����_OU�=��qn�{$}�IMAG��iˀ�0P�qIM��Ơ�IN�q���RGOVRDȡ:���|�aP~���Р�0L_6p0���i��RB���0e��M���EDѐ*F� ��N`M*���o�'�˱SL�`�ŀw x $OwVSL�vSDI��DEXm�g�e�9w�$����V� ~�N���@w����Ûǖȳ�M��͐�q<��� �x HˁE�F�AT+US���C�0à�ǒ��BTM����I
f���4����(�ŀy DˀEz�g���PE�r�����
���EXE��V��E�Y�8$Ժ ŀz @ˁ��3UP{�h�$�p��XN���9�H�� �PG"�{ h? $SUB��c��@_��01\�MPW�AI��P����LO��<�F�p�$R�CVFAIL_C�f�BWD"�F����DEFSPup | Lˀ`�D�� U�UNI��S�b��R`���_L�pAP��̐���ā}���� B�~���|��`ҲNN�`KET��y���P� $�~���0SIZE��ଠ{����S<�OR��FORMAT/p � F��ᖫrEMR��y�UqX���@�PLI7�~ā  $�P_SWI��Ş�_PL7�AL_ S�ސR�A��B��(0C��Df�$E�h����C_=�U�� � � ���~�J3�0�����TIA4��5��6��MOM������h �B�AD��*��* PU70NARW��W ���V����� A$PI�6���	�� )�4l�}69��Q�|��c�SPEED�PGq�7�D�>D�� ���>tMt[��SAM�`痰>��MOV���$�@�p�5��5�D�1�$2�������{�2��Hip�IN?,{� �F(b+=$�H*�(_$<�+�+GAMM�f�1>{�$GET��Đ�H�D����
^pLI�BR�ѝI��$H�I��_��Ȑ*B6Eď�*8A$>G086LW =e6\<G9�686��R���ٰV��$�PDCK�Q�H�_����;"��z�.%��7�4*�9� ��$IM_SR�O�D�s"���H�"�L	E�O�0\H��6@�� �ŀ�P~�qUR_SCR����AZ��S_SAV�E_D�E��NO��CgA�Ҷ��@�$�� ��I��	�I� %Z[ � ��RX" ��m�� �"�q�'"�8� Hӱt�W�UpS���*�M��O㵐.' }q��Cg���@ʣ����тM�AÂ� �� $PY��3$WH`'�NGp��� H`��Fb��Fb��Fb��PLM���	� 0h�H�J{�X��O��z�Z�e8T�M���� pS��C��O__0_B_t�a��_%�� |S� ���@	�v��v �@���w�v��EM��%��es�B�ː��ftPn��PM��QU� �U�Q��Af�wQTH=�HOL��oQHYS�ES�F,�UE��B��O#��  -�P0�|�gAPQ���ʠu���O��ŀ�ɂv�-�A;ӝGROG��a2D��E�Âv�_�ĀZ�INFO&��+����b�Ȝ�OI킍 ((@SLEQ/�#@������o���S`�c0O�0�01E�Z0NUe�_�AUT<�Ab�COPY���(��{��@M��N������1�P�
� ��RG4I�����X_�Pl�C$�����`�W���P��j@�G���E�XT_CYCtb����p����h�_NA�!$�\�<��RO�`]�� �s m��POR�㸅����SRVt�)l����DI �T_l� ��Ѥ{�ۧ��ۧ �ۧU5٩6٩7٩8��Ҝ�S�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,(@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#q��QSwKIP�� ĕ�Zx�O�`NT!� ��P_x���ǚ@�b �p1�1�1Ǹ�?�  �?��>��>�&�>��3�>�9�J2R�;쐖 4��EX� TQ����ށ�Q����[�KFд�w�RD�CIf� �U`�X}�R�#%M!*�0�)�~�$RGEAR_0sIO�TJBFLG�L�igpERa��TC݃�������2TH2N<��� 1�b��uGq T�0 ����M���`Ib�����REF�1�� yl�h��ENAB��lcTPE?@���! (ᭀ����Q�#�~��+2 H�W���2�Қ����"�4�F�X�j�3�қ{��������
j�4�Ҝ��
��.�P@�R�����5�ҝu�@����������j�6�����(:Lj�7�ҟo�����j�8�Ҡ���"4Fj�SMSKJ�����a��E�A���MOTE�������@ "1��Q�IIO�5"%I��tRd�9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C��>%/S232%�Sb�i�DEVICEUS�#�R�RPARIT|�!OPBIT�Q���OWCONT�R��Qⱓ�RCU�� M�SUXTAS�K�3NB��0�$TATU�P�P� @@R쐦F�6�_�PC}��$FREEFR�OMS]p�ai�GE�TN@S�UPDl�A6RB�'��SP%0��ߧ� !m$USA���az9�L��ERI�0���pRY$�5~"_�@��P�1�!N�6WRK��D9��F9ХFRIEND�Q4bUF��&�A@oTOOLHFMY5��$LENGTHw_VT��FIR�p�qC�@�E� IUF�IN�R���RGyI�1�AITI:�bxGX��I�FG2�7�G1a����3�B�GP1RR�DA��O_� o0e�I1RER�đ�3&����TC���AQJV ��G|�.2���F� �1�!d�9Z�8+5K�+5౑E�y�L0�4�XS �0m�LN�T�3�Hz��89��%�4�3G���W�0�W�RdD �Z��Tܳ��K�a3d���$cV 2����1��I1H�02*K2sk3K3Jci �aI�i�a�L��SL���R$Vؠ�BV�EVPk�]V*R��� �,6 Lc���9V2F{/P:Bֵ�PS_�Et�$prr�C�ѳ$A0���wPR���v�U�cS�k�� {����3���# 0���VX`�!�t�X`��0P�Ё�
z�uSK!� �-q�R��!0���z�N�J AX�!h�A�@LxlA��A�THIC�1��������1TFE����q>�IF_CH��3A�I0�����G�1�x������9�nɆ_JF҇PR(����RVAT�� �-p��7@����sDO�E��COU(���AXIg��OF�FSE+�TRIG �SK��c���Ѽ�e�[��K�Hk���8�IGM�Ao0�A-��ҙ�ORG_UNEV�Ξ� �S�쐮Od �$�������GROU��ݓTO�2��!ݓDSP��JcOG'��#	�_P'��2OR���>P6KEPl�IR�0�P�M�RQ�AP�Q��Ep�0q�e���SYSG���"��PG��BRK *Rd�r�3�-�������ߒ<pAD��ݓJ�OBSOC� N�DUMMY14�p�\@SV�PDE_O�P3SFSPD_WOVR��ٰCO�L�"�OR-��N�0b.�Fr�.��OV�CSFc�2�f��F���!4�S��RA�"LC�HDL�RECOQV��0�W�@M��յ�RO3��_��0� @�ҹ@V�ERE�$OFSf�@CV� 0BWDG��ѴC��2j�
�TR��!��E_FD}Oj�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��2_�Gxǋ�AM��k�0J0������_M��2x{�#�8$CA��{Й���8$HBKX|1c��IO��.�:!aPPA"�N�3��^�F���:"�DVC_DB�C��d�w"�Ј��!��1���ç�3�����ATIO� ��q0�UC�&CAB�BS�PⳍPȲȖ��_0c�SUOBCPUq��S�P a aá�}0�Sb��c���r"ơ$HW_C ���:c��IcA�A-��l$UNIT��l���ATN�f����C�YCLųNECA���[�FLTR_2_FI���(��}&���LP&�����_SC-T@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb�r�v: _T��PRO��,O�� EM�_��98u�q u�q���DI�0e�RAI�LAC��}RMƐL!OԠdC��:anq��Xwq����PR��SLQI�pfC��30	���FUNCŢ�rRI�NkP+a�0 ��!RA� >R 
Я��ԯWAR�BLFQ��A�����DA�����LDm0�aB9��nqBTIvrbؑ����PRIAQ1�"AFS�P�!����P�`%b���M�I1U�DF_j@��y1°�LME�FA�@HR�DY�4��Pn@RS�@Q�0"�MULS�Ej@f�b�q ��X��ȑ���$�.A$�1$c1�Ó���� x�~�EG� ݓ�q!A1R����09>B�%���AXE��RO%B��W�A4�_�-֣CSY���!6��&S�'�WR���-1���SCTR��5�9�E�� 	5B��=QB�90�@6������OT��0o 	$�ARAY8�w20���	%��FI��;�$LI�NK�H��1�a_�63�5�q�2XYZ"��;�q�3@��1)�2�8{0B�{�D��� CFI���6G��
�{�_�J��6��3aOP�_O4Y;5�QTB�mA"�BC
�z�DU�"�66CTURN 3�vr�E�1�9�ҍGFL�`���~ �@�5�<:7�� 1�J?0K�Mc�68Cpb�vrb�4�ORQ�� X�>8�#op�������wq�Uf�����TOV	E�Q��M;�E#�UK#�UQ"�VW�ZQ�W ���Tυ� ;����Q H�!`�ҽ��U�Q�Wke0K#kecXER���	GE	0��S�dA WaǢ:D���7!�!AX�rB!{q�� �1uy-!y�pz �@z�@z6Pz\Pz � z1v�y�y �+y�;y�Ky�[y �ky�{y��y�q�yoDEBU��$� ���L�!º2WG`  CAB!�,��SV���� 
w���m��� w����1���1���A�� �A��6Q��\Q���!�pm@��2CLAB3B��U�����S � ÐER���� O� $�@� Aؑ!p�PO��Z�xq0w�^�_MRAȑ_� d  T��-�ERR��ÏT)Yz�B�I�V3@�cNΑTOQ�d:`L� ��d2�p ��˰[! /� p�`T}0i��_V1�r�a'�
4�2-�2<����@Pq�����F�$W���g��V_!�l�$��P����c��q"�	�V FZN_CFG_!� 4��?º�|��ų����@�ȲW ��'��\$� � n���Ѵ��9c�Q��(��FA�He�,�XE�DM�(�����!s��Q�g�P{RV HEL}Lĥ� 56��B_BAS!�RSQR��ԣo �#S��T[��1r�%��2ݺU3ݺ4ݺ5ݺ6ݺ�7ݺ8ݷ��ROO0I䰝0�0NLK!�C�AB� ��ACK��IN��T:�1�@p�@ z�m�_PU!�CO� ��OU��P�� Ҧ) ��޶��T�PFWD_KAR�ӑ��RE~��P8��(��QUE������P
��CSTOPI_AL�����0&p���㰑�0SEMl�db�|�M��d�TY|�3SOK�}�DI����p�(���_TM\�MANRQ�ֿ0E�+�|�$KEYSWITCH&	����HE
�BEAT4����E� LEҒ��
�U��FO�����_O_HOM�O�7REF�PPRz�(�!&0��C+�OA��ECO��B�rI�OCM�D8׵�p]���8�` � D�1$����U��&�MH��<�P�CFORC���� ��OM�  �� @V��|�U�,3P� 1-�`� 3�-�4��NPX_�ASǢ� 0ȰA�DD����$SI}Z��$VARݷ. TIP]�\�2�A򻡐���]�_�$ �"S꣩!Cΐ��OFRIF⢞�S�"�c���NF��V ��n` � x�`SI��TES�R6SSGL(T�2P&��AU�<� ) STMTQZ�Pm 6BW�P*S�HOWb��SV|�\$�� ���A00P�a�6�@@�J�T�5�	U6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	f0 u�	�0u�	�@u�[Pu%121?1�L1Y1f1s2��	2�	2�	2�	2��	2�	2�	22�2%222?2�L2Y2f2s3�P)3�	3�	3�	3��	3�	3�	33�3%323?3�L3Y3f3s4�P)4�	4�	4�	4��	4�	4�	44�4%424?4�L4Y4f4s5�P)5�	5�	5�	5��	5�	5�	55�5%525?5�L5Y5f5s6�P)6�	6�	6�	6��	6�	6�	66�6%626?6�L6Y6f6s7�P)7�	7�	7�	7��	7�	7�	77�7%727?7�,i7Y7Fi7s�v�VP�UPD��  ��|�԰މ�YSLOǢ� � z��и���o��E��`>�^t��АAL1Uץ����CU���w=FOqID_L�ӿu�HI�zI�$FI�LE_���t��$�`�JvSA��� h����E_BLCK��#�C,�D_CPU<�{�<�o����txJr��R ��g
PW O� ��LA��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ� ��TBCu�C� ��X -$�LE�Ni��v������I���G�LOW_AXMI�F1��t2X�AM����D�
 ��I��s ��}�TOR�D���Dh��� L=���⇒�s���#�_M�A`�ޕ��ޑTCV����T���&���ݡ����J�����J$����Mo���J�Ǜ R�������2��`� v�����F�JK��CVKi�Ρv�Ρ3���J0�ңJJڣJJ�AALң�ڣ���4�5z�&�NA1-�9���␅�L~��_Vj�������� ` �GROU�pD��B�NFL�IC��REQUwIREa�EBUA�0�p����2¯����c�� \^��APPR��C����
�EN�CL9Oe��S_M v��,ɣ�
���� ���MC�&���g�'_MG�q�C� �p{�9���|�BRKz�GNOL��|ĉ R�Ї_LI|��Ǫ�k�J����P
���ڣ��� ��&���/���6��6���8������G� ��8�%�W�<2�e�PATHa�z�@p�z�=�vӥ�ϰ�x�CN=�CA�����6p�IN�UC��bqZ��CO�UM��YZ������qE%���2�������PAYLOA��J2L3pR_A	N��<�L��F�B�6��R�{�R_F2LS3HR��|�LOG�������ӎ���ACRL�_u�������.���H��p�$H{���FWLEX
��J�� :�/��� �6�2�����;�M�_�F16����n���������ȟ��Eҟ��� ��,�>�P�b��� d�{������������$5�T��X��v� ��EťmFѯ� ������&�/�A��S�e�D�Jx�� �� ������j�4pA�T����n�EL  ��%øJ���ʰJ�E��CTR�Ѭ�T�N��F&��HAN/D_VB[
�pnK�� $F2{�6� �rSW$#�U��� $$Mt�h�R��08��@<b 35��^6A�p3�k��q{9�t�A�̈p��A��A��ˆ0��U���D��Dʴ�P��G��ISTЙ�$A��$AN��DY ˀ�{�g4�5D���v� 6�v��5缧�^�@��P�����#�,�p5�>�(#�� &0��_�ER!V9�SQAS�YM��] �����px��ݑ���_SHl� ������sT�(����(�:�JA���S�ci\r��_VI�#Oh|9�``V_UNI��td�~�J���b�E�b ��d��d�f��n��� ������uN����D��H�������"CqEN� a�DI���>�Obt�'��Cqx�� ��2IxQA����q��-��s� �� ����� �^�OMME�h�rr�QTVpPT�P  ���qe�i����P��x ��yT�Pj� �$DUMMY9��$PS_��R�Fq�0$:� ����!~q� XX����K�STs�ʰ�SBR��M21_�Vt�8$SV_E�Rt�O��z���CLRx�A  O�r?p? �Oր � D ?$GLOB���#LO��Յ$�o���P�!SYSADqR�!?p�pTCHM0 � ,����oW_NA��/��e�����TSR~��l (: ]8:m�K6�^2m�i7 m�w9m��9���ǳ��� ����ŕߝ�9ŕ�� �i�L���m��_�_��_�TD�XSCRE��ƀ�� ��ST�F���}�pТ6��C�] _v AŁ� 9T����TYP�r�@K��u�!u���-O�@IS�!��tvC�UE{t� �����H�S���!RSM�_�XuUNEXCcEPWv��CpS_�� {ᦵ�ӕ���÷����COU ��� [1�O�UET�փr|���PROGM� {FLn!$CU��cPO*q��c�I_�p}H;� � 8��.N�_HE
p��Q�~�pRY ?����,�J�*��;�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�# m+�q��TR�IP)�m�UNjp{t� QP��XuoWARNWu�R�WTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� D�C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!& �VS�HIF��|s�P �p�6�s���R���OSURW�pRGADIz��2�_�q��h�g! �q)�L�Uza$OUTP�UT_BM��I�ML�oR6(`)�@T;IL<SCO�@Ce�;��9��F�� T��a��o�>�3�P����w�2u��tp�V�zu��%�DJ�U��|#�WAIET������%O{NE��YBOư� �� $�@p%�C�SBn)TPE��NEC��x"�$�t$���*B_T��R���%�qR� ���sB�%�tM�+��t�.耰F�R!݀��OPm�M�AS�_DOG�
OaT	�D����C3S�|	�O2DELAY���e2JO��n8E��S s4'#J�aP6%�����Y_��O2� �2�x��5��`? ���ZABCS�� � $�2��J�
0�  �$$CLA}S�����A�B���'@@VIRT8��O.@ABS�$��1 <E�� <  *AtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@��R�d�v�����M@[�A�XLր�&A�dC  ���IN��ā��GPRE������LARMRECOV <I䂥��NG�� \K	 =#�
J�\�M@�PPLIC�?�<E�E�H�andlingT�ool �� 
�V7.50P/2{8 *A�Hy���
�_SW�� �UP*A� ��F�0ڑ����A����� 20��*A��:�����FB 7DA�5�� '@�Iy@��No�ne������ ���T��*A4�9xx��P_���V����g�U[TOB ����~��HGAPON8@蕮LA��U��D 1-<EfA����������� Q 1EשI Ԁ�� Ԑ�:�i�n����#B�)B ����\�HE�Z�r�?HTTHKY��$B I�[�m�����	�c� -�?�Q�o�uχϙϫ� ���������_�)�;� M�k�q߃ߕߧ߹��� �����[�%�7�I�g� m����������� ��W�!�3�E�c�i�{� ��������������S /A_ew�� �����O+ =[as���� ���K//'/9/W/ ]/o/�/�/�/�/�/�/ �/G??#?5?S?Y?k? }?�?�?�?�?�?�?CO OO1OOOUOgOyO�O �O�O�O�O�O?_	__`-_K_Q_��(�TO4��s���DO_CLE�AN��e��SNM ; 9� �9o�Ko]ooo�o�DSP�DRYR�_%�HI��m@&o�o�o# 5GYk}���`�"���p�Ն �ǣ�qXՄ��ߢ��g�PLUGGҠ�Wߣ���PRC�`B`"9��o�=�OB��o^e�SEGF��K�� ����o%o����#�85�m���LAP�oݎ ����������џ������+�=�O�a���T�OTAL�.���U�SENUʀ׫ �X���R(�RG_S�TRING 1~��
�M���Sc�
��_ITwEM1 �  nc� �.�@�R�d�v����� ����п�����*��<�N�`�r�I/�O SIGNAL���Tryou�t Mode��Inp��Simu�lated�O�ut��OVE�RR�` = 10�0�In cy�cl���Pro?g Abor������Status��	Heartb�eat��MH �FaulB�K�AlerUم�s߅ߗߩ������������ �S���Q��f�x� ������������� �,�>�P�b�t�������,�WOR������ V��
.@Rd v��������*<N`PO��6ц��o�� ���//'/9/K/ ]/o/�/�/�/�/�/�/8�/�/�DEV�*0 �?Q?c?u?�?�?�? �?�?�?�?OO)O;O�MO_OqO�O�O�OPALTB��A���O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo8(o:o�OGRI�p�� ra�OLo�o�o�o�o�o �o*<N`r ������`o��RB���o�>�P�b� t���������Ώ��� ��(�:�L�^�p����PREG�N��.� �������*�<�N� `�r���������̯ޯ����&����$A�RG_��D ?	����i���  	]$��	[}�]}����Ǟ�\�SBN_�CONFIG �i�������C�II_SAVE � ��۱Ҳ\�T�CELLSETU�P i�%H?OME_IO�͈�?%MOV_�2ώ8�REP���V�U�TOBACK
��ƽFRA;:\�� �Ϩ���'` ��������� ����$��6�c�Z�lߙ��Ĉ�������������!� ����M�_�q���� 2���������%�7� ��[�m��������@� ������!3E$���Jo����\���INI�@���ε��MESS�AG����q��ODE_D$����O,0.��PAUS��!�i� ((Ol������ �� /�//$/Z/�H/~/l/�/�'akTSK  q������UPDT%�d�0;WSM_C5F°i�еU�>'1GRP 2h�93+ |�B��A�/S��XSCRD+11
N1; ����/ �?�?�? OO$O��� �?lO~O�O�O�O�O1O �OUO_ _2_D_V_h_��O	_X���GROU�N0O�SUP_N5AL�h�	�ĠV�_ED� 11;
� �%-BCKEDT-�_`�!oEo$���a��o��e���ߨ���eA2no_˔o�o�b����ee�o"�o�oED3 �o�o ~[�5GED4�n#��� ~�j���ED5 Z��Ǐ6� ~���}���ED6����k�ڏ� ~G���!�3�ED7 ��Z��~� ~�V�şןED8F�&o��Ů�}����i�{�ECD9ꯢ�W�Ư
}03�����CRo�� ���3�տ@ϯ����P~�PNO_DEL�_��RGE_UNUS�E�_�TLAL_OUT q�c�QWD_ABOR� ��΢Q��ITR_R�TN����NON�Se���CA�M_PARAM �1�U3
 8�
SONY XC�-56 2345�67890�H �� @���?}���( АVڪ|[r؀~�X�H�R5k�|U�Q�߿�R�57����Aff���KOWA S_C310M|[r�}̀�d @6� |V��_�Xϸ���V� �� ���$�6��Z�l���CE_RIA_UI857�F�1���R|]��_�LIO4W=� ��P<~�F<�GP ]1�,���_�GYk*C*  ���C1� 9� @Ң G� �CLC]�� d� l� s�R�� ��[�m� v� � �� �� +C�� �"�|W���7�HEӰONFI�� ��<G_PRI 1�+P�m®/ ��������'CHKPAUS� w 1E� ,� >/P/:/t/^/�/�/�/ �/�/�/�/?(??L?�6?\?�?"O��x���H�1_MOR��� ��PBZ�?����5 	  �9 O�?$OOHOZK�2D	���=9"�Q?5�5��C�PK�D3P������a�A-4�O__|Z
�O G_�7�PO�� ��6_��Y,xV�ADB���=�'�)
mc:cpmidbg�_`��S?:�  7;�P��Ŀ��Up�_)o�S g �C@��	f��P�_mo8j�  ׏`�Oko�oV9i�(�I(�JOk�g�o�o�li�j�Okf�oGq:I�ZD�EF f8��)��R6pbuf.t�xtm�]n�@�����# 	`(Ж�A=�L���zMC�21��=��9���4��=�n׾�Cz  �BHBCCPUeB���CF�;�.<C���C�5rSZE@D�n�yDQ��D���>��D��;D����F���>F�$G�}RB�GMzր��SY��!�vJqG���Em�(�U.��(�(��<�Lq�G�x2��Ң ��� a�D�j���E�S\E@EX�E�Q�EJP F��E�F� G��ǎ^F E��� FB� H�,- Ge��H�3Y���  >�33 ���NxV  n2xQ@��#5Y��8B� A�ASTo<#�
� �_�'�%��wRSMOF�S���~2�yT1>�0DE �O@b� 
�(�;�"� � <�6�z�R��X�?�j�C4��SZ�m� W��{�m�CR��B-G�Cu�@$��q��T{�FPROG %i�����c�I��� �Ɯ�f�K�EY_TBL  �vM�u� �	
��� !"#�$%&'()*+�,-./01c�:�;<=>?@AB�C�pGHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������p����͓���������������������������������耇��������������������!j�LCK��.�j����STAT���_A�UTO_DO����W/�INDT_ENB߿2R��9�+��T2w�XSTOP�\߿2TRLl�LE�TE����_SCREEN i�kcsc��U���MMENU 1� i  < g\��L�SU+�U��p3 g������������ 2�	��A�z�Q�c��� ������������. d;M�q�� ����N% 7]�m��� /��/J/!/3/�/ W/i/�/�/�/�/�/�/ �/4???j?A?S?y? �?�?�?�?�?�?O�? O-OfO=OOO�OsO�O �O�O�O�O_�O_P_�Sy�_MANUAyL��n�DBCOU��RIG���DBN�UM�p��<���
��QPXWORK 1!R�ү�_oO�.o@oRk�Q_AWA�Y�S��GCP r��=��df_AL�P�db�RY�������X�_�p 1"�� , 
�^���o �xvf`MT�I^�rl@|�:sONTIM�כ����Zv�i
�õ�cMOTNEN�D���dRECOR/D 1(R�a��ua�O��q��sb �.�@�R��xZ���� ���ɏۏ폄���#� ��G���k�}�����<� ş4��X���1�C� ��g�֟��������ӯ �T�	�x�-���Q�c� u����������>�� ��)Ϙ�Mϼ�F�� �ϧϹ���:������� %�s`Pn&�]�o��ϓ� ~ߌ���8�J����� 5� ��k����ߡ�� J�����X��|��C� U����������0������	��dbTOL�ERENCqdB�ܺb`L�͐PCS_CFG )�k�)wdMC:\�O L%04d.C�SV
�Pc�)sA� �CH� z�P�)~���hMRC_OUT *�[��`+P SGN �+�e�r��#��10-MAY-20 08:57*V�27-JANj2�1:48�k P;���)~��`pa�m���PJPѬV�ERSION �SV2.0�.�6tEFLOG�IC 1,�[ 	DX�P7)�PF.�"PROG_ENqB�o�rj ULSew� �T�"_WRS�TJNEp�V�r`dE�MO_OPT_S�L ?	�es
 	R575)s 7)�/??*?<?'�$TO  �-��?�&V_@pEX�Wd��u�3PATH ;ASA\�?�?\O/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C���SqqF�PMAqU� t/XrMSWR�.�i6.|S/�Z!D_N�O0__T_�C_x_g_�_�tSBL__FAUL"0�[^3wTDIAU 16M�6p�A1�234567890gFP?BoTo foxo�o�o�o�o�o�o �o,>Pb�SZ�pP�_ ���_ s�� 0`���� �)�;�M�_�q����������ˏݏ��|)U3MP�!� �^��TR�B�#+�=�PM�EfEI�Y_TEM=P9 È�3@�3�A v�UNI�.(Y�N_BRK 2�Y)EMGDI_�STA�%WЕNC�2_SCR 3��1o"�4�F�X�fv ���������#��ޑ14����)�;������ݤ5��� ��x�f	u�ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/߭P�b�t�� �� xߞ߰���������
� �.�@�R�d�v��� �����������*� <�N���r��������� ������&8J \n������ ��"`�FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/4? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O ?�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�O�O�o�o�o
 .@Rdv�� �������*� <�N�`�r����o���� ̏ޏ����&�8�J� \�n���������ȟڟ�����H�ETMO�DE 16���� ��ƨ
�R�d�v�נRROR�_PROG %fA�%�:߽�  ���TABLE  �A������#�L�R�RSEV_NUM�  ��Q���K�S���_AUT�O_ENB  ���I�Ϥ_NOh� �7A�{�R� W *���������	���^�+��Ŀֿ���HISO�͡I�}�_ALM 18A�� �;�����+�e�wωϛϭϿ�r�_H���  A����|��4�TCP_VER !A��!����$EXTL�OG_REQ�9�{�V�SIZ_�QԿTOL  ͡D}z��=#׍�?XT_BWD���иr���n�_DI�� 9��}�z�͡<m���STEP����|4��OP_DO����ѠFACTO�RY_TUN�d�G�EATURE �:����l��Handlin�gTool �� � - CEn�glish Di�ctionary���ORDEA�A Vis�� M�aster���9�6 H��nalo�g I/O���H�551��uto �Software� Update � ��J��mati�c Backup~��Part&��ground E�dit��  8\�apCame�ra��F��t\j�6R�ell���LwOADR�omm���shq��TI" ��co��
! yo���pane��� 
!��ty�le selec]t��H59��nD�~��onitor��48����tr��R�eliab���a�dinDiagnos"����2��2 ual Che�ck Safet�y UIF lg�\a��hance�d Rob Se�rv q ct\���lUser F�rU��DIF��E�xt. DIO 6��fiA d��wendr Err YL@��IF�r�ನ  �П�90��F�CTN Menu�Z v'��74� T�P In��fac�  SU (�G=�p��k E�xcn g�3��High-Sper wSki+�  sO��H9 � mmuni]c!�onsg�te�ur� ����V��y��conn���2��EN��Inc=rstru����5.fdKA�REL Cmd.� L?uaA� O~�Run-Ti� 'Env����K� ��u+%�s#�S/W���74��Licen�seT�  (A�u* ogBook�(Sy��m)��"�
MACR�Os,V/Off�se��ap��MH�� ����pfa5�M�echStop �Prot��� d��b i�Shif����j545�!x�r ��#��,K��b ode Swiwtch��m\e�!�o4.�& pr�o�4��g��M?ulti-T7G����net.P{os Regi���z�P��t Fu9n���3 Rz1���Numx �����9�m�1�  Adju<j��1 J7�7�*� ����6tatu�q1EIKRD�Mtot��scove�� ��@By<- }uest1�$G�o� � U5\SNPX b"���<YA�"Libr��㈶�#�� �$~@h�p�d]0�Jts i?n VCCM����ĕ0�  �u!��2 �R�0�/I�08~��TMILIB�M� J92�@P�A�cc>�F�97�TgPTX�+�BRSQselZ0�M8 Rm��q%��692��Unexceptr �motnT  CcVV�P���KC�����+-��~K  I�I)�VSP CSXC�&.c�� e�"��� t�@We�w�AD Q�8bv9r nmen�@�KiP� a0y�0��pfGridAplay !� nh�@*��3R�1M-10iA�(B201 �`2�V"  F���sci�i�load��8�3 M��l����G�uar�d J85��0�mP'�L`���s�tuaPat�&]$C�yc���|0ori�_ x%Data'Pqu���ch�1���g`� j� RLJa�m�5���IMI �De-B(\A�cP"� #^0C  e�tkc^0assw�o%q�)650�Ap�U�Xnt��PvKen�CTqH�5�0�YELLOW� BO?Y��� Arc�0vis��C�h�WeldQci�al4Izt�Op�� ��gs�` 2@�a6��poG yRjcT1 NE�#HTf� xyWb��! �p��`gd`���p\� �=P��JPN ARCP*PR�A�� �OL�pSup̂fil�p��J�� n��cro�670�1�C~E�d��SS�pe.�tex�$ �P� �So7 t� ssa%gN5 <Q�BP:� 2�9 "0�QrtQCr��P�l0dpn������rpf�q�e�ppm�ascbin�4psyn�' pstx]08�HEL�NCL VIS �PKGS �Z@M�B &��B J8�@IPE GET_VAR FI?S_ (Uni� LU��OOL: ADD��@29.FD�TC4m���E�@DVp����`A�ТNO WT?WTEST �� �V�!��c�FOR ^��ECT �a!� �ALSE ALA�`�CPMO-13�0��� b D: H�ANG FROM�g��2��R709� DRAM AV�AILCHECK�S 549��m�V�PCS SU֐L_IMCHK��P�0~x�FF POS� �F�� q8-12 CHARS��ER6�OGRA ���Z@AVEH�AME��.SV��Вאqn$��9�m "y��TRCv� SHA�DP�UPDAT �k�0��STATI���� MUCH ����TIMQ MOTN-003���@OBOGUI�DE DAUGH໱�b��@$tou�� �@C� �0��PA�TH�_�MOVE�T�� R64��V�MXPACK M�AY ASSERyTjS��CYCL`��TA��BE CO�R 71�1-�AN���RC OPTI�ONS  �`��A�PSH-1�`fi	x��2�SO��B��XO򝡞�_T��	�i�j�0j��du�byz �p wa��y�٠H�I������U�pb X?SPD TB/�F�_ \hchΤB0����END�CE�06�\Q�p{ sma'y n@�pk��L} ��traff#��	� ��~1fro�m sysvar/ scr�0R� ��Nd�DJU���H��!A��/��SET GERR�D�P7�����NDANT S�CREEN UNREA VM �P�D�D��PA���R~�IO JNN�0��FI��B��GRwOUNנD Y��Т٠�h�SVIP� 53 QS��DI�GIT VERS���ká�NEW�� �P06�@C�1IMCAG�ͱ���8� �DI`���pSSU�E�5��EPLAN� JON� DELL���157QאD��CALLI���Q��m���IPND}�IMG N9 PZ�{19��MNT/���ES ���`LocR Hol߀=��2�P�n� PG:��=�M��can����С�: 3D mE2view d X���ea1 �0b�po;f Ǡ"HCɰ��ANNOT AC�CESS M c�pie$Et.Qs �a� loMdFle�x)a:��w$qmo+ G�sA9�-'p~0̿�h0pa��eJ AUTO-�0��!�ipu@Т<ᡠIA�BLE+� 7�a F�PLN: L�p�l m� MD<�V�I�и�WIT H�OC�Jo~1Qu�i��"��N��US�B�@�Pt & r�emov���D�vAxis FT_7�PGɰCP:�O�S-144 � h� s 268QՐO�ST�p  CRA�SH DU��$P~��WORD.$��LOGIN�P��P�:	�0�046 i�ssueE�H�:� Slow st�c�`6�����z��IF�IMPR��SPOT:Wh4����N1STY��0V�MGR�b�N�CA�T��4oRRE�� �� 58�1��:N%�RTU!Pe -M .a�SE:�@pp���$AGpL��m@�all��*0a�OC�B WA���"3 �CNT0 T9DW�roO0alarm8�ˀm0d t�M��"0�2|� o�Z@O�ME<�� ��E%  ;#1-�SRE��M��st}0g   �  5KANJI~5no MNS@��INISITA7LIZ'� E�f�cwe��6@� dr�@� fp "��SC�II L�afai�ls w��SY�STE[�i�� � � Mq�1QGro8�m n�@vA�����&��n�0q��R�WRI OF L|k��� \ref"��
�up� de-r�ela�Qd 03�.�0SSchőb�etwe4�INDo ex ɰTPa�#DO� l� �ɰ�GigE�sope�rabil`p l�,��HcB��@]�lye�Q0cflxz�8Ð���OS {�����v4pfigi GL�A�$�c2�7H� wlap�0ASB� �If��g�2 l\�c�0�/�E�� �EXCE 㰁�P����i�� o0��G�d`]Ц�fq�l lsxt��EFal����#0�i�O�Y�n�CL�OS��SRNq1NT^�F�U��FqKP~�ANIO V7/�¥�1�{����DBa �0��ᴥ�ED��DET|�'� �b�F�NLINEb�B�UG�T���C"RL�IB��A��ABC? JARKY@���� rkey�`IL����PR��N��ITG+AR� D$�R �Er *�T��a�U�0��h�[�ZE V�� TASK p7.vr�P2" .�XfJ�srn�S谥d�IBP	c���B/��BUS��UNN�� j0-�{��cR�'���LOE�DIVS�CULs$cb����BW!��R~�W`�P�����IT(঱t�ʠ�OF��UNE�Xڠ+���p�FtE���SVEMG3`N�ML 505� D�*�CC_SAFE��P*� �ꐺ� PE�T��'P�`�F  �!���IR����c Ri S>� K��K��H GUNCHGz��S�MECH��IM��T*�%p6u���tPORY LE�AK�J���SP�EgD��2V 74\GRI��Q�g��oCTLN��TRe `@�_�p ���EN'�IN������$���r��T3)�i�STO��A�s�L��͐X	���q��Y� ��CTO2�J m��0F<�K����DU�S��O���3 9�J F��&���SSVGN�-1#I���RSRwQDAU�Cޱ� �T6��g��� 3�]���BR�KCTR/"� �q\�j5��_�Q�S�qI{NVJ0D ZO�P ݲ���s��г�Ui ɰx̒�a�DUAL�� J50e�x�RV�O117 AW�T�H!Hr%�N�247�%�52��|�&aol� ���R���at�Sd��cU���P,�LER��iԗQ0�ؖ  S!T���Md�Rǰt�_ \fosB�A�0@Np�c����{�U���ROP 2�b�pB>��ITP4M��b !AUt c0< � �plete�N@�� z1^qR635� (AccuCa�l2kA���I) �"�ǰ�1a\�Ps ��ǐ� bЧ0P������ig\cba?cul "A3p_ �1��ն���eta�ca��AT���PC��`�����_p�.�pc!Ɗ��:�cicrcB���5�tl��Bɵ�:�fm+�Ί��V�b�ɦ�r�upf�rm.����ⴊ�x�ed��Ί�~�ped�A�D �}b�ptl�ibB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆Ϙ���c�Ӳ�5�1j>�����tcȐ�Ϣ	�r����mm 1���T�sl^0��T�m�ѡ�#�rm3��u8b Y�q�std}��3pl;�&�ckv�=߆r�vf�䊰��9�v1i����ul�`�04fp�q �.f���� daq; i Da�ta Acqui+si��n�
��4T`��1�89���22 DMCM oRRS2Z�75���9 3 R710,�o59p5\?T "��1 (D�T� nk@���� ����E Ƒȵ��Ӹ��etdmm ��ER�����gE��1�q\mo?۳�=( G���[(

�2�` �! �@JMAC�RO��Skip/Offse:�a���V�4o9� &qR6C62���s�H��
 6Bq8����9~Z�43 J77� =6�J783�o `��n�"v�R5�IKCBq2 PT�LC�Zg R�3; (�s, �������03�	зJ���\sfmnmc? "MNMC�����ҹ�%mnf�FM�C"Ѻ0ª etm�cr� �8����� ,K�D�V�   874\prdq>�,jF0���axi�sHProcess Axes e�wrol^PRA
��Dp� 56 J81�j�59� 56o6�� ���0w�690 998� [!IDV�1��2(x2��2ont �0�
����m2����?C��etis "ISD��9�� F/praxRAM�P�8 D��defB�,��G�isbasicHB�@޲{6�� W708�6��(�Acw:������D
�/,��AMOX�� ��DvE ��?;T��>Pi� RACFM';�]�!PAM�V �W�Ee�U�Q'
bU�75�.�ceN�e� nterfa�ce^�1' 5&!5�4�K��b(Dev am±�/�#���/<�Tazne`"DNEWE����btpdnui� �AI�_s2�d_rsono���bAs�fjN��bdv_arFvf�xhpz�}w��shkH9xstc��gAponlGzv{�ff��r���z��3{q'Td>pcOhampr;e�p� ^5977��	܀�4}0��mɁ�/�����l�f�!�pcchmp�]aMP&B�� �m�pev�����p�cs��YeS�� M/acro�OD��16Q!)*�:$�2U"_,x��Y�(PC ���$_;������o��J�g�egemQ@GEM�SW�~ZG�gesn�dy��OD�ndda��S��syT�Kɓ�Csu^Ҋ���n�m��<�L��  ���9:�p'ѳ޲��spotplusp���`P-�W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\f�eatu 0FEA�WD�oolo�s�rn'!2 p���a؝As3��tT.� (?N. A.)��!�e!�J# (j�,`��oBIB�oD -��.�n��k9�"K���u[-�_���p� "PSEqW����?wop "sEЅ� &�:�J������y�|� �O8��5��Rɺ��� ɰ[��X������ـ%�(
ҭ�q HL �0k�
�z�a!�B�Q�"(g�Q����� ]�'�.�����&���<�0!ҝ_�#��tpJ�H� ~Z��j�����y���� ��2��e������Z�� ��V��!%���=�]�p͂��^2�@iRV� Kon�QYq͋JF0B� 8ހ�`�	(^>�dQueue���X�\1�ʖ`�+F1tpv�tsn��N&��ftupJ0v �RDV�	�f��J1 Q���v��en��kvst�k��mp��btk�clrq���get����r��`kack�XZ��strŬ�%�st0l��~Z�np:!�`����q/�ڡ6!l��/Yr�mc�N+v�3�_� ����.�v�/\jF���� �`Q�΋ܒ�N50 (FRA��+�����fraparm���Ҁ�} 6�J6�43p:V�ELSE�
#�VAR $�SGSYSCFG�.$�`_UNITS 2�DG~°@�4�Jgfr��4A�@FRL-��0ͅ�3ې���L �0NE�:�=�?@�8 �v�9~Qx304��;�BPRSM~QA��5TX.$VNUM_OL��5��DJ�507��l� Functʂ"qwAP��琉�3 H�ƞ�kP	9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TP�PR���QA�prnaSV�ZS��AS8D�j510U�-�`cAr�`8 ��ʇ�DJR`�jYȑH  ��Q �PJ6�a2�1��48AA�VM 5�Q�b0 �lB�`TUP xb?J545 `b�`�616���0V�CAM 9�CwLIO b1�s5 ���`MSC8��
rP R`\s�STYL MNI�N�`J628Q  �`NREd�;@�`�SCH ��9pDCSU Mete�`�ORSR Ԃ�a0�4 kREIO�C �a5�`542�b9vpP<�nP�a�`�R�`7�`�M?ASK Ho�.r�7 �2�`OCO :��r3��p�b�p���r0X��a�`13\�mn�a39 HR�M"�q�q��L�CHK�uOPLG� B��a03 �q.��pHCR Ob�pC�pPosi�`fP6� is[rJ554��òpDSW�bM�D8�pqR�a37 }Rjr30 �1�s4 �R6�m7��52�r5 �2.�r7 1� P6����Regi�@T^�uFRDM�uSaq�%�4�`930�uS�NBA�uSHLB�̀\sf"pM�N{PI�SPVC�oJ520��TC�`�"MNрTMIL��IFV�PAC �W�pTPTXp6�.%�TELN N� Me�09m3�UECK�b�`U�FR�`��VCOR^��VIPLpq89q�SXC�S�`VVF��J�TP �q��Rw626l�u S�`�Gސ�2IGU�I�C��PGSt�\ŀH863�S�q������q34sŁ6�84���a�@b>�3� :B��1 T��9�6 .�+E�51 �y�q53�3�b1 ̛��b1 n�jr9 <���`VAT ߲�q�75 s�F��`�sA�WSM��`TOP u�ŀR52p���a�80 
�ށXY �q���0 ,b�`8855�QXрOLp}��"pE࠱tp�`LCyMD��ETSS�挀6 �V�CPEs oZ1�VRCd3�
�NLH�h��0011m2Ep��3 f��p���4 /165CR��6l���7PR���008 tB��9 o-200�`U0�p�F�1޲1 ��޲2 L"���p��޲4���5 \hmp޲6 RBCF�`ళ�fs�8 �Ҋ��~�J�?7 rbcfA�L��8\PC����"�32�m0u�n�K�Rٰn�5� 5EW
n�99 z��40 kB���3 ��6ݲ�`00�iB/��6�u��7�u��8 µ������s�U0�`�t �1 0�5\rb��2 E@���K���j���5˰��60��a�HУ`:Ł63�jAF�_���F�7 ڱ݀H�8�eHЋ�&�cU0��7�p���1u��8u��9 c73������D7� r��5t�97 ��E8U�1��2��1�)1:���h��1np�"���8(�U1��\pyl��,࿱v ��B�854��1V���D�-4��im��1�<����>br�3pr�48@pGPr�6 B����$�p��1����1�`͵�155ض157 �2��62�S����B��1b��2����1Π2"�2���B6`�1<c�4 7B�5i DR��8_�B/���187 uJ�8 ;06�90 rBn��1 (��202 /0EW,ѱ2^��2��90�U2�p�2��S2 b��4��2�a�"RB����9\�U�2�`w�l���4 6	0Mp��7������b�,s
5 ��3����<pB"9 3 ����l�`ڰR,:7 �2��V�2��5���2^H��a^9���qr�����n�5����5᥁""�8a�Ɂ}�5B���5����`UA���� ���86 �6 S�0�5�p�2�#�52�9 �2^�b1
P�5~�2`���&P*5��8��5��u�r!�5��ٵ544��%5��R�ąP nB^,z�c (�4���L���U5J�V�5��1�1^��%�����5 b21��gA���58W82� r�b��5N�E�589�0r� 1�95  �"������c8"a��|�L ���!J"5|6���^!�6��B�"8P�`#��+�8%�6B��AME�"1 iCN��622�Bu�6V���d� 4��84�`A�NRSP�e/S� C�5� �6� ��� \� �6� �V� 3�t��� T20CA�R��8� Hf� 1D�H�� AOE� ��� ,K|�� a�0\�� �!64K���ԓrA� �1 (M{-7�!/50T� [PM��P�Th:1�C��#Pe� �3�0� 5>`M75T"� �D�8p� �0Gc� u�4|��i1-710i�1B� Skd�7j�?6�:-HS,� �RN�@��UB�f�X�=m7C5sA*A6an���!X/CB�B2.6A �0 ;A�CIB�A�2�QF1�U�B2�21� /70�S� �4����Aj1��3p���r#0 B2\m*A@C��;bi"�i1K�u"A~AAU� imm7c7��ZA@HI�@�Df�A�D5*A��E� 0TkdR1�35�Q1�"*�@�Q�1�QC )P�1*A�5*A�EA�5XB�4>\77
B7=Q �D�2�Q$B�E7�C�D%/qAHEE�W7�_|` jz@� 2�0�Ejc�7�`�E"l7�@7@�A
1�E�V~`�W2%Qr�R9ї@0L_�#�����"A���b��H3s=rA/2�R5nR 4�74rNUQ1ZU�A�sw\m9
1M92L2��!F!^Y�ps� 2c1i��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHsXBSt62�q`s������ ��Pxq3530_*A3I)�2�db�u0�@� '4TX�m0�pa3i1A3s0Q25�c��st�r�VR1%e�q0
��j1 ��O2 �A�UEiy�@.�‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?P Q��qA!Pvs� 5	1 5aU���?PŅ���ဝQ9A6�zS*�7�qb5�1����Q��'00P(��V7]u�a itE1���ïp?7� �!?�z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ�޵y00\ry�"R�2BL�tN  ���� �1DVA��2�qeR�5���_b�3�X]1m1l�cqP1�a�E�Q� 5�F����!5���@M-16Q�� f���r���Q�e� ��� PN�L�T_�1��i1��945�3��@�e�|�b1l>F1u*AY2�
�R8�Q����RJ�J13�D}T� 85
Qg� /0��*A!P�*A�Ð�d����2ǿپ6t�6=Q���Pȓ��� AQ� g�*ASt]1 ^u�ajrI�B����~`�|I�b��yI�\m�Qb�I�uz�A�c3Apa\9q� B6S��S��m���}�85`N�N�  �(M�� �f1���6����161j��5�s`�SC���U��A����5\se�t06c����10��y�h8��a6��6x��9r�2HS �� �Er���W@}�a��IlB���Y�ٖ�m�u �C����5�B��B��h`�F���X0���A :���C�M��AZ��@��4�6i����� e�O�-	���f1��F  �ᱦ�1F�Y	���GT6HL3��U66~`Ȗ��U�dU�9D20Lf0��Qv� ��fjq ��N������0v
� ���i	�	��72l�qQ2������� \�chngmove�.V��d���@2l_arf	�f ~��6������9C��Z���~���kr41@ S���0��V��t�����U�p7nu�qQ%�A]��V�1\"�Qn�BJ�2W� EM!5���)�#:��64��F�e50S �\��0�=�PV�� �e������E������m7shqQSH"U��)��9�!A���(���� �,K��ॲTR11!��,�60e=��4F�����2��	 R-����������@�Ж��4���LS0R�)"�!lOA��Q�X) %!� 16�
U /��2�"2�E�9p���2>X� SA/i��'�
7F�H�@!B�0�� �D���5V��@2cV E��p��T��pt갖��1L~E�#�F�Q��9�E�#De/��RT��59���	�A�EiR���|����9\m20챃20��+�-u�19r4 �`�E1�=`O9`� �1"ae��O�2��_\$W}am41�4�3��/d1c_std ��1)�!�`_T��r~�_ 4\jdg�a �q�PJ%!~`-�r�+�bgB��#c300D�Y�5j�QpQb1�`bq��vB��v25�Up�����qm43�  �Q<W�"PsA��e ����t�i�P�W .��c�FX.�e4�kE14�44�~o6\j4�443sxj��r�j4up�� �\E19�h�PA�T�= :o�APf��coWol!\�2a��2A;_	2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a�:88J9X�l5�m�1a첚��*���(85�&�������P6���R,52&A����,fA9IfI50\u�z�OV
�v��}E�֖J���Y>� 16�r�C�Y��;��1��L ���Aq�&ŦP1��vB�)e�m�����1pĻ �1DV��27��F�KAREL �Use S��FC�TN��� J970�FA+�� (�Q޵0�p%�)?�Vj9F?(��j�Rtk208 C"Km�6Q�y�j��iæPr�9�s#��v��krcfp�RCF�t3���Q��kcctme�!ME�g����^6�main�dV�� ��ru��kDº��c���o����J�dt��F �»�.vrT�f�����E%�!��\5�FRj73B�K����UER�HJ�O  �J�� (ڳF���F �q�Y�&T��p�F�z��19�tkvBr���V�Bh�9p�E�y�<�k�������;�v���"CT��f����)�
І ��)�V	�6���!� �qFF��1q���=��� ��O�?�$"���$���je���TCP A�ut�r�<520 �H5�J53E19�3��9��96�!8���9��	 �B574V��52�Je�(�� Se%!Y�����u���ma�Pqtool��ԕ������co�nrel�Ftro�l Reliab�le�RmvCU!��H51����� a�551e"�CNRE¹I�c�&���it�l\sfut?st "UTա��"X�\u��g@�i�D6Q]V0�B,Eѝ6A� �Q�)C���X���Yf�I�1|6s@6i��T6IU��vR��d�
$e%1��2�C58�E6��8�Pv�iV�4OFH58SOeJ� mnvBM6E~O58�I �0�E�#+@�&�F�0 ���F�P6a���)/++��</N)0\tr1x�����P ,K�ɶ��rmaski�ms�k�aA���ky'd�h�	A	�P�sDisp_layIm�`v��~��J887 ("A��+Heůצprd�s��Iϩǅ�h�0p�l�2�R2��:�Gt�@��PRD�TɈ�r��C�@Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��Px^@�P�firmQ� ���Pp�2�=bk�6�r��3��6��tppl��PL���O�p<b�ac�q	��g1J�U�d0�J��gait_9e���Y�&��Q���	�S�hap��erat�ion�0��R6�7451j9(`sGen�ms�42-f�Ár�p�5����2�rsgl�E��p�G���qF�205p�5S���ՁN�retsap�BP�O��\s� "GC�R�ö? �qngda�G��V��st2axU��Aa]��b�ad�_�btpu�tl/�&�e���tp�libB_��=�2.p����5���cird��v�slp��x�hex��v�re?�Ɵx�gkey�v�pm���x�us$�6�gcr��F������[�q27�j92�v�ollismqSk�9O��>�� (pl.���t��p!o��29$Fo8���cg7no@�tptwcls` CLS�o�b�\�km�ai_
�!s>�v�o	�t�b��x�ӿ�E�H��6~�1enu501�[�m��utia|$c�almaUR��Ca�lMateT;R5	1%�i=1]@-��/V�� ��Z�� �fq1�9 "K9E�L����z2m�CLMTq��S#��et �LM�3!} �F�c�ns�pQ�c���c_mo4q��� ��c_e���F��su��ޏ �_ �x@�5�G�join�@i�j��oX���&cW0v	 ���N�ve��C�clm�&Ao# �|$�finde�0�STD ter� FiLANiG���R��
��8n3��z0Cen���r,������J��� �� ���K��Ú�=�К�_Ӛ��r� "FNDR�� 3��}f��tguid��`��N�."��J�tq��  �������������J����_������c���	m�Z��\fndr.��n#>
B2�p��Z�CP Ma�����38A��� c
��6� (���N�B ������� 2�$�	81��m_���"ex�z5�.Ӛ��c���bSа�ef�Q��	��RBT~;�OPTN � +#Q�*$�r*$��*$r *$%/s#C�d/.,P�/|0*ʲDPN���$���$*�Gr�$ko Exc�'IF�$�MASK�%93 {H5�%H558�$_548 H�$4-1��$��#1(�$�0 E�$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3��9j0"M�49�4 � ��4�4tp�sh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E�\���5�A�4��3a�dq\�5K979�":E�ajO l "�DQ^E^�3i�Dq� ��4ҲO ?R�? ��q�5��T��3rAq�O�Lst�5~��7�p�5��REJ#�2�@a�v^Eͱ�F���4��.��5y N� �2il�(in�4��31 aJH1�2Q4�251ݠ��4rmal� �3) �REo�Z_�æOx�����4��^F�?onor Tf��7_ja�UZҒ4l��5rmsAU�Kkg���4�$HCd\�fͲ�e�ڱ�4�REM���4y�ݱ"u@�RER593�2fO��47Z��5lity,�U��e"DGil\�5��o ��7987�?�25 �3hk910�3���FE�0=0P_�Hl\mhm�5��qe�=$��^�
E��u�IAymptm�U��BU��vste�y\�3��me� b�DvI�[�Qu�:F�U�b�*_�
E,�su$��_ Er��oxx���4huse�E-�?�sn�������FE��,�box�����c݌,"��������z��M��g��pdspw)�	��9��� b���(��1�� �c��Y�R�� �>�P� ��W��������'��0ɵ�[��͂����  � ,KN@� �A��bumpšf��B*�Box%��7Aǰ�60�BBw���MC� u(6�,f�t I�s� ST��*���}B�����w��"BBF
�>�`���)���\bbk968� "�4�ω�bb��9va69����etbŠ��X�����#ed	�F��u�f�& �sea"������'�\��,���b�ѽ"�o6�H�
�x�$�f���!y���Q[�!� tperr�f�d� TPl0o� R/ecov,��3D���R642 � 0���C@}s� N@��(NU�rro���yu2�r��  �
�  ����$$�CLe� �������������$~z�_DIGIT��.������ .�@�R�d�v������� ��������*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_��_ oo$j��+c:PRODUCTM��0\PGSTKD��V&ohozf99���D���$F�EAT_INDE�X��xd���  
�`IL�ECOMP ;����#��`�cS�ETUP2 <��e�b�  �N �a�c_AP2�BCK 1=�i  �)wh0?{%&c����Q� xe%�I�m�� �8��\�n����!� ��ȏW��{��"��� F�Տj���w���/�ğ S���������B�T� �x������=�үa� �����,���P�߯t� �����9�ο�o�� ��(�:�ɿ^���� �ϸ�G���k� �ߡ� 6���Z�l��ϐ�ߴ� ��U���y����D� ��h��ߌ��-���Q� ��������@�R��� v����)�����_��� ��*��N��r� �7��m�@&�3\�i
pP� 2#p*.V1Rc�*��`� /��PC/|1/FR6:/"].��/+T�`�/ �/F%�/�,�`r/?��*.F�8?	�H#&?e<�/�?;STM �2�?�.K �?��=iPen�dant Panel�?;H�?@O�7�.O�?y?�O:GIF �O�O�5�OoO�O_:JPG _J_�56_�O�_�_�	PANE�L1.DT�_@�0�_�_�?O�_2�_�So�WAo�_o�o�Z3 qo�o�W�o�o�o)�Z4�o[�WI���
TPEINSO.XML��0�\���qCust�om Toolb�ar	��PAS�SWORDy�FRS:\L�� �%Passwo�rd Config���֏e�Ϗ�B 0���T�f�������� ��O��s������>� ͟b��[���'���K� �򯁯���:�L�ۯ p�����#�5�ʿY�� }��$ϳ�H�׿l�~� Ϣ�1�����g��ϋ�  ߯���V���z�	�s� ��?���c���
��.� ��R�d��߈���;� M���q������<��� `������%���I��� �����8����n ���!��W�{ "�F�j| �/�Se��/ �/T/�x//�/�/ =/�/a/�/?�/,?�/ P?�/�/�??�?9?�? �?o?O�?(O:O�?^O �?�O�O#O�OGO�OkO }O_�O6_�O/_l_�O �__�_�_U_�_y_o  o�_Do�_ho�_	o�o -o�oQo�o�o�o�o @R�ov��; �_���*��N� �G������7�̏ޏ m����&�8�Ǐ\�� ���!���E�ڟi�ӟ ���4�ßX�j����� ���įS��w�������B�#��$FIL�E_DGBCK �1=��/���� ( ��)
SUMMA�RY.DGL����MD:������Diag Sum�mary��Ϊ
C?ONSLOG������D�ӱCon�sole log�E�ͫ��MEMCHECK:�!ϯ����X�Memory� Data��ѧ��{)��HAD�OW�ϣϵ�J����Shadow C?hangesM�'��-��)	FTAP7Ϥ�3ߨ���Z��mment TB�D��ѧ0=4)�ETHERNET��������T�ӱE�thernet �\�figurat�ionU�ؠ��DCSVRF�߽߫������%�� ve�rify all���'�1PY���DIFF�����[����%��diff]������1R�9�K���� ���X=��CHGD������c��r�����2ZAS� ��GD����k��z��FY�3bI[� �/"GD����s/����/*&UPDATES.� ��/��FRS:\��/�-ԱUpda�tes List��/��PSRBWLOD.CM(?���"�<?�/Y�PS_ROBOWEL��̯�? �?��?&�O-O�?QO �?uOOnO�O:O�O^O �O_�O)_�OM___�O �__�_�_H_�_l_o �_�_7o�_[o�_lo�o  o�oDo�o�ozo�o 3E�oi�o�� �R�v���A� �e�w����*���я `���������O�ޏ s������8�͟\�� ���'���K�]�쟁� ���4���ۯj����� �5�įY��}���� ��B�׿�x�Ϝ�1� ��*�g�����Ϝ��� P���t�	�ߪ�?��� c�u�ߙ�(߽�L߶� �߂���(�M���q�  ���6���Z���� ��%���I���B������2�����h�����$FILE_� P�R� ��������M�DONLY 1=�.�� 
 � ��q��������� �~%�I�m �2��h� �!/�./W/�{/
/ �/�/@/�/d/�/?�/ /?�/S?e?�/�??�? <?�?�?r?O�?+O=O �?aO�?�O�O&O�OJO �O�O�O_�O9_�OF_�o_
VISBCK�L6[*.VD�v_�_.PFR:\��_�^.PVis�ion VD file�_�O4oFo\_ joT_�oo�o�oSo�o wo�oB�of�o �+����� ��+�P��t���� ��9�Ώ]�򏁏��(� ��L�^�������5� ��ܟk� ���$�6�ş�Z��~�����
M�R_GRP 1>�.L��C4 w B���	 W������*u����RHB ���2 ��� ��� ���B� ����Z�l���C���D�ি����Ŀ��J�8�L���J�a�F�5U��R�e����ֿ �Gn�E��.�E88�-���?:u�{@ �����@A�A��a�f�?h!A����r��E�� F�@ ������ھ���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6�\b��B�Y<%���AD��=�@�0eߋ�NҞ�A��߲� v���r������
�C� .�@�y�d������ ��������?�Z�l�v��BH�� ��R�?�VE��������
0�PJ��P��H��ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�OPгߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������/[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U��0
//./A�#��� �~/����/�/�/ �/� ?2?D?V?h?�/ ?�?�?�?�?�?�?� ��@O?dO�/�O�O �O�O�?�O�O__*_ MON_�Or_�_�_�_�_ 	OO-O�_A_&ouOJo \ono�o�o=o�o�o�o �oo�o4FXj |�_�_�_o�7o ��0�B�T�#x��� �������e����� ,�>�����ŏ�� �Ο������:� L�^�p�����'���ʯ ܯ� �O�a�s����� l���������ƿؿ�� ��� �2�D�g��z� �Ϟϰ����#�5�G� I��}�R�d�v߈ߚ� iϾ��������)߫��<�N�`�r��XST_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��FFF9E3��?�FRS:D�EFAULT�<�FANUC W�eb Server�:
�����<kO�}O�O�O�O�O��WR�_CONFIG ;O�� �?���IDL_CPU_kPC@�B���7P�BHUMIN�(\��<TGNR_I�O������PNP�T_SIM_DO�mVw[TPMOD�NTOLmV �]_�PRTY�X7RTO�LNK 1P�� ��_o!o3oEoWoio>�RMASTElP�|�R�O_CFG�oƙiUO��o�bCY�CLE�o�d@_A�SG 1Q����
 ko,>Pbt ����������sk�bNUM��x��K@�`IPCH�o���`RTRY_C�N@oR��bSCRQN����Q��� �b�`�bR���Տ���$J23_DS/P_EN	���~�OBPROC�ܱU�iJOGP1S�Y@��8�?р!�T�!�?*�PO�SRE�zVKANJI_�`��o_�� ��T�L�6͕����CL_LGP<�_����EYLOGGINʧ`��LA�NGUAGE ,YF7RD w����LG��U�?⧈J�x� �����=P���'0��$� NMC:\RS�CH\00\��L�N_DISP �V��
��������O�C�R.RDzVT=#��K@9�BOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ�{
�Å��ۯ_MOx�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f��xұ]�l��I��p�����������b���3��´  �
`�>����bϸ�z��꜐rg�Jm��
� B߀H�˱]Ӂt�q�	� �p�  P�pQ�p��p|  �Ъ�g���c�	'�� � ��I�� �  �����:�È
���=���"�s���	�ВI  �n @B�cΤ�\��ۤ��tq�y߁rN<���  '������@2��@������/�C��C>�C�@ C���z���
�A���   @�<�P�R�
h�BD�b�A��j�����������Dz۩���������j��(� �� -���C���'�7������q�Y����� �??�ff ��g|y ������q:a��
>+�  PƱj�(�����7	���|�?˙���xZ�p<
�6b<߈;����<�ê<�? <�&Jσ��AI�ɳ+���?offf?I�?&��k�@�.��J<?�`�q�.� �˴fɺ�/��5/� ���j/U/�/y/�/�/ �/�/�/?�/0?q��F�?l??�?/�?+)�?�?�E��� E�I�G+� F��?)O�?9O_O`JO�OnO�Of�BL޳B�?_h�.��O�O�� %_�OL_�?m_�?�__�_�_�_�_�
�h�yÎg>��_�Co�_goRodo�o�GA�ds�q�C�o�o�o|����$]�Hq���D��pC���pCHmZZ7t����6q�q��ܶN'��3A�A�AR�1AO�^?��$�?�K�0���
=ç>�����3�W
=�s#�W��e�צ��@����{�����<���(�B�u���=B0�������	L��H��F�G���G���H�U`E����C�+���I�#�I��H�D�F��E��RC�j=���
I��@H��!H�( E?<YD0q� $��H�3�l�W���{� �������՟���2� �V�A�z���w����� ԯ��������R� =�v�a���������� ��߿��<�'�`�K� ��oρϺϥ������ ��&��J�\�G߀�k� �ߏ��߳�������"� �F�1�j�U��y�� ����������0���T�?�Q����(�1�3�3/E�����5�������q3ǭ8�����q4M�gs&IB+�2D�a���{�^^	����(��uP2P7Q4_A��M0bt��R�����,�/   �/� b/P/�/t/�/ *a)_ 3/�/�/�%1a?��/?;?M?_?q?  �?�/�?�?�?�?O~ 2 F�$�v'Gb�/�A��@�a,�`�qC��C@�o�O�2���OF� D�zH@�� F�P D���O�O�ys<O!_3_E_W_i_s�?���@@pZJ.t22!2~
 p_�_�_ �_	oo-o?oQocouo��o�o�o�o��Q ���+��1��$�MSKCFMAP�  �5� �6�Q�Q"~�c�ONREL  �
q3�bEX_CFENB?w
s�1uXqFNC_QtJOGOVLIM?w�dIpMrd�bKEY�?w�u�bRUN�|�u�bSFSPDTY�avJu3s�SIGN?QtT1�MOT�Nq�b_�CE_GRP 1-p�5s\r��� j�����T��⏙�� ����<��`��U��� M���̟��🧟�&� ݟJ��C���7����� ��گ�������4�V��`TCOM_CF/G 1q}�Vp�􂿔�
P�_ARC�_\r
jyUAP�_CPL��ntNO�CHECK ?{ 	r� �1�C�U�g�yϋϝ� ����������	��({�NO_WAIT_�L�	uM�NTX��r{�[m�_ER�RY�2sy3� A&�������r�cx� ��T_MO��}t��, �,$�|k�3�PARAM��u{��V[���!�u?�� =9@345678901� �&���E�W�3�c������{������� �����=�UM_?RSPACE �V�v��$ODRD�SP���jxOFF�SET_CART�ܿ�DIS��PEN_FILE� �q��c֮�OPTI�ON_IO��PWORK v_�ms �P(�R�Q
�j.j	 �ЖHj&6$� RG�_DSBL  Ċ5Js�\��RI_ENTTO>p9!sC��Pq=#��UT_SIM_D�
r�b� V� LCT ww�bc���U)+$_PEXE�d&RATp �vju��p��2X�j)TU�X)TX�##X d-�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O?O�H2�/oO�O�O�O��O�O�O�O�O_]�< ^O;_M___q_�_�_�_ �_�_�_�_o���X��OU[�o(�꘯(���$o��, ��IpB` �@D�  Ua?��[cAa?��]a]�D�WcUa쪋l;�	l�mb�`�xJ�`�����a�< ��`�� ��b, H(���H3k7HSM�5G�22G���Gp
��
�!�c�'|, CR�	>�>q�GsuaT��3���  �4 spBpyr  ]o�*S�B_����j�]��t�q� ��rna �,����6  ��P�Q�|N��M�,k�!�	'� �� ��I� �  ��%�=��ͭ���ba�	���I  �n @��~����p����� �N �U�[�'!o�:q�pC\�C�@@sBq�|�z�� m�
�A\�*�h@ߐ�n����Z�B\��A���p�G �-�qbz��P��t�_�������( �� -��恊�n�ڥ[A"]Ѻ�b4�'!��(p? �?�ff� ��
����OZ�R���8��z���>΁  	Pia��(�ವ@����ک�a�c�dF#?�嚥�x����<
6�b<߈;܍��<�ê<� <�&�o&�)��A�lcΐI�*�?f7ff?�?&c����@�.uJ<?�`��Yђ^� nd��]e��[g��Gǡd <����1��U�@�y� dߝ߯ߚ����߼�	� ��-������&��"�E�� E��G+� Fþ����� �������&��J�5��bB��AT�8�ђ ��0�6���>���J� n�7��[m�0���h��1��>��M�I
��@��A�[��C�-�)��?�A��� /�YĒ�a�Jp��vav`CH/�������}!@I��Y�'�3A��A�AR1AO��^?�$�?�����±
=���>����3�?W
=�#����+�e��ܒ������{����<�����.(�B�u���=B0������	��*H�F�G����G��H�U�`E���C�+��-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�?O �?3OOWOBOTO�OxO �O�O�O�O�O�O_/_ _S_>_w_b_�_�_�_ �_�_�_�_oo=o(o aoLo�o�o�o�o�o�o �o�o'$]H �l������ �#��G�2�k�V��� z���ŏ���ԏ��� 1��U�g�R���v��� ��ӟ�������-���(�������y�a����Q�<c�,!3�8�}���,!4Mgs����ɢ�IB+կ篴a���{���A�@/�e�S���w��P!�	P�������7��0ӯ�ϑ�R9�K�`��oχϓϥ�  ���χ����)��M� ���������{߉ߛ���ߒߤ�������  )�G�q�_����2 F;�$�&Gb���n�a�[ZjM!C�s��@j/�A�S���F�� Dz��� F�P D��W����)������������x?���@U@
9�E�E���E��
  v������ �*<N`�*�P ���˨�1���$PARAM�_MENU ?�-�� � DEFP�ULSEl	W�AITTMOUT��RCV� �SHELL_W�RK.$CUR_oSTYL�,�OPT�/PTB�./("C�R_DECSN���,y/�/ �/�/�/�/�/?	??�-?V?Q?c?u?�?�U�SE_PROG �%�%�?�?�3C�CR�����7_HOST !�#!�44O�:T̰�?�PCO)ARC�O�;_�TIME�XB� � �GDEBU�GV@��3GINP?_FLMSK�O�IqT`��O�EPGAPe �L��#[CH�O^�HTYPE����?�?�_�_�_�_�_ oo'o9obo]ooo�o �o�o�o�o�o�o�o :5GY�}�� �������1��Z��EWORD ?}	7]	RS`�_	PNS�$斂JOE!>�TE�s@WVTRACEC�TL 1x-�� ��e ���Ӱ��ɆD/T Qy-��䀿D � ��7ӱ4�P  :�L :�GP:�D :�@ �:�8�8�	8�
�8�8�8�8��8�8�X@:�8�*8�8�8�8���:�8�8�x�:��8�P�:�d :�8��8���:�
�:�!8�"�8�#8���:�%8�&�8�'8�(8�)8�*�8���:�,8�-8�.*8�/8�08�18�,� >�P�b�t��������� Ο�����(�:�L� ^�p���������L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�(�p��������� ������ $6H Zl~����� �� 2DVh z������� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_d��_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п�_��� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p�������� //$)�$�PGTRACEL�EN  #!  ��" ��8&_UP z/���g!o S!�h 8!_CFG7 {g%Q#"!�x!�$J �#|"DEFSPD |�,�!!J �8 IN~ TRL }�-�" 8�%�!PE__CONFI� ~g%��g!�$\�%�$LID�#�-�74GRP 1��7Q!�#!A ����&ff"!A�+33D�� D�]� CÀ A)@+6�!�" d�$�9��9*1*0� 	 �+9�(�&�"�? ��	C�?�;B@3AO��?OIO3OmO"!>�?T?�
5�O�O��N�O =��=#�
�O_�O_J_ 5_n_Y_�O}_�_y_�_<�_�_  Dzco" 
oBo�_Roxoco �o�o�o�o�o�o�o�>)bM��;�
V7.10be�ta1�$  �A�E�rӻ�A " �p?!G���q>���r�܁0�q�ͻqBQ��qA\�p�q�4T�q�p�"�BȔ 2�D�V�h�w��p�?�?)2{ȏw�׏ ���4��1�j�U��� y�����֟������ 0��T�?�x�c����� ��ү����!o�,�ۯ P�;�M���q�����ο ���ݿ�(��L�7��p�+9��sF@  �ɣͷϥ�g%����� �+�!6I�[߆����� �ߵߠ���������!� �E�0�B�{�f��� ����������A� ,�e�P���t������� �����=(a L^������ �'9$]�Ϛ� �ϖ�������/ <�5/`�r߄ߖߏ/> �/�/�/�/�/?�/1? ?U?@?R?�?v?�?�? �?�?�?�?O-OOQO <OuO`O�O�O�O�O�� �O_�O)__M_8_q_ \_n_�_�_�_�_�_�_ o�_7oIot���o �o���o�o�o(/! L/^/p/�/{*o�� �������A� ,�e�P�b��������� �Ώ��+�=�(�a� L���p������Oߟ� ��� �9�$�]�H��� l�~�����ۯƯ��� #�No`oro�on��o�o �o�oԿ���8J \ng����vϯϚ� ������	���-��Q� <�u�`�r߫ߖ��ߺ� ������;�M�8�q� \��������z���� ��%��I�4�m�X��� |�����������:� L�^���Z������� ����$�6�H� Swb���� ���//=/(/a/ L/�/p/�/�/�/�/�/ ?�/'??K?]?H?�? ��?�?f?�?�?�?O �?5O OYODO}OhO�O �O�O�O�O�O&8J 4_F_����_�_� �_�_"4-o�O*o coNo�oro�o�o�o�o �o�o)M8q \������� ��7�"�[�m��?�� ��R�Ǐ���֏�!� �E�0�i�T���x��� �����_$_V_ �2��l_~_�_�����R�$�PLID_KNO�W_M  �T������SoV ��U͠�U��
�� .�ǟR�=�O�����m�ӣM_GRP 1���!`0u��T@Rٰo�ҵ�
�� �Pзj��`���!� J�_�W�i�{ύϟϱ����������߱�MR������T��s�w� s��ߠ޴߯߅��� �߻�����A���'� ���������� ����=���#����������}������S��S�T��1 1��U�# ���0�_ A .��,>Pb� �������3 (iL^p��P���2*N���<-/3/)/;/M/4f/x/�/�/5�/�/�/�/A6??(?:?7S?e?w?�?8�?�?�?��?MAD  �d#`PAR�NUM  �w�%OSCH?J �ME
�G`A�Iͣ�EUPD`OrE
a�OT_CMP_��B@�P�@'˥TER_wCHK'U��˪?R$_6[RSl�¯��G_MOA@�_�U_�_~RE_RES_G ��>�oo8o+o \oOo�oso�o�o�o�o��o�o�o�W �\ �_%�Ue Baf�S � ����S0�� ��SR0��#��S�0 >�]�b��S�0}������RV 1�����rB�@c]��t�(�@c\����D�@c[�$���RT?HR_INRl�DA���˥d,�MASS69� ZM�MN8�k��MON_QUEUE ���˦��x�� RDNPUbQN8{�P[��END���_�ڙEXE�ڕ�@B�E�ʟ��OPTI�OǗ�[��PROG�RAM %��%���ۏ�O��TAS�K_IAD0�OCFG ���tO��Š�DATA���Ϋ@��27�>�P�b� t���,�����ɿۿ������#�5�G���IN+FOUӌ������ �ϭϿ��������� +�=�O�a�s߅ߗߩ߀���������^�jč�� yġ?PDI�T �ίc���W�ERFL
��
RGADJ �n�A����?����@�~��IORITY{��QV���MPDSP(H�����Uz����oOTOEy�1�R� (!AF4��E�P]���!t�cph���!u�d��!icm���ݏ6�XY_ȡ�R��ۡ)� a*+/ ۠� W:F�j��� ���%7[�B�*��POR�T#�BC۠�����_CARTRE�P
�R� SKSTyAz��ZSSAV����n�	2500H863���r�$�!�R�����q�n�}/�/�'� UR�GE�B��rYWFF� DO{�rUVWV���$�A�WRUP_�DELAY �|R��$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?�3AQSKIP!�vn�l#x 	1/ +O+ OROdOvO9Hn� �O�G�O�O�O�O�O_ �O_D_V_h_._�_z_ �_�_�_�_�_
o�_.o @oRoovodo�o�o�o �o�o�o�o*<�Lr`���n��?$RCVTM������pDCR!��LЈqC`N��C���C�Q�?��>r���<|�{4M�g��&��/��Z���t����l4�{�4Oi��O� <
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E0�kATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960�iW+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�MD�$bR  ��ϰ�P{_�P_INTVAL�@�����JR_OPT�ION�V �E�BpVAT_GRPw 2����G(y_Ho �e_ vo�o�oYo�o�o�o�o �o*<�bOoND pw������ 	���?�Q�c�u��� ��/���ϏᏣ���� )�;���_�q������� ��O�ɟ���՟7� I�[�m�/�������ǯ ٯ믁��!�3���C� i�{���O���ÿտ� ��ϡ�/�A�S�e�'� �ϛϭ�oρ������ �+�=���a�s߅�G� �߻����ߡ���'� 9�K�]��߁���� y����������5�G��Y��E�$SCAN�_TIM�AYue�w�R �(�#�((�<0.aWaPaP
T�q>��Q��o������OO"2/���d;2"BaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>HE�̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:L!`O�UT",REC 1�Z� d �  	  	������

 �Z�{0 H6lZ�~�� ���� //D/2/ h/z/\/�/�/�/�/�/ �/�/?�/,?R?@?v? d?�?�?�?�?�?�?�? OO(ONO<OrOTOfO �O�O�O�O�O�O_&_ _J_8_Z_\_n_�_�_ �_�_�_�_�_"ooFo 4oVo|o^o�o�o�o�o �o�o�o0TB xf����(� ��,��P�>�`��� h���������Ώ�� (�:��^�L���p��� ����ܟ���� �6� $�Z�H�~���r����� دƯ����2��&� h�V���z�����Կ� ȿ
�����.�d�R� �Ϛ�|ϾϬ������ ���<��`�N�pߖ� �ߺߨ���������8�&�\�J�l��jV� 1�w Pl��	� � ��F��
TYPE�VFZN_CF�G �x��d7�GRP� 1�A�c ,�B� A� D;�� B���  B�4RB21^HELL:�(
 X����%RSR���� E0iT�x�� ����/S�ew�  ���%w������#�����A�2#�d�����HK 1���  ���m/h/z/�/�/�/ �/�/�/�/
??E?@?�R?d?�?�?�?�?��OMM ����?���FTOV_ENB� ���+�HOW_R�EG_UIO��I_MWAITB�.JKOUT;F��LIwTIM;E���O�VAL[OMC_UN�ITC�F+�MON�_ALIAS ?�e�9 ( he �s_(_:_L_^_��_ �_�_�_�_j_�_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]n��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� ���������ӟ~��� 	��-�?��c�u��� ����V�ϯ����� �;�M�_�q������ ��˿ݿ����%�7� I���m�ϑϣϵ�`� ������ߺ�3�E�W� i�{�&ߟ߱������� ����/�A�S���w� ����X������� ���=�O�a�s���0� ������������' 9K]���� b���#�G Yk}�:��� ���/1/C/U/ / f/�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_O
O�O�O�O �O�OvO�O__%_7_��C�$SMON_�DEFPRO ����`Q� *SY�STEM*  d�=OURECAL�L ?}`Y (� �}.xcop�y fr:\*.�* virt:\tmpback�Q�=>inspir�on:1228 ��R�_�_�_	o  }/�Ua�_�_�P�_ao�so�od
xyzrate 61 +o@=oOo�o�oe�g>�X4064 �o�o ]o��o�b+=O����)y207�6��\�n���i3��Ts:orderfil.dat�l@*�ӏ���	�`*�Rmdb:�o*�ˏ\� n���i�_�o.�O��� ��o����7�Пa� s�������3�N�߯� ��(�:�̯]�o��� ����9�ʟۿ���� $���H�Y�k�}ϐ��� ��Ư������� ���`D�U�g�yߋ�}6����emp��192�.168.4��4?6:3892��������}.��*.d�������`�r��1 +�=�O������� ���2 ����c��u����4 �:prwgst�`.dg����U�����
�ť�c?onslog����� ��ew�	io���<N���2���errall.ls����fx� }9�߲�=S���/}0 ߻���b/t/�/�߫9R 8736 W/�/�/�/ �/�)�/`?r?�?�� ��;?M?�?�?O�'� �4�?�?cOuO�O�� 5/�'�O�O�O/"/�O �(�Ob_t_�_����3̆=_6 U_�_�_
o }5 ϱ_�_�_goyo �o�O�O9_T_�o�o	 _�o@_�ocu��_ -o?o�_���o� �No_�q����o�o1 �oݏ��&��J�[�m�����$SN�PX_ASG 1ߺ������� P 0 �'%R[1�]@1.1����?���%֟��&�	� �\�?�f���u����� ���ϯ��"��F�)� ;�|�_�������ֿ�� ˿���B�%�f�I� [Ϝ�Ϧ��ϵ����� ��,��6�b�E߆�i� {߼ߟ���������� �L�/�V��e��� ����������6�� +�l�O�v��������� ������2V9 K�o����� ��&R5vY k�����/� �<//F/r/U/�/y/ �/�/�/�/?�/&?	? ?\???f?�?u?�?�? �?�?�?�?"OOFO)O ;O|O_O�O�O�O�O�O �O_�O_B_%_f_I_ [_�__�_�_�_�_�_ �_,oo6oboEo�oio {o�o�o�o�o�o�o L/V�e�� ������6���+�l�O�v�������PARAM ������ �	���P����O�FT_KB_CF�G  ヱ���P�IN_SIM  ���C�U�g������RVQSTP_DSB,�򂣟�����SR �/��� & MULT�IROBOTTA�SK�����T�OP_ON_ER/R  ����PTN /��@�A	�RI�NG_PRM� ���VDT_GR�P 1�ˉ�  	������������ Я�����*�Q�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߣ� �߲����������� 0�B�i�f�x���� ���������/�,�>� P�b�t����������� ����(:L^ p�������  $6HZ�~ �������/  /G/D/V/h/z/�/�/ �/�/�/�/?
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8___\_���VPRG_COUNT��@���R'ENBU��UM�S���__UPD 1�>/�8  
s_� oo*oSoNo`oro�o �o�o�o�o�o�o+ &8Jsn��� ������"�K� F�X�j���������ۏ ֏���#��0�B�k� f�x���������ҟ�� ����C�>�P�b��� ������ӯί������UYSDEBU)G�P�P�)�d�YH�SP_PASS�U�B?Z�LOG [��U�S)�9#�0�  ��Q)�?
MC:\��6���_MPC���U�$��Qñ8� �Q趿SAV ���ج�ǲ&�ηSV�;�TEM_TIM�E 1��[ (�m��&����}YT1SVGUNS�P֕U'�U���AS�K_OPTIONДP�U�Q�Q��BC?CFG ��[u�� n�A�a�` a�gZo��߃ߕ��߹� ������:�%�^�p� [��������� � ����6�!�Z�E�~�i� ��������&����� ��&8��nY� }�?��ԫ � �(L:p^� ������/ / 6/$/F/l/Z/�/~/�/ �/�/�/�/�/�/2?8  F?X?v?�?�??�? �?�?�?�?O*O<O
O `ONO�OrO�O�O�O�O �O_�O&__J_8_n_ \_~_�_�_�_�_�_�_ o�_ o"o4ojoXo�o D?�o�o�o�o�oxo .TBx��j �������� ,�b�P���t�����Ώ ��ޏ��(��L�:� p�^�������ʟ��� �o��6�H�Z�؟~� l�������د���ʯ  ��D�2�h�V�x�z� ��¿���Կ
���.� �>�d�Rψ�vϬϚ� �Ͼ�������*��N� �f�xߖߨߺ�8��� ������8�J�\�*� ��n���������� ��"��F�4�j�X��� |������������� 0@BT�x� d�����> ,Ntb���� ��/�(//8/:/ L/�/p/�/�/�/�/�/ �/�/$??H?6?l?Z? �?~?�?�?�?�?�?O �&O8OVOhOzO�?�O �O�O�O�O�O
__�O @_._d_R_�_v_�_�_ �_�_�_o�_*ooNo <o^o�oro�o�o�o�o �o�o J8n $O�����X����4�"�X�B�v���$TBCSG_G�RP 2�B��  �v�� 
 ?�   ������׏�������@1��U�g�z���ƈ��d, ���?~v�	 HC��d��>����e�CL  B���Пܘ��w���\)���Y  A�ܟ$�B�g�B�Bl�i�X��ɼ���X��  DA	J���r�����C�����үܬ���D�@ v�=�W�j�}�H�Z����ſ���������v�	V3.0�0��	m61c�	*X�P�u�g�&p�>���v�(:��� ��p͟�  O����p�����z�JCFG �B���� �����������=��=�c�q�K�qߗ߂� �ߦ��������'�� $�]�H��l����� ��������#��G�2� k�V���z��������� �����p*<N ���l����� ��#5GY} h����v�b�� >�// /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?d?R?t?v?�? �?�?�?�?O�?*OO :O`ONO�OrO�O�O� �O�O�O_&__J_8_ n_\_�_�_�_�_�_�_ �_�_�_oFo4ojo|o �o�oZo�o�o�o�o�o �oB0fT�x �������,� �P�>�`�b�t����� Ώ�������&�L� �Od�v���2�����ȟ ʟܟ� �6�$�Z�l� ~���N�����دƯ� � �2��B�h�V��� z�����Կ¿���� .��R�@�v�dϚψ� ���Ͼ�������<� *�L�N�`ߖ߄ߺߨ� ���ߚ�������\� J��n������� ���"���2�X�F�|� j��������������� .TBxf� ������ >,bP�t�� ���/�(//8/ :/L/�/�ߚ/�/�/h/ �/�/�/$??H?6?l? Z?�?�?�?�?�?�?�? O�?ODOVOhO"O4O �O�O�O�O�O�O
_�O _@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<oro`o�o�o�o�o �o�o�o&�/>P �/������ ���4�F�X��(� ��|�����֏���� Ə0��@�B�T���x� ����ҟ������,� �P�>�t�b������� ��������:�(� ^�L�n�������2d �����̿�$�Z�H� ~�lϢϐ��������� �� ��0�2�D�zߌ� �߰�j���������� 
�,�.�@�v�d��� �����������<� *�`�N���r������� ������&J\ �t��B��� ���F4j| ��^����/��  2 6# �6&J/6"�$TB�JOP_GRP �2���?  ?�X,i#��p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�x�'�!�!>���
5�59>�0+1�33=�CL� �fff?+0?�ffB� J1�%Y?d7�.���/>��2�\)?0�5����;��hCY� ��  @� �!B� � A�P?�?�3EC�  D�!�,�0�*BOߦ?�3JB���
:���Bl�0��0�$�1�?O6!?Aə�AДC�1sD�G6�=q�E�6O0�p��B�Q�;�A�� �ٙ�@L3D	��@�@__�O�O>BÏ\JU�OHH�1ts}�A@33@?1� C�� �@�_�_&_8_>��D�UV_0��LP�Q30<{�zR� @�0�V�P!o3o �_<oRifoPo^o�o�o �oRo�o�o�o�oM (�ol�p~���p4�6&�q5	�V3.00�#m761c�$*(��$�1!6�A� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,IR�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^S@;Q��|8�E`rz@/&�8�6&�<��1�w�^$ES�TPARS  �*({ _#HR��AB_LE 1�p+Z�6#|�Q� � 1�|��|�|�5'=!|�	�|�
|�|�˕6!�|�|�|���RDI��z!ʟܟ� ��$���O������ ¯ԯ�����S��x# V���˿ݿ��� %�7�I�[�m�ϑϣ� �����������U-�� ��ĜP�9�K�]�o���-�?�Q�c�u���6�N�UM  �*z!� >  Ȑ�����_CFG ������!@b IMEBF_TT����x#��a�VER��b�w�a�R 1�p+
' (3�6"1 ��  6!����������  �9�$�:�H�Z�l�~� ���������������^$��_��@x�
�b MI_CHAN�m� x� kDBGLV;0o�x�a!n �ETHERAD �?�� �y��$"�\&n ROUmT��!p*!�*�SNMASK��x#�255.�h�fx^$OOL�OFS_DI���[ՠ	ORQCTRL �p+;/�� �/+/=/O/a/s/�/ �/�/�/�/��/�/�/�!?��PE_DET�AI��PON_�SVOFF�33P_MON �H��v�2-9STRTC_HK ����42VTCOMPA�Ta8�24:0FPR�OG %�%�MULTIROB�OTTO!O06�P�LAY��L:_IN�ST_MP GL�7YDUS���?�2L�CK�LPKQUIC�KMEt �O�2SC�RE�@�
tps��2�A�@�I���@_Y���9�	S�R_GRP 1Ҿ� ��� \�l_zZg_�_�_�_�_�_�^�^�oj�Q'O Do/ohoSe��oo�o �o�o�o�o�o! WE{i�������	1234�567��!���X��E1�V[
 �}�ipnl/a�g?en.htmno���������ȏ~�P�anel setup̌}�?��0�B�T�f� ��񏞟 ��ԟ���o���� @�R�d�v������#� Я�����*���ϯ ůr���������̿C� �g��&�8�J�\�n� ����϶��������� uϣϙ�F�X�j�|ߎ� �����;��������0�B��*NUALR�Mb@G ?�� [���������� �� ��%�C�I�z�m�������v�SEV � ����t�E?CFG Ձ=]�/BaA$   B�/D
 ��/C� Wi{�����@�� PRց;C �To\o�I�6?K0(%����0 �����//;/ &/L/q/\/�/�/�/lƇD �Q�/I_��@HIST 1׾�9  (�0� ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1 Ec0p?0�?�?�?/C�'=?O>71n?�?	OO-O�1y3�?O5edit[2?MULTIRf?O��O�O2O� FOP=962vO __$_6_�O�O�A36�O�_�_�_ �_IR�_�_�_oo+o =o�_aoso�o�o�o�o Jo�o�o'9I|��a81�ou��� ���o���)�;� M��q���������ˏ Z�l���%�7�I�[� ��������ǟٟh� ���!�3�E�W���� ������ïկ�v�� �/�A�S�e�Pb�� ����ѿ������+� =�O�a�s�ϗϩϻ� ������ߒ�'�9�K� ]�o߁�ߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y��� v�����������	 �?Qcu��( ����)� M_q���6� ��//%/�I/[/ m//�/�/�/D/�/�/ �/?!?3?�/W?i?{? �?�?�?�����?�?O O/OAOD?eOwO�O�O �O�ONO`O�O__+_ =_O_�Os_�_�_�_�_ �_\_�_oo'o9oKo �_�_�o�o�o�o�o�o jo�o#5GY�o�}������?���$UI_PAN�EDATA 1������  	�}��0�B�T�f�x��� ) �����4�ۏ���� #�5���Y�@�}���v� ����ן�������1���U�g�N������ �1��Ïȯگ� ���"�u�F���X�|� ������Ŀֿ=���� ��0�T�;�x�_Ϝ� �ϕ��Ϲ������,���M��j�o߁ߓ� �߷������`��#� 5�G�Y�k��ߏ��� �����������C� *�g�y�`��������� F�X�	-?Qc ����߫���� ~;"_F� �|�����/ �7/I/0/m/�����/ �/�/�/�/�/P/!?3? �W?i?{?�?�?�?? �?�?�?O�?/OOSO eOLO�OpO�O�O�O�O �O_z/�/J?O_a_s_ �_�_�_�O�_@?�_o o'o9oKo�_oo�oho �o�o�o�o�o�o�o# 
GY@}d�� &_8_����1�C� �g��_��������ӏ ���^���?�&�c� u�\�������ϟ��� ڟ�)��M����� ������˯ݯ0��� ��7�I�[�m������ ����ٿ�ҿ���3� E�,�i�Pύϟφ���0����Z�l�}���1� C�U�g�yߋ�)߰� #������� ��$�6� ��Z�A�~�e�w��� ��������2��V��h�O����v�p��$�UI_PANEL�INK 1�v��  ��  ��}12�34567890 ����	-?G� ��o�����a ��#5G�	�����p&���   R�����Z� �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?.O@O ROdOvO�O O�O�O�O �O�O_�O�O<_N_`_0r_�_�_�0,���_ ��_�_�_ o2ooVo hoKo�ooo�o�o�o�o �o�o��,>r} ��������� ���/�A�S�e�w� �������я���t v�z����=�O�a� s�������0S��ӟ� ��	��-���Q�c�u� ������:�ϯ��� �)���M�_�q����� ����H�ݿ���%� 7�ƿ[�m�ϑϣϵ� D��������!�3�E� �_i�{�
�߂����� �������/��S�e� H���~��R~'�'� a��:�L�^�p��� ������������  ��6HZl~�� �#�5��� 2 D��hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?�/ �?�?�?�?�?�?m?O O&O8OJO\O�?�O�O �O�O�O�O�O[�_�� 4_F_)_j_|___�_�_ �_�_�_�_o�_0oo Tofo��o��o��o �o�o,>1b t����K�� ��(�:����{O ������ʏ܏�uO� $�6�H�Z�l������� ��Ɵ؟����� �2� D�V�h�z�	�����¯ ԯ������.�@�R� d�v��������п� ��ϕ�*�<�N�`�r� ���O�Ϻ�Io������ ���8�J�-�n߀�c� �߇����߽����o 1�oX��o|���� ���������0�B� T�f������������ ��S�e�w�,>Pb t��'���� �:L^p� �#���� // $/�H/Z/l/~/�/�/ 1/�/�/�/�/? ?�/ D?V?h?z?�?�?�??? �?�?�?
OO.O��RO dO�߈OkO�O�O�O�O �O�O_�O<_N_1_r_ �_g_�_7OM�m��$UI_QUI�CKMEN  >��_Ao�bRESTORE� 1�?  �|��Rto�o�im�o�o�o�o �o:L^p� %������o� ���Z�l�~����� E�Ə؏���� �Ï D�V�h�z���7����� ��/���
��.�@�� d�v�������O�Я� ����ßͯ7�I��� m�������̿޿��� �&�8�J��nπϒ� �϶�a�������Y�"� 4�F�X�j�ߎߠ߲� �����ߋ���0�B�T�gSCRE`?�#mu1s]co`u2��3��U4��5��6��7��y8��bUSERq�dv��Tp���ks����4��5��6��7���8��`NDO_�CFG �#k � n` `PDA�TE ����NonebSE�UFRAME  ��TA�n�RTO?L_ABRTy�l�Α�ENB����GR�P 1�ci/aCz  A�����Q@�� $6HR�d��`U�����MSK  �����MNv�%�U�%����bVISCAN�D_MAX�I���FAIL_�IMG� �PݗP#���IMREGN�UM�
,[SI�Z�n`�A�,~VONTMOU��@���2���a��a��~��FR:\� � MC{:\�\LOG�7B@F� !�'/�!+/O/�Uz �MCV�8#U�D1r&EX{+�S|�PPO64_���0'fn6PO��LIb�*�#9V���,f@�'�/�� =	�(SZV��.����'WAI��/STAT 	����P@/�?�?�:�$�?�?��2DW�P  ��P yG@+b=��� H��O_JMPE�RR 1�#k
 � �2345678901dF�ψO{O �O�O�O�O�O_�O*_�_N_A_S_�_
� M�LOWc>
 �_�TI�=�'M�PHASE  ���F��PSHI[FT�1 9�]@<�\�Do�U#oIo �oYoko�o�o�o�o�o �o�o6lCU �y����� �@�	�V�-�e2����	VSFT1�2�	VM�� ��5�1G� ���%A_�  B8̀̀E�@ pكӁ˂�у���z�ME@�?��{��!c>&%�aM�1��k�0�{ �$�`0TDINEND��\�O� �z���S��w��P��=�ϜRELE�Q���Y���\�_ACT�IV��:�R�A ���e���e�:�R�D� ���YBOX� �9�د�6���02���1�90.0.�83v��254�:�QF�	 �X��j��1�ro�bot���  � p�૿�5pc��̿������7�����-�f�ZABC�����,]@U��2 ʿ�eϢωϛϭϿ� ���� ���V�=�zߐa�s߰�E�Z��1� Ѧ