��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�FPCUR�EQ1 � �$SOFT; T_�ID�TOTAL7_EQ� $� � �NO�PS_SP�I_INDE���$�X�SCRE�EN_NAME ��SIGN���� PK_�FIL	$TH{KYMPANE��  	$DUM?MY12 � u�3|4|GRG_�STR1 � �$TITP$I��1�{�P����5�6�U7�8�9�0���z�����1��1�1 '1
'2�"GSBN_CF�G1  8 �$CNV_JNT�_* |$DAT�A_CMNT�!?$FLAGS�*�CHECK�!�A�T_CELLSE�TUP  P� $HOME_�IO,G�%�#M�ACRO�"REPyR�(-DRUN� 5D|3SM5H �UTOBACKU�0 $E�NAB��!EVI�C�TI �� D� DX!2ST�� ?0B�#$INT�ERVAL!2DISP_UNIT!2�0_DOn6ERR��9FR_F!2I�N,GRES�!�0Q_;3!4C_W�A�471�:OFF_� N�3DELHL�OGn25Aa2?1i1@N?�� -JM�H W+0�$Y �$DB� 6CO5MW!2MO� 21�\D.	 \rVE�1$F��A{�$O��D�B�CT_MP1_F�E2�GC1_�3�B�2FX�D�#
 d �$CARD_EX�IST4$FS?SB_TYPuA?HKBD_S�B�1�AGN Gn �$SLOT_NUyMJQPREV,D�BU� g1G ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�AE�TE_OKRUSބP_CRQ$�;4�V� 0LACIw1�RAPk �1x@�ME@$D��V�Q�Pv�A{'o�BL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa�!ip;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I�9�TY�D,P*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6���7��8��9�CO�$ <� $6x8K3 1w`O_M�@�C_ t � E#f6NGP�ABA�  �c��ZQ���`���@n!r��� ��P�0��,��x�p�PzP�b26����"J�_)R��BC�J��3�JVP��tBS��}�Aw��"�tP_*0O�FSzR @� RcO_K8���aIT�3���NOM_�0�1�ĥ34 ��T Ԑ� $���AxP��K}EX�� �0g0I01��p��
$TFa��C$7MD3��TO�3�0yU� �� �)Hw2�C1|�EΡg0�wE{vF�vF����p@�a2 
P�$A`PU�3Nc)#�dR*�AX�!�sDETAI�3BU�FV��p@1 |X�p۶�pPIdT� +PP[�MZ�Mg�Ͱ�j�F[�SIMQS@I�"0��A.�����Nlw Tp|zM�x�P�B�FACTrbHPEW7�P1Ӡ��v��MCd� �$*1JB�p<�*1GDECHښ�H����b� � +PN�S_EMP��$GP���,P_��3�p2�@Pܤ��TC��|r ��0�s��b�0�� �B0���!
���JR� ��_SEGFR��Iv *�aR�TkpN&S,��PVF4��� &k�Bv�u�cu� �aE�� !2��+�MQ��E�SIZ�3�����T��P�����aRSINF�����kq�� ������LX������F�CRCMu�3CClpG��p���O}�� �b�1�������2�V�DxIC��C���r��`��P��{� EV ��zF_��F�pNB0�?������A�! �r�Rx�� ��V�lp�2��aR�t��,�g�RTx #�5�5"2��uA�R���`CX�$LG�p��B�1 `s�P�tB�aA�0{�У+0R���tME�`!BupCfrRA 3tAZ��h��pc�OT�FC�b�`�`FNp���1��ADI+�a%��b �{��p$�pSp�c�`aS�P��a,QMP6䒁`Y�3��M'�pUt��aU  $>�TITO1�S�S�!���$�"0�DBPX�WO��!��$cSK��2p�DB��"�"@�PR8�� 
� ���# �>�q1$��$��+�L9$?(�V�R%@?R4C&_?�R4ENE��'�~?(�� RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@����C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!��DCS_)  `IS#� �� @�s3S�AQ汯 4R�x�ZSW�AQ�p�@1UW���cTNTV)�5RV 
a���|c�éWƃ���JB��x0��SAF�Eۥ�V_SV�bEOXCLUU�;��'ONL��cYg�~a�z�OT�a{�HI_�V? ��R, M�_ #*�0� ��_z�2�o CdSGO  +�rƐm@�A�c ~b���w@��V�i�b>�fANNUNx0�$��dIDY�UABc �@Sp�i�a+ �j�f�"��pOGIx2,��c$F�b�$ѐOT�@�A $DUM�MY��Ft��Ft±�� 6U- ` !�HE�|s��~bc|�B@ SUFFI��[4PCA�Gs�5Cw6CqibMSW�U. 8!�KEYI��5�TM�1�s�qLoA�vINޱw�(�!�, / D��HOST�P!4���<����<�°<��p<�EMp'���Z�� SBL� �UL��0   �	��E�� T�0?1 � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0�QS�����#��SAV �����c�S< 9�`��fP$�0E!� YwN_B�#2 0�`DI�d�pO|�m��#�$F�R_IC�� �ENC2_Sd3  ��< 3�9���� cgp����B4�"��2�A��ޖ5���`ǻ��@Q@K&D-!�a�A�VER�q����D3SP
���PC_�q���"�|�ܣ�VALMU3�HE�(�M�sIP)���OPPm �TH�*���S" T�/�Fb�;�d����d D�qЗ1�6 H(rLL_DUǀ�a�@��k���֠OT�"U�/����@@NOAUTO70�$}�x�~�R@s��|�C͠��IC� 2z�L�� 8H *��L� ���Բ@sv��` � �� ÿ���Xq��cq����q���q��7��8J��9��0���1�U1 �1-�1:�1G�U1T�1a�1n�2|ʩ2��2 �2-�2�:�2G�2T�2a�2*n�3|�3�3� �U3-�3:�3G�3T��3a�3n�4|'�����9 < ���z�ΓKI����H硵BaFEq@{@�: ,��&a? P_P?��>�����E�@���!QQ��z;fp$TP�?$VARI����n,�UP2Q`< W�߃TD��g���`��x�����_BAC�"G= T2����$)�,p+r³�p IFI�� �p�� q M�P"��Fl@``>t �;��6����ST ����T��M ����0	��i���F����������kRt ����FO�RCEUP�b܂FWLUS
pH(N��x� ��6bD_CM�@E�7N� (�v�P.��REM� Fa@��@j���
K�	9N���EFF/��f�@IN�QOV���OVA�	TRO�V DT)��DTMX:e �P:�/��Pq�vXpCLN _�p��@ ��	_|��_T: �|��&PA�QDI����1��0�Y0R�Qm�_+qH���M����CL�d#�RIqV{�ϓN"EAR/�IO�PCP��BR��CM�@N 1b{ 3GCLF���!DY�(��a�#5T�DG���� �%�%�FSS� )�? �P(q1�1�`_(1"811�EC1�3D;5D6�GRA����@�����PW��ON2EBU�G�S�2�C`gϐ_?E A ��?�����TERM�5B<�5��ORIw�0�C�6 �SM_�-`���0D�5����TA�9E�5����UP��F� -�QϒA�P�3�@B�$SEGGJ� EL��UUSEPNFI��pBx��1@��4>D�C$UF�P��!$���Q�@C���G�0T�����SNST�j�PATۡg��AP'THJ�A�E*�Z% qB\`F�{E��F�q�pA�RxPY�aSHFT�͢qA�AX_SHOQR$�>��6 @$GrqPE���OVR����aZPI@P@$U?r *aAYLO���j��I�"��Aؠ��ؠERV��Qi�[Y)��G��@R��i�e��i�Rz�!P�uASYM����uqAWJ�G)��E ��Q7i�RD�U[d�@ i�U��C�%UP���P����WOR�@M��]k0SMT��G��cGR��3�aPA�@���p5�'�H � uj�A�TOCjA�7pP]Pp$OP@d�O��C�%�p�YO!��RE.pR�Cb�AO�?��Be5p�R�EruIx'QG�e$7PWR) IMdu�R�R_$s��5��B �Iz2H8�=�_AD�DRH�H_LENAG�B�q�q:�x�R��So�J.�SS��SK������ ��-ãSE*���rSN�M-N1K	�j�5�@r�֣OL��\�WpxW�Q�>pACRO�p ���@H ����Q� N��OUPW3�b_>�I��!q�a1����� ���|��������`-���:���iIOX2S=�D�e��]���L $��p�!_�OFF[r_�PRM�_�I�aTTPu_�H��M (�p�OBJ�"�pG�$�H�LE�C��ٰN� � 9�*�AB%_�T��
�S�`�S6��LV��KRW"du�HITCOU?B-Gi�LO�q�����d� Fpk�GpSS� ���HWh�wA���O.��`INCP}UX2VISIO�� !��¢.�á<�á-¿ �IOLN)�P� 87�R'�[p$�SL�bd PUTM_��$dp�Pz x�� F_AS2Q/�$LD���D�DaQT U�0]P�A������PHYG灱Z�̫P4�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp���x�X�ٶ��UJ��S��v��NE�WJOG�GN �DIS��r�KĠL��3T |��AV���`_�CTR!S^�FgLAGf2r�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_H��Dq��N?���V��EE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�B�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S S�n���_BUFF�1XY��PT�$�� �v��fĘ�1�A�rYY��P ���\��pOS1�2��3���0Z �  ��aiE�*���IDX�dP�RhrO��+��A&ST��R���Yz�<! Y$EK&CK+���Z&�m&�5�0[ L ��o�0��]PL�6pwq��t^����w��7�_ \ �`��瀰��7��#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3b�DM�R7��LDR5<4R5ORG.���e2 (`���V�8.��T<�4�d^ �q�<4��-4
R5S�`T00m��0D}FRCLMC!D`�?�?3I@��MIC���d_ d���RQzm�q�DSTB	��  �Fg�HAX�;b �H�LEXC#ESZr��rBMup�a`��B;d�!rB`�j�`a��F_A�J���$[�O�H0K�db� \��ӂS�$MB既LIБ}SREQUIR�R>q�\Á�XODEBU��oAL� MP�c�ba��P؃ӂ!BoAND���`�`ad�҆�c�cDC1��IN�����`@�(hB?Nz�@q��o��UwPST8� e�r7LOC�RI�p�EX�fA�p��AoA�ODAQP�f Xf��ON��[rMF�� ���f)�"I��%�e���T� �FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y��RFЭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?:�uD�)P:�`��	@Ði �@CU���V�T0�eRR2�j Dɐ�Qނ�B?d$CALI�@F��G�s�2�RINt��v�<��NTE���kE���,��b����_Nl��ڂ��kDtׄRm�DIViF�DH�@ـn�c$V��'c!$��$Z�����~��[��oH ��$BELTb��!A/CCEL+��ҡ��IRC�t����yT/!��$PS�@
#2L�q�Ɣ83��𧗙�� ��PATH��������3̒Vp�A�_�Q�.�4�B�C�ᐈ�_MGh�$�DDQ���G�$FWh��p��m�����b��DE��PPABN�ԗROTSPEED����00J�Я8���@���$USE�_��P��s�SYh��c�A >qYNu@9Ag��OFF�q�7MOUN�NGg�K�sOL�H�INC*���a��q��Bj�L@�BENCS��q�Bđ���D��IN#"��x���4�\BݠVEO�w�Ͳ�23_UPE�߳LOWL���00����D���BwP��� ��1RCʀƶMOSIV�JRMO���@GPERCH  �OV��^��i�<! �ZD<!�c��d@�P���V1�#P͑��L`���EW��ĸUP��8����TRKr�"AYLOA'a�� Q�-�̒<�1Ӣ`0 ��RcTI$Qx�0 MO�� �МB R�0J��D��s��H����b�DUM�2(�S_BCKLSH_C̒��>�=� q�#�U��ԑ���2�t�]ACLALvŲ�18n�P�CHK00'%SD�RTY4�k���y�1�q_6#2�_U�M$Pj�Cw�_�SC�L��ƠLMT_J'1_LO��@���q��E�����๕����SPC��7����&��PCo���H� �PdU�m�C/@�"XT_�.c�CN_��N��e�&��SFu���V�&#@����9�̒��=�C�u�SH6#��c����1 �Ѩ�o�0�͑
��_�3PAt�h�_Ps�W�_10��4�R�01D�V�G�J� L�@J�O�GW���TORQU��ON*�Mٙ�sRH�љ��_W��-�_@=��C��I��I��I�II�F�`�J�LA.�1[�VC��0�D(RO1U�@i�B\JRKU��	@?DBL_SMd�B�M%`_DLC�BGRV��C��I���H_� �*CO1S+\�(LN�7+ X>$C�9)I�9)u*�c,)�Z2 HƺM1Y@!�( "TH&-�)�THET0�NK�23I��"=�A CB6CB=�C�A�B(2`61C�616SBC��T25GTS QơC ��aS$" �4c#�7r#$DUD�EX�1@s�t�(R�6��(QQ|rN�f$NE�DpIB �U�\B5��$!��!A��%E(G%(!LP!H$U�2׵�2SXpC c%pCr%�2�&�C�J�&�!�VAHV6H3�YLV�hJVuKV�KV�KV*�KV�KV�IHAHZF�`RXM��wXuKH�KH��KH�KH�KH�IOJ2LOAHO�YWNOhJUOuKO�KO�KO�KO�KO�&F�2#1i�c%�d4GSPBAL�ANCE_�!�cLmEk0H_�%SP���T&�bc&�br&PFULC�hr�grr%Ċ{1ky�UTO_?��jT1T2Cy��2N&�v�ϰctw�g�pP�0Ӓ~���T��O�|��� INSEGv��!�REV�v!���D3IF��1l�w�1m�0OB�q
��Ɠ�MIϰ1��LC�HWAR����AB�&u�$MECH`,1� :�@�U�AX:��P��Y�G$�8pn �
Z��|���ROBFR�CR��N����MSK_�`f�p WP Np_��R����΄ݡ�1��ҰТ`΀ϳ��΀"�IN�q��MTCOM_�C@j�q  �L��p��$NOR�E³5���$�r� 8� GR�E�S�D�0ABF�$XYZ_DA5A���DEBU�qI��Q��s �`$�COD��� ��k�F��f�$BUFIN�DXР����MO�R��t $-�U ��)��r�B���������Gؒu � ?$SIMULT ���~�� ���OBJE|�` �ADJUS>��1�AY_Ik��Dp_����C�_FIF�=�T� ��Ұ�� {��p� �����p�@�ŝD�FRI��ӥT&��RO� ��E���=��OPWO�ŀ�v0��SYSByU�@ʐ$SOP�ȸ��#�U"��pPR�UN�I�PA�DpH�D����_OU��=��qn�$}�I�MAG��ˀ�0Pf�qIM����IN��q���RGOVRDȡ:���|�P~���Р�0L_6p���i��SRB���0��M���EDѐF� ��N�`M*����̰S�L�`ŀw x �$OVSL�vSDI��DEXm�g�eĐ9w�����V� ~�N ���w����Ûǖȳ�M�����q<��� x HˁE�F�ATUS���Cp�0àǒ��BTM��*��If���4����\(�ŀy DˀEz�g���PE�r�����
���EXE��V���E�Y�$Ժ ŀz @�ˁ��UP{�h�$�p��XN���9ԼH� �PG"�{� h $SUB���c�@_��01\�M/PWAI��P���ՓLO��-�F�p��$RCVFAILs_C�-�BWD"�|F���DEFSPup | Lˀ`�D�p� U�UNI���S���R`���_L�pP��̐���ā}��� B�~���|��`:ҲN�`KET��y����P� $�~���0SIZE�ଠ�{���S<�OR��FORMAT/p � XF���rEMR���y�UX���LI�7�ā  $>�P_SWI����@��_PL7�ALO_ �ސR�A���B�(0C��Df��$Eh����C_�=�U� � �c ���~�J3�0�����TIA4��5:��6��MOM������ �B�A�D��*��* PU70NRW��W �@�U����� A$PI�6���	�� )�4l�}69���Q���c�SPEED�PGq�7�D�>D� ���>tMt[��SAM�`痰8>��MOV���$���p�5��5�D�1�$2�������d{�Hip�IN?, {�F(b+=$�H*�(x_$�+�+GAMM�f|�1{�$GET���ĐH�D����
^pL�IBR�ѝI��$HI��_��Ȑ*B6�E��*8A$>G086LW=e6\<G9�686���R��ٰV��$PDCK�Q�H�_����;"��z�.%�7�4*�9� ��$IM_SRO�D�s"���H�"�LE�O�0\H���6@���U� �ŀ��P�qUR_SCR�ӚAZ��S_SA�VE_D�E��NO��CgA�Ҷ��@�$ ����I��	�I� %Z [� ��RX" ��m� ��"�q�'"�8 �Hӱt�W�UpS��рM��O㵐.' }q��Cg���@ʣ�����S�M�AÂ� �� $PY��3$WH`'�NGp��� H`��Fb��Fb��Fb��PLM���	� 0h�H�J{�X��O��z�Z�e8T�M���� pS��C��O__0_B_t�a��_%�� |S� ���@	�v��v �@���w�v��EM��%���dt�B�ː��ftPn��PM��QU� �U�Q��A-�wQTH=�HOL��oQHYS�ES�F,�UE��B��O#��  -�P0�|�gAPQ���ʠu���O��ŀ�ɂv�-�A;ӝGROG��a2D��E�Âv�_�ĀZ�INFO&��+����b�Ȝ�OI킍 ((@SLEQ/�#@������o���S`�c0O�0�01E�Z0NUe�_�AUT<�Ab�COPY���(��{��@M��N������1�P�
� ��RG4I�����X_�Pl�C$�����`�W���P��j@�G���E�XT_CYCtb����p����h�_NA�!$�\�<��RO�`]�� �s m��POR�㸅����SRVt�)l����DI �T_l� ��Ѥ{�ۧ��ۧ �ۧU5٩6٩7٩8��Ҝ�S�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,(@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#qX� �Q�SKIP�� Ĵ��x�O�`NT!���P_x���ǚ@ �b�p1�1�1Ǹ� ?� �?��>��>�&��>�3�>�9�J2�R;쐖 4��EX� TQ����ށ�Q����[�KFд�w�R;DCIf� �U`�X}�R�#%M!*�0��)��$RGEAR_�0IO�TJBFLG��igpERa��TC�݃������2TH2yN��� 1�b���Gq T�0 �$���M���`Ib���C�EF�1��� l�h��ENAB��lcTPE?@��� !(ᭀ����Q�#�@~�+2 H�W���2������"�4�F�X�j�3�қ{��������j�4�Ҝ��
��P.�@�R�j�5�ҝu�@����������j�6�����(:L�P
��7�ҟo���\�� ��8�����"4Fj�SMSK������a��E�A��MOT-E������@ "�1��Q�IO�5"%I(��P�QRd�Wi@��  �����X�gp�i�쐤��Y"$DS?B_SIGN4A�Q�i�̰C�ШP��S�232%�Sb�iDEVICEUS#|�R�RPARIT򱾈!OPBIT�Q���OWCONTR`��Q�ѓ�RCU� �M�SUXTASK��3NB��0�$TAT�U�P�1� @@쐦�F�6�_�PC}�$�FREEFROMqS]p�ai�GETN@�S�UPDl�ARB�� SP%0����� !m$US�A���az9�L�ER1I�0f��pRY�5~"�_�@f�P�1�!�6WRK��D9�F9�~�FRIEND�Q�4bUF��&�A@TO�OLHFMY5�$�LENGTH_VT��FIR�pqC�@��E� IUFINt�R���RGI�1��AITI:�xGX���I�FG2�7G1`a����3�B�GPRR�DA��O_� o0e�I1�RER�đ�3&���T�C���AQJV �G(|�.2���F��1�! d�9Z�8+5K�+5��E��y�L0�4�X T�0m�LN�T�3Hz���89��%�4�3G��W$�0�W�RdD�Z���Tܳ��K�a3d��=$cV 2���1���I1H�02K2
sk3K3Jci�aI��i�a�L��SL��R$)Vؠ�BV�EVk�]V*R��� �,6Lc����9V2F{/P:B��P5S_�E��$rr�C��ѳ$A0��wP!R���v�U�cSk�� p{�@#�2��� 0��D�VX`�!�tX`��P�0P�Ё�
�uSK!/� �-qR��!�0���z�NJ AX�!h�A�@LlA��A�/THIC�1�������1TFE���q>��IF_CH�3A�I00�����G1�x�������9�Ɇ_J�F҇PR(���R�VAT�� �`-p��7@����DO�E���COU(��AX�Ig��OFFSE+�TRIG�SK��c@���Ѽ�e�[�K�Hk�<��8�IGMAo0�A�-��ҙ�ORG_�UNEV��� ��S�쐮d ��$������GROU��ݓTO2��!ݓwDSP��JOG'�L�#	�_P'�2OR�p��>P6KEPl�#IR�0�PM�RQ�AP�Q��E�0q�e����SYSG��"��PG��BRK*Rd�r�3�-�������ߒ<p�AD��ݓJ�BSO�C� N�DUM�MY14�p\@SV��PDE_OP3S�FSPD_OVR�����CO��"�OIR-��N�0.�Fr�l.��OV�SFc�2�f��F��!4�S���RA�"LCHDL>�RECOV��0��W�@M�յ�R�O3��_�0�s @�ҹ@VERE��$OFS�@CV� 0BWDG�ѴC��X�2j�
�TR�!���E_FDOj�MOB_CM��U�B ��BL=r0�w�=q�tV@fQ��x0sp��_�Gx���AM��k�J0������_M��2{�#�8$CA�{Й���8$HBK|1c�ыIO��.�:!aPPA"�N�3�^�F����:"�DVC_DB �C��d�w"����!�Ց1���ç�3����ATIO� �q0�qUC�&CAB� BS�PⳍP�Ȗ���_0c�SUBCP	Uq��S�Pa aáĀ}0�Sb��c��r"ơ$HW_C��� :c��IcA�A-�l$U�NIT��l��AT�N�f����CYCL�ųNECA��[�F�LTR_2_FI`���(��}&��LP&������_SCT@SF�_��F����G���FqS|!�¹�CHAA�/����2��RSD��x"ѡb�r�: _T���PRO��O�� E%M�_��8u�q� u�q��DI��0e�RAILAC4��}RMƐLOԠdC��:anq��wq����+PR��SLQ�pf�C�ѷ 	��FUN9CŢ�rRINkP+a0�0 ��!RA� >R� 
Я�ԯW3AR�BLFQ���A�����DA`�����LDm0 �aB9��nqB�TIvrbؑ���PR�IAQ1�"AFS�P �!�����`%b����M�I1U�DFa_j@��y1°LME�{FA�@HRDY�4��Pn@RS@Q�0">�MULSEj@f�<b�q �X���ȑ���$.A$��1$c1Ó��߰� x~�EG0vpݓ�q!AR����09>B�%��A�XE��ROB��Wd�A4�_�-֣SY��h�!6��&S�'WR��r�-1���STR���5�9�E�� 	5B��=QB90�@6X������OT�0o ;	$�ARY8�w2h0���	%�FI��~;�$LINK��H��1�a_63�t5�q�2XYZ"� �;�q�3@��1�2�8%{0B�{D��� CFI��6G�0�
�{�_J��86��3aOP_O4Y;5�QTBmA"�B�C
�z�DU"�66CTURN3�vr�E`�1�9�ҍGFL�`@���~ �@�5<:7�^� 1�?0K�	Mc�68Cb�vrb�4�ORQ��X�>8 �#op������wq�Uf�8����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W���Tυ � ;����QH�!`�� ���U�Q�WkeK#kec�XER��	GE	0��S�dAWaǢ:D����7!�!AX �rB!{q��1u y-!y�pz�@z�@ z6Pz\Pz� z1 v�y�y�+y� ;y�Ky�[y�ky��{y��y�q�yDEBU��$����L�`!º2WG`  AB!��,��SV���� 
w���m���w����1 ���1���A���A��6Q ��\Q���!�m@��2.CLAB3B�U��x���S ? Ð�ER���� � i$�@� Aؑ!p�PO��Z�q0w�^��_MRAȑ� d�  T�ĴER1R��TYz�B��I�V3@�cΑTO	Q�d:`L� �d2��]�X�C[! �� p�`T}0i��_�V1�r�a'�4�2B-�2<����@P�����F�$W��g��5V_!�l�$�P����c��q"�	V F�ZN_CFG_!� 4��?º�|�ų��0��@�ȲW �P��\$� �n���Ѵ��09c�Q��(�FA�He�,�XEDM�(���H��!s�Q�g�P{R�V HELLĥ�� 56�B_BAS!�RSR��ԣo E�#S��[��1r�U%��2ݺ3ݺ4ݺU5ݺ6ݺ7ݺ8ݷ��ROOI䰝0�03NLK!�CAB� n��ACK��IN��T:�1�@�@ z�m�7_PU!�CO� ��OU��P� Ҧ) ���޶��TPFWD�_KARӑ��R�E~��P��(�Q�UE�����P
��C�STOPI_AL �����0&���㰑�0GSEMl�b�|�M��6d�TY|�SOK�}�DI�����(����_TM\�MANR�Q�ֿ0E+�|�$�KEYSWITCaH&	���HE
�OBEAT��cE� �LEҒ���U��F�O�����O_HOuM�O�REF�P�PRz��!&0��Cr+�OA�ECO��xB�rIOCM�D8׵����8�` G� D�1����U���&�MH�»P�CFO3RC��� ����OM�  � @�V��|�U,3P� 1(-�`� 3-�4���NPX_ASǢ�; 0ȰADD�����$SIZ��$�VARݷ TIPR]�\�2�A򻡐@���]�_� �"S��!Cΐ��FRIF�⢞�S�"�c���N�F��V ��` � x6�`SI�TES�R.6SSGL(T�2P�&��AU�� ) ST�MTQZPm 6ByW�P*SHOWb���SV�\$�w� ���A00P �a�6�@�J�TT�5�	6�	7�	8�	9�	A�	� �@!�'��0�F� 0u�	f0u�	�0u��	�@u[Pu%1�21?1L1Y1�f1s2�	2�	2��	2�	2�	2�	2��	222%2�22?2L2Y2�f2s3P)3�	3��	3�	3�	3�	3��	333%3�23?3L3Y3�f3s4P)4�	4��	4�	4�	4�	4��	444%4�24?4L4Y4�f4s5P)5�	5��	5�	5�	5�	5��	555%5�25?5L5Y5�f5s6P)6�	6��	6�	6�	6�	6��	666%6�26?6L6Y6�f6s7P)7�	7��	7�	7�	7�	7��	777%7�27?7,i7Y7�Fi7ss'� P��UPD�� � ��|�԰
,pY�SLOǢ� � z��и���o�E��`p>�^t��АALUץL����CU���wFOq�ID_L�ӿuHI��zI�$FILE1_���t��$`�^�vMsSA��� h��~�E_BLCK��#�C,�D_CPU <�{�<�o����t����R ��
�PW O� ��L�A��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ� �T�BCu�C� ��X -$�LEN@i��v������I���G�LOW_AXI��F1��t2X�M�����D�
 ��I�� 9��}�TOR��"��Dh��� L=�������s���#�_MA�`�ޕ��ޑTCV����T���&��@ݡ����J�����J����Mo���J�Ǜ ��)�����2�Ѓ �v�����F�JK��V�Ki�Ρv�Ρ3��J�0�ңJJڣJJ�AALң�ڣ���4�5z�&�N1�-�9���␅�L~�_�Vj�������{ ` �GROU�p�D��B�NFLI�C��REQUI;REa�EBUA��p����2¯����x�c�� \��/APPR��C����
�EN�CLOe��S_M v�,��
���� ���MC�&���g�_MG�q�C� �{ȸ9���|�BRKz�N�OL��|ĉ R��_CLI|��Ǫ�k�J����P
���ڣ�����&���/���6��6���8�������# ��8�%�W�2�e�PATHa�z�pӠz�=�vӥ�ϰ�x�CN=�CA�����p�IN�UC��bq��-CO�UM��YZ������qE%���2����~��PAYLOA���J2L3pR_AN��<�L��F�B�6�R��{�R_F2LSHR��|�LOG��р���ӎ���ACRL_@u�������.���H�p��$H{���FL�EX
��J�� :�/�����6�2�����;�M�_�F16����n���������ȟ��Eҟ���� �,�>�P�b���d� {������������5���T��X��v��� EťmFѯ��� ����&�/�A�S��e�+p�x�� � �������j�4pATر���n�EL  ԁ%øJ���ʰJEΧ�CTR�Ѭ�TN���F&��HAND_VB[
�pK�7� $F2{�6�, �rSWi�D�U��� $$Mt�h�R��08��@<b 35��^6A�p3�k��q{9�t�A�̈p��A��A��ˆ0��U���D��Dʴ�P��G��ISTЙ�$A��$AN��DY ˀ�{�g4�5D���v� 6�v��5缧�^�@��P�����#�,��5�>�D�J�� �&0�_�ER!V9�SQA'SYM��] ������x��ݑ���_SH l�������sT�(����(�:�JA���S�c�ir��_VI�#�Oh9�``V_UNI��td�~�J���b�E �b��d��d�f��n�@��������uN���9D��H�������"CqEN� a�D	I��>�Obt2Dpx��� ��2IxQA ����q��-��s �� ������ ��OMME��rr/�TVpPT�P ���qe�i����P�x ���yT�Pj� $�DUMMY9�o$PS_��RFq�s  ��:� �8��!~q� X�����K�STs�ʰSB}R��M21_Vt�8$SV_ERt�qO��z���CLRx�EA  O�r?p? Oր� � D $�GLOB���#LO ��Յ$�o��P�!wSYSADR�!�?p�pTCHM0 �� ,����W_NA��/�e����D�SR��l (:]8:m�K6� ^2m�i7m�w9m��9�� �ǳ��ǳ���ŕߝ�9 ŕ���i�L����m��_�_�_�T2��?TXSCRE�ƀ5�� ��STF���#}�pТ6�C�] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��tC�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$��VSHIF��|s�P�p�6��s���R���OSU�RW�pRADIz��2�_�q�h�g!� �q)�LUza�$OUTPUT_3BM��IML�oRp6(`)�@TIL<'SCO�@Ce�; ��9��F��T��a ��o�>�3�����Bw�2u�P{t���%�DJU��|#�/WAIT����ک�%ONE��Y�BOư ��� $@p%�C�SB�n)TPE��NEC���x"�$t$���*B_T��R��%�qR� $���sB�%�tM�+���t�.�F�R!݀��O�Pm�MAS�_DUOG�OaT	�D�����C3S�	�O2DELcAY���e2JO�� n8E��Ss4'#J�aP60%�����Y_��O2�$��2���5��`?{ sqZABCS�?�  $�2���J�
B��$$CL�AS������AB���'@@VIRqT��O.@ABS��$�1 <E�� < *AtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��.� @�R�d�v�����M@[�GAXLրK�*B�dC7  ���IN��ā���PRE������LARMRE?COV <I䂶��NG�� \K	? A   J�\��M@PPLIC�?�<E�E��Handling�Tool �� �
V7.50P/�28[�  ��c���
�_SW UP*A� F��F0ڑ����A��~�� 20���*A���:����o�FB 7wDA5�� �'@?�c@���None������� ��T'~*A4�bxl�E_��V����g�UTOB�ค����?HGAPON8@���LA��U��D 1<EfA����������� Q 1"שI Ԁ��Ԑ��:�i�n����#B{)B ����\�HE�Z�r�HTTHKY��$BI� [�m�����	�c�-� ?�Q�o�uχϙϫϽ� �������_�)�;�M� k�q߃ߕߧ߹����� ���[�%�7�I�g�m� ������������ W�!�3�E�c�i�{��� ������������S /A_ew��� ����O+= [as����� ��K//'/9/W/]/ o/�/�/�/�/�/�/�/ G??#?5?S?Y?k?}? �?�?�?�?�?�?COO O1OOOUOgOyO�O�O �O�O�O�O?_	__-_0K_Q_��(�TO4�s����DO_CLEA�N��e��SNM  9� �9oKo�]ooo�o�DSPDgRYR�_%�HI��m@&o�o�o#5 GYk}����0"���p�Ն �ǣ��qXՄ��ߢ��g�PLUGGҠ�Wߣ��WPRC�`B`9��o�=�OB��oe�/SEGF��K���� ��o%o����#�5�m���LAP�oݎ�� ��������џ������+�=�O�a���TO�TAL�.���USWENUʀ׫ �X����R(�RG_STRING 1���
�M��S�c�
��_ITE;M1 �  nc�� .�@�R�d�v������� ��п�����*�<��N�`�r�I/O SIGNAL���Tryout� Mode�I�np��Simul�ated�Ou�t��OVER�R�` = 100��In cyc�l���Prog� Abor���~��Status��	Heartbe�at��MH F�aulB�K�AlerUم�s߅ߗߩ߻����������  �S���Q��f�x�� ������������� ,�>�P�b�t�������,�WOR������V� ��
.@Rdv ��������*<N`PO ��6ц��o��� ��//'/9/K/]/ o/�/�/�/�/�/�/�/�/�DEV�*0� ?Q?c?u?�?�?�?�? �?�?�?OO)O;OMO�_OqO�O�O�OPALTB��A���O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o:o�OGRI�p��ra �OLo�o�o�o�o�o�o *<N`r�������`o��R B���o�>�P�b�t� ��������Ώ���� �(�:�L�^�p����PREG�N��.��� �����*�<�N�`� r���������̯ޯ����&����$AR�G_��D ?	����i���  	$���	[}�]}����Ǟ�\�SBN_C�ONFIG �i�������CI�I_SAVE  ���۱Ҳ\�TC�ELLSETUP� i�%HO�ME_IO�͈�%MOV_�2�8��REP���V�UT�OBACK
��ƽFRA:\�� �Ϩ���'` ��������� ����$�6��c�Z�lߙ��Ĉ�� �����������!凞 ��M�_�q����2� ��������%�7��� [�m��������@��������!3E$���Jo��������INI�@���ε��MESSA�G����q��OD�E_D$���Ox,0.��PAUS��!�i� ((Ol������� � /�//$/Z/H/�~/l/�/�'akTSK  q������UPDT%�d�0;WSM_CF°i�еU�'1�GRP 2h�93� |�B��A�/S�XoSCRD+11
1;' ����/�? �?�? OO$O��߳? lO~O�O�O�O�O1O�O UO_ _2_D_V_h_�O�	_X���GROUN�0O�SUP_NA�L�h�	�ĠV_�ED� 11;
 ��%-BCKEDT-�_`�!oEo$����a��o������ߨ���e2 no_˔o�o�b���eep�o"�o�oED3 �o�o ~[�5GED4�n#�� ~p�j���ED5Z� �Ǐ6� ~���}���ED6����k�ڏ ~pG���!�3�ED7�� Z��~� ~�V�şן�ED8F�&o��Ů�}����i�{�ED!9ꯢ�W�Ư
}3�����CRo���� �3�տ@ϯ����P�P?NO_DEL�_�R�GE_UNUSE��_�TLAL_OU�T q�c�QW?D_ABOR� ����Q��ITR_RT�N����NONS�e���CAM�_PARAM 1��U3
 8
�SONY XC-�56 23456�7890�H �� @���?�>��( АV�|[�r؀~�X�HR�5k�|U�Q�߿�R5y7����Aff���KOWA SC�310M|[r��>��d @6�|V ��_�Xϸ���V���  ���$�6��Z�l���CE_RIA_I�857�F�1���R|]��_LeIO4W=� ��P�<~�F<�GP 1.�,���_GxYk*C*  �V�C1� 9� @� iG� �CLC]� Ud� l� s�R� T��[�m� v� �� �� �� C�� �"�|W��7�{HEӰONFI� ���<G_PRI 1�+P�m®/���������'C�HKPAUS�  ;1E� ,�>/ P/:/t/^/�/�/�/�/ �/�/�/?(??L?6?h\?�?"O������H�1_MOR��� �0�5 	 �9 O�?$OOHO6K��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`ϖ�S:�(����Yp0�_)o�S`�BBia�P�_mo8j�(�aKoo�o9i�(�E�og�o�o�m�o�f�oGq:I�ZDE�F f8��)��R6pbuf.txAtm�]n�@�����# 	`(Ж�A=L����zMC�21B�=��9���4�=��n׾�Cz  B�HBCCo�C|���CqD���C���C��{iSZE@D���F.��F���E⚵F,�E�ٙ�E@F�N��IU��I?O��I<#I6��I�SY����vqG���Em��(�.��(�(���<�q�G�x2���2� �� a�D�j����E�e��EX�E�Q�EJP F��E�F� G��ǎ^F E��� FB� H�,- Ge��H�3Y���  >�33 ���NxV  n2xQ@��#5Y��8B� A�ASTo<#�
� �_�'�%��wRSMOF�S���~2�yT1>�0DE �O c�
�(�;�"�  Q<�6�z�R���?,�j�C4��SZm�E W��{�m�C��)B-G�C�`@$�q���T{�FPROG %i����c��I��� �Ɯ�f�KEY_TBL  �v�M�u� �	
��� !"#$�%&'()*+,�-./01c�:;�<=>?@ABC��pGHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����p����͓��������������������������������������������������?������!j��LCK��.�j���S�TAT���_AU_TO_DO���W�/�INDT_EN�B߿2R��9�+�Ty2w�XSTOP\��2TRLl�LET�E����_SCR�EEN i_kcsc��U���MMENU 1 ~i  <g\ ��L�SU+�U��p3g� ������������2� 	��A�z�Q�c����� ����������. d;M�q��� ���N%7 ]�m���/ ��/J/!/3/�/W/ i/�/�/�/�/�/�/�/ 4???j?A?S?y?�? �?�?�?�?�?O�?O -OfO=OOO�OsO�O�O �O�O�O_�O_P_Sy��_MANUAL���n�DBCOU�R�IG���DBNUIM�p��<���
�Q�PXWORK 1!R�ү�_oO.o�@oRk�Q_AWAYz�S��GCP ��9=��df_AL�P߄db�RY�������X_�p 1"�� , 
�^���o xvJf`MT�I^�rl@��:sONTIM��M����Zv�i
õ��cMOTNEND����dRECORD 1(R�a��ua�O��q��sb� .�@�R��xZ������ �ɏۏ폄���#��� G���k�}�����<�ş 4��X���1�C��� g�֟��������ӯ� T�	�x�-���Q�c�u� ���������>��� �)Ϙ�Mϼ�F�࿕� �Ϲ���:�������%� s`Pn&�]�o��ϓ�~� ����8�J�����5�  ��k����ߡ��J� ����X��|��C�U� ���������0������	��dbTOLEoRENCqdBȺb�`L�͐PCS_?CFG )�k)wdMC:\O �L%04d.CS�V
�Pc�)sA V�CH� z�P�)~���hMRC_�OUT *�[��`+P SGN �+�e�r��#�1�0-MAY-20� 10:33*V1�7-FEBj9:�09�k PQ��8��)~�`�pa�m��P�JPѬVERSION S�V2.0.8�.|EFLOGIC� 1,�[ 	�DX�P7)�PF."PROG_ENB�o\�rj ULSew �T��"_WRSTJ�NEp�V�r`dEMO�_OPT_SL �?	�es
 	R575)s7)�/�??*?<?'�$TO�  �-��?&V�_@pEX�Wd�u��3PATH ASA\�?�?O/{�ICT�aFo`-��gdse�gM%&ASTBF_TTS�x�Y^C��StqqF�PMAU� \t/XrMSWR.�i�6.|S/�Z! D_N�O0__T_C_x_�g_�_�tSBL_F�AUL"0�[3wTDIAU 16M6p��A1234567890gFP?BoTofoxo �o�o�o�o�o�o�o�,>Pb�S�pP�_ ���_s� � 0`�����)� ;�M�_�q����������ˏݏ��|)UMP��!� �^�TRp�B�#+�=�PMEfE~I�Y_TEMP9 È�3@�3A v��UNI�.(YN_?BRK 2Y)�EMGDI_ST�A�%WЕNC2_�SCR 3�� 1o"�4�F�X�fv����������#��ޑ14 ����)�;�����:ݤ5����� x�f	u�ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� �P�b�t�� ��xߞ� ����������
��.� @�R�d�v����� ��������*�<�N� ��r������������� ��&8J\n �������� "`�FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/4?,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O?�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �O�O�o�o�o
. @Rdv���� �����*�<�N� `�r����o����̏ޏ ����&�8�J�\�n� ��������ȟڟ�����H�ETMODE� 16���+ ��ƨ
R�d��v�נRROR_P�ROG %A�%��:߽�  ��TA�BLE  A�������#�L�RRS�EV_NUM  y��Q��K��S���_AUTO_?ENB  ��I��Ϥ_NOh� 7�A�{�R�  *U�������������^�+��Ŀֿ迄�H�ISO�͡I�}�_A�LM 18A� e�;�����+鿀e�wωϛϭϿ��_\H���  A����|��4�TCP_V_ER !A�!�����$EXTLOGo_REQ��{��V�SIZ_�Q�TOoL  ͡Dz���A Q�_BW�D����r���n�_D�I�� 9���}�z�͡m���STE�P����4��OP_�DO���ѠFA�CTORY_TU�N�dG�EATU�RE :�����l�Hand�lingTool� ��  - C�English� Diction�ary��ORDE�AA Vis��� Master����96 H��n�alog I/O����H551��u�to Softw�are Upda�te  ��J��m�atic Bac�kup��Part�&�groun�d Edit�� � 8\apC_amera��F���t\j6R�ell����LOADR�o�mm��shq��T7I" ��co���
! o���pa�ne�� 
!���tyle se�lect��H59��nD���onit�or��48����t�r��Reliab����adinDiagnos"�����2�2 ual �Check Sa�fety UIF� lg\a��ha�nced Rob� Serv q �ct\��lUse�r FrU��DI�F��Ext. D�IO ��fiA �d��endr E�rr L@��IF��r��  �П�9�0��FCTN M�enuZ v'��7}4� TP In���fac  SU_ (G=�p��_k Excn g��3��High-S�per Ski+� � sO�H9 � mm�unic!�onsg�teur� �����V����coknn��2��EN���Incrstr�u���5.fd�KAREL C�md. L?ua�A� O�Run-;Ti� Env����K� ��+%�s#�S�/W��74��Li�censeT� � (Au* ogB�ook(Sy��m�)��"
M�ACROs,V/�Offse��ap���MH� ����pf�a5�MechStop Prot��� d�b i�S�hif���j54�5�!xr ��#��,��qb ode �Switch��mK\e�!o4.�&� pro�4��g���Multi-�T7G��net.�Pos Re�gi��z�P��t� Fun���3 9Rz1��Numx ������9m�1�  A�djuj��1 J�7�7�* ����6t�atuq1EIKoRDMtot��_scove�� ���@By- }ues�t1�$Go� � U5\�SNPX b�"���YA�"LibAr����#�� �$�~@h�pd]0�Jt�s in VCC!M�����0�  �u!Ξ�2 R�0�/I��08��TMIL{IB�M J92�@�P�Acc>�F�9=7�TPTX�+�B�RSQelZ0�M8� Rm��q%��69�2��Unexce{ptr motnT  CVV�P���KC����+-��~K�  II)�VSP� CSXC�&.c��� e�"�� t�@�Wew�AD �Q�8bvr nmeYn�@�iP� a0�y�0�pfGrid~Aplay !� �nh�@*�3R�1M-1�0iA(B2015 �`2V"  F����scii�loa�d��83 M��l�����Guar�d 'J85�0�mP'�L`����stuaPat�&]$Cyc���|0�ori_ x%Dat�a'Pqu���ch��1��g`� j� RLJam�5���I_MI De-B(\A^�cP" #^0C�  etkc^0a�sswo%q�)65�0�ApU�Xnt\��Pven�CTq�H�5�0YEL?LOW BO?Y���� Arc�0vis���Ch�Weld�Qcial4Izt��Op� ��gs�` �2@�a��poG yRjT1 NE�#3HT� xyWb��#! �p�`gd`����p\� =P��JPN� ARCP*PRx�A�� OL�pwSup̂fil�pp��J�� ��cro�6�70�1C~E�d��SuS�pe�tex�$Y �P� So7 t� /ssagN5 <Q�B�P:� �9 "0�Qr�tQC��P�l0dpn�笔�rpf�q�e��ppmasc�bin4psyn��' ptx]08�H�ELNCL V�IS PKGS �Z@MB &��B� J8@IPE �GET_VAR �FI?S (Uni�� LU�OOL: �ADD�@29.F�D�TCm���E�@D�Vp���`A�ТNO� WTWTEST� �� ��!��c�F�OR ��ECT ��a!� ALSE �ALA`�CPMO�-130��� b D�: HANG F�ROMg��2��R�709 DRAM� AVAILCH�ECKS 549���m�VPCS S�U֐LIMCHK���P�0x�FF P�OS� F�� q�8-12 CH�ARS�ER6�OG�RA ��Z@AVE�H�AME��.SV���Вאn$��9�m� "y�TRCv� �SHADP�UPD�AT k�0��ST�ATI��� MU�CH ���TIM�Q MOTN-0�03��@OBO�GUIDE DAUGH���b��@$Gtou� �@C� �0���PATH�_�M�OVET�� R6�4��VMXPAC�K MAY AS�SERTjS��CY�CL`�TA��BE COR 71�1�-�AN��RC O�PTIONS  ��`��APSH-1N�`fix��2�SO���B��XO򝡞�_TP��	�i��0j��du�{byz p wa���y�٠HI������U��pb XSPD T�B/�F� \hch�ΤB0���END�C�E�06\Q�p{ s>may n@�p�k��L ��traff#�	� ��~1�from sysvar scr�0qR� ��d�DJU����H�!A��/��S?ET ERR�D��P7����NDAN�T SCREEN� UNREA V�M �PD�D��PA����R�IO J�NN�0�FI��B���GROUNנD� Y�Т٠�h�S�VIP 53 QS���DIGIT V�ERS��ká�NE�W�� P06�@C�1IMAG�ͱ���8� DI`���p�SSUE�5��EP�LAN JON� gDEL���157QzאD��CALLI�ॡQ��m���IPN�D}�IMG N9� PZ�19��MN;T/��ES ���`wLocR Hol߀�=��2�Pn� PG:t��=�M��can������С: 3D �mE2view d3 X��ea1 �0�b�pof Ǡ"H�Cɰ�ANNOT� ACCESS �M cpie$Etn.Qs a� loMd�Flex)a:��w^$qmo G�sA9�a-'p~0��h0pa���eJ AUTO-�0��!ipu@Т<ᾡ�IABLE+� �7�a FPLN: �L�pl m� M�D<�VI�и�WI�T HOC�Jo�~1Qui��"��N���USB�@�Pt & remov����D�vAxis F�T_7�PGɰCP�:�OS-144� � h s 26�8QՐOST�p  �CRASH DU���$P��WORD�.$�LOGIN̈P��P:	�0�046 issueE��H�: Slow� st�c�`6Й���໰IF�IM�PR��SPOT:�Wh4���N1STY<��0VMGR�b�N�CAT��4oRR�E�� � 58t�1��:%�RTU!Pre -M a�SE:�@!pp���AGpL��9m@all��*0va�OCB WA����"3 CNT0 �T9DWroO0al�arm�ˀm0d �t�M�"0�2|� o�Z@OME<�� ���E%  #1-�SR�E��M�st}0g �    5KA�NJI5no M�NS@�INIS�ITALIZ'� E�f�we��6@� �dr�@ fp "~��SCII L�afails w�>�SYSTE[��i��  � Mq�1�QGro8�m n@�@vA����&��n᰼0q��RWRI O�F Lk��� \r�ef"�
�up� d�e-rela�Qd� 03.�0SSc}hőbetwe4�IND ex ɰTPa�DO� l�y �ɰGigE�s�operabil.`p l,��HcB�̚@]�le�Q0cf�lxz�Ð���OS� {����v4pfigi GLA�$�c2��7H� lap�0A[SB� If��g�2 l\c�0�/��E�� EXCE �㰁�P���i�� Do0��Gd`]Ц�fq��l lxt��EFal��#0�i�O�Y��n�CLOS��SR�Nq1NT^�F�U�FqKP�ANIO V7/ॠ1�{����DB �0��ᴥ�;ED��DET|�'�� �bF�NLINEb�BUG�T���C"RLIB��A���ABC JARK�Y@��� rkey��`IL���PR��N\��ITGAR� D$��R �Er *�T���a�U�0��h�[�Z�E V� TAS�K p.vr�P�2" .�XfJ�srn8�S谥dIBP	c�v��B/��BUS��UNN� j0-�{�d�cR'���LOE�wDIVS�CULs0$cb����BW!���R~�W`P�����ITd(঱tʠ�OF���UNEXڠ+���p��FtE��SVEM�G3`NML 50�5� D*�CC_SAFE�P*� �ꐺ� PET��'P�`�gF  !���IR����c i S>� K���K�H GUN�CHG��S�MEKCH��M��T*��%p6u��tPORY_ LEAK�J����SPEgD��2Vw 74\GRI�x�Q�g��CTLN��TRe @�_�p ���EN'�IN�����0�$���r��T3)�iԗSTO�A�s�L���͐X	���q��Y� ��TO2�J m���0F<�K����DU��S��O��3 �9�J F�&���SSVGN-1#I���'RSRwQDAU�Cޱ � �T6�g��� 3�]�~��BRKCTR/"� �q\j5��_�QܺS�qINVJ0D ZO�Pݲ���s��г��Ui ɰ̒�a�DU{AL� J50e��x�RVO117 AW�TH!Hr%�N�7247%�52��|�&aol ���R���at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���Md��Rǰt� \fosB�A�0Np�c�����{�U��ROP 2��b�pB��ITP4aM��b !AUt �c0< � plete��N@� z1^qR�635 (Acc_uCal2kA���I) "�ǰ�1a\�Ps��ǐ� bЧ0�P򶲊���ig\�cbacul "A3p_ �1��ն���_etaca��AT����PC�`�����_p�.pc!Ɗ��:�circB���5��tl��Bɵ�:�fm+�Ί�V�b�ɦ�r�?upfrm.����ⴊ�xed��Ί�~�'pedA�D �}b�ptlibB�� ߆_�rt��	Ċ�_0\׊ۊ�6�fm�݊��oޢ�e��̆Ϙ���c��Ӳ�5�j>�����tcȐ��	�r����emm 1��T�sl^0���T�mѡ�#�rm�3��ub Y�q�st�d}��pl;�&�c1kv�=�r�vf�䊰���9�vi����u�l�`�0fp�q �.yf��� daq; �i Data Ac_quisi��n��
��T`��1�8�9��22 DMCM RRS2Z��75��9 3 Rg710�o59pq5\?��T "���1 (D�T� n k@��������E Ƒȵx��Ӹ�etdmm F��ER����gE<��1�q\mo?۳ �=(G���[(

�2�` ! �@J�MACRO��Sk�ip/OffseP:�a��V�4o9� &qR662���Rs�H�
 6Bq8�����9Z�43 J�77� 6�J783�o ��n�"v��R5IKCBq2� PTLC�Zg� R�3 (�s,� �������03��	зJԷ\sfm�nmc "MNM�C����ҹ�%mnf�FMC"Ѻ0ª etmcr� �8����� ,��qD�q �  874\prdq>,jF0����axisHPro�cess Axe�s e�rol^P�RA
�Dp� 56 �J81j�59� 5�6o6� ���0w�6�90 98� [!IDV�1��2(x2��2ont�0�
�����m2���?C��etis "ISD��x9�� FpraxRA�M�P� D��de�fB�,�G�isb/asicHB�@޲�{6�� 708�6
��(�Acw:�����@�D
�/,��AMOX��  ��DvE��?;T��>Pi� RAFM';�]�!PAM�V�W�Ee�U0�Q'
bU�75�.��ceNe� nterface^�1' �5&!54�K��b(Devam±�/�#��Э/<�Tane`"D�NEWE���btpd/nui �AI�_s~2�d_rsono����bAsfjN��bdv_arFvf�xhp�z�}w��hkH9xs�tc��gAponlGzv{�ff��r ���z�3{q'Td~>pchampr;re�p� ^5977� �	܀�4}0��mɁ�/������lf�!�pcc7hmp]aMP&B<�� �mpev������pcs��YeS~�� Macro�O	D��16Q!)*�:$��2U"_,��Y�(PC ��$_;������o|��J�gegemQ@�GEMSW�~ZG�g�esndy��OD�n�dda��S��syT�Kɓ�su^Ҋ����n�m���L��  �	��9:p'ѳ޲���spotplus�p���`-�W�l�J�s⽱t[�׷p�key �ɰ�$��s�-Ѩ�m�~��\featu 0�FEAWD�oolo�srn'!2 �p���a�As3��tT�.� (N. A.)��!e!�J# (j�,��oBIB�o�D -�.�n��k9�"K��u[-�_���}p� "PSEq�W����wop "sEЅ�&�:�J����� �y�|��O8��5��R ɺ���ɰ[��X�� �����%�(
ҭ�q HL�0k�
�z�a !�B�Q�"(g�Q �����]�'�.����ɀ&���<�!ҝ_�#��tpJ�H�~Z��j����� y������2��e��� ���Z����V��!%���=�]�͂��^2�@i[RV� on�QYq͋JF0� 8ހ�`�	�(^�dQueue���X\1�ʖ`�+F1�tpvtsn��N�&��ftpJ0v �R�DV�	f��J1 Q4���v�en��k/vstk��mp��~btkclrq���get�����r��`kack8�XZ�strŬ�%��stl��~Z�np:!�`���q/��ڡ6!l�/Yr�mc�N+v3�_� ���l�.v�/\jF��� �`Q�΋ܒ��N50 (FRA���+��͢frap�arm��Ҁ�} 6��J643p:V�E�LSE
#�VA�R $SGSYS�CFG.$�`_U?NITS 2�DG0~°@�4Jgfr��4A�@FRL-��0ͅ�3 ې���L�0NE�:� =�?@�8�v�9~Qx3�04��;�BPRS�M~QA�5TX.$VNUM_OL��85��DJ507��l�? Functʂ"q�wAP��琉�3 HH�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6 N�kAP����S��"TPPR���Q.A�prnaSV�ZSx��AS8Dj510U�-�`cr�`8 ��ʇ��DJR`jYȑH � �Q �PJ�6�a21��48AAVM 5�Q�b0 lB�`TUP� xbJ5459 `b�`616���0VCAM 9��CLIO b1��5 ���`M�SC8�
rP R`\�sSTYL �MNIN�`J62�8Q  �`NRExd�;@�`SCH ���9pDCSU Me�te�`ORSR �Ԃ�a04 kR_EIOC �a5�`542�b9vpP<� nP�a�`�R�`7�`��MASK H�o�.r7 �2�`O'CO :��r3��p�b�p���r0X��a�`�13\mn�a39 HRM"�q�q�ҿLCHK�uO�PLG B��a03� �q.�pHCR �Ob�pCpPosi��`fP6 is[rJ�554�òpDSWĤbM�D�pqR�a37� }Rjr0 �1�s4i �R6�7��52�rs5 �2�r7 1� �P6���Regi��@T�uFRDM��uSaq%�4�`93�0�uSNBA�uSwHLB̀\sf"p�M�NPI�SP{VC�J520���TC�`"MNрT�MIL�IFV�P�AC W�pTPT�Xp6.%�TEL�N N Me�0�9m3UECK��b�`UFR�`��V�COR��VIPL:pq89qSXC�S�`�VVF�J�TP ��q��R626l�u� S�`Gސ�2�IGUI�C��PG�St�\ŀH863`�S�q�����q34sŁ684���a��@b>�3 :B��1 \T��96 .�+E�g51 y�q53�3f�b1 ���b1 n��jr9 ���`VAT9 ߲�q75 s�F�<�`�sAWSM��`�TOP u�ŀR582p���a80 
�ށgXY q���0 ,b��`885�QXрO�Lp}�"pE࠱tp��`LCMD��ET3SS���6 �V��CPE oZ1�V�RCd3
�NLH�h���001m2Ep��3� f��p��4 /1�65C��6l���7zPR��008 tB~��9 -200�`�U0�pF�1޲1 ��޲2L"���p��޲y4��5 \hmp~޲6 RBCF�`0ళ�fs�8 �Ҋ���~�J�7 rbc	fA�L�8\PC�����"�32m0u�n�K�R�ٰn�5 5EW�
n�9 z��40Y kB��3 ��6ݲ��`00iB/��6$�u��7�u��8 µ������sU0�`�t �1 05\rb��2 E���K���j�2��5˰��60��a�HУ`:�63�jAF�_����F�7 ڱ݀H�80�eHЋ��cU0��I7�p��1u��8u��9 73�������D7� ��5t�9+7 ��8U�1��2J��1�1:���h���1np�"��8(�U1��\pyl��,࿱�v ��B�854��1hV���D�4��im�с1�<���>br�3�pr�4@pGPr�6 !B���цp��1�����1�`͵155ض1g57 �2��62�S����1b��2����1Π"�2���B�6`�1<c�4 L7B�5 DR��8_�{B/��187 u�J�8 06�90� rBn�1 (��202 0EW,ѱ�2^��2��90�U2��p�2��2 b��4:��2�a"RB����9\�U2�`w�l���O4 60Mp��7��`����b�s
5 ���3����pB"9 3a ����`ڰR,:�7 �2��V�2��5@���2^��a^9��B�qr����n�5����5᥁"�8a�Ɂ}Չ5B���5����`U�A���� ��86 �6 S�0��5�p�2�#�529 �2^�Tb1P�5~�2`P���&P5��8��5��u�!�5��ٵ5+44��5��R�ąPa nB^z�c (�a4�����U5J�
V�5��1�1^��%������5 b21���gA��58W8-2� rb��5N�E�G5890r� 1�95 �"������c 8"a��|�L ���!J"E5|6��^!�6���B�"8�`#��+�8�%�6B�AME�"1w iC��622�B�u�6V��d� 4��8�4�`ANRSP�e?/S� C�5� �6� ��� \� �6� ��V� 3t��� TG20CA�R��8� pHf� 1DH�� AOE�� �� ,�|�� �0\�� �!64K��ԓrA� �1� (M-7�!/50T�[PM��P�Th:1�C�#Pe� �3��0� 5`M75T1"� �D8p� �0Gc�� u�4��i1-710i�1� Skd�7j�z�?6�:-HS,�  �RN�@�UB�f�X�=m75sA*A6a�n���!/CB�B2.6A �0;A�CIB�A�2P�QF1�UB2�21� �/70�S� �4��� �Aj1�3p���r�#0 B2\m*A@C@��;bi"i1K�u"A~A�AU� imm7c7@��ZA@I�@�Df�Ab�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A��EA�5B�4>\77
B7=Q�D�2�Q$B�E)7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E"l7�@7�A
1�E�V~`��W2%Q�R9ї@0L_�#����"A����b��H3s=rA/2 �R5nR4�74rNUQ1�ZU�A�s\m9
1M�92L2�!F!^Y�ps�� 2ci��-?�qhimQ�t  w043�C�p�2�mQ�r�H_ �H20��Evr�QHsXBSt62�q`s����� ��P�xq350_*A3I)�2�d�u0�@� '4kTX�0�pa3i1�A3sQ25�c��s�t�r�VR1%e�q0 
��j1��O2 �A �UEiy�.�‐ �0C2h20$CXB79#A�����M Q1]�~�� 9 �Q��?PQ��qA!Pvs � 5	15aU���?P�Ņ���ဝQ9A6�zS*�7�qb5�1��8��Q��00P(��V7]u�aitE1���ïp�?7� !?�z��rbUQRB1PM=�Qa9p��H��QQ�25L��@�����Q��@L���8ܰ��y00\r�y�"R2BL�tN�  ��� �1D�q�2�qeR�5���_b�3�X]1/m1lcqP1�a�ED�Q� 5F����!5���@M-16Q�� f� ��r��Q�e� ��� PN�LT_�1��i1��9453��@�e�|�b1l>F1u*AY2�
��R8�Q���RJ�J3�D}T� 85
Qg�/0��*A!P� *A�Ð𫿽�2ǿپ6t�6=Q���P�X���� AQ� g� *ASt]1^u�ajrI�B ����~�|I�b��yI�\m�Qb�I�uz�A��c3Apa9q� B6S���S��m���}�85�`N�N�   �(M���f1���6��P��161��5�s`҃SC��U��A����5\set06c��f��10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C����5�B��B��h`�F��� X0���A:���C�M��!AZ��@��4�6i����� e�O�-	���f 1��F �ᱦ�1F�8Y	���T6HL3��BU66~`���U�dU�9D20Lf0��Qv�  ��fjq��N������ 0v
� ��i	�	��72lqQ2�������� \chngmOove.V��d��|��@2l_arf 	�f~��6���� ��9C�Z���~���kr41 S���0��V���t�����U�p7nuqQ%�A]��V�1\�Qn�BJ�2W�EM!5���)�#:�64��F�e50S�\��0�=� PV���e�������E�����m7shqQSH"U��)��9�!A��(���� ,�q�����TR1!��,�6�0e=�4F�����2��	 R-������ �����Ж��4���LSR�)"�!lO�A��Q�) %!� 16�
U/��2�"2�E��9p���2X� SA/Ai��'�
7F�H�@ !B�0��D���5V� �@2cVE��p��T��pt갖�1L~E�#�Fd�Q��9E�#De/��RT��59���	�A�E�iR������9\m20�20��+�-u�19r4�`�E1�=` O9`�1"ae��O��2��_$W}am41��4�3�/d1c_std��1)�!�`�_T��r�_ 4\jdg�a�q�PJ%!~` -�r�+bgB��#c'300�Y�5j�QpQb1�bq��vB��v�25�U�����qm43� �Q<W�"Ps� �A��e����t� i�P�W.��c�F�X.�e�kE14�4y4�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf��`coWo!\�2a��K2A;_2��QW2�`bF�(�V11�23�`���X5�Ra21�J�*9�a:88J9X�l5�m1a첚��*���(85�&��������P6���R,52&A����,fA9IfI'50\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP 1��vB)e�m�����ު1p� �1D��q�27�F�KAR�EL Use S���FCTN��� �J97�FA+�� �(�Q޵�p%�)?�Vj�9F?(�j�Rtk208 "Km�6Q�yB�j��iæPr�9�sx#��v�krcfp��RCFt3���Q��k�cctme�!ME�g����6�mainj�dV�� ��ru��kDº�c���o����&J�dt�F �»��.vrT�f�����E�%�!��5�FRj73�B�K���UER�HJn�O  J�� (ڳF���F�q�Y�&T��`p�F�z��19�tkvBr���V�h�9p�E�y�<�k������;�v���"CT��f���� )�
І��)�V	�6� ���!��qFF��1q� ��=�����O�?�$"����$��je���TC�P Aut�r�<5�20 H5�J5�3E193��9��96�!8��9��	 �B�574��52�J:e�(�� Se%!Y������u��ma�Pqtool�ԕ�����~�conrel�F�trol Rel�iable�RmvCU!��H51�����8 a551e"�CNRE¹I��c�&��it�l\s�futst "UaTա��"X�\u�� g@�i�6Q]V0�B,Eѝ6A� �Q�)C ���X��Yf�I�1|�6s@6i��T6I U��vR�d�
$e%1���2�C58�E6��8`�Pv�iV4OFH58SOteJ� mvBM6E~O58�I�0�E�#+@� &�F�0���F�P6a����)/++�</N)0\�tr1�����P ,��qɶ�rmask�i�msk�aA���k�y'd�h	A	�P�sD�isplayIm��`v����J887# ("A��+Heůצprds��Iϩǅ�Uh�0pl�2�R2���:�Gt�@��PRD �TɈ�r�C�@Fm��D��Q�AscaҦ� �V<Q&��bVvbrl �eې@��^S��&5U�f�j8710�yl 	��Uq���7�&�p��p��P^@�P�firmQ����Pp�2�=b�k�6�r�3��6��t7ppl��PL���O�p<b�ac�q	��g1�J�U�d�J��gait_9e��Y�&��Q����	�Shap��e?ration�0��R67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G����qF�205p�5pS���Ձ�retsap��BP�O�\s� O"GCR�ö? �q/ngda�G���V��st2axU��Aa]��bad�_�btputl/�&�e�>��tplibB_���=�2.����5���c3ird�v�slp���x�hex��v�re8?�Ɵx�key�v�cpm��x�us$�6�gcr��F�����8�[�q27j92�v��ollismqSk��9O�ݝ� (pl�.���t��p!o��2 9$Fo8��cg7no@ƿtptcls` C�LS�o�b�\�km�ai_
�s>�v�o	��t�b���ӿ�E�H��6�1enu5�01�[m��uti|a|$calmaUR���CalMateNT;R51%�i=1]@ -��/V� ��Z�� �tfq1�9 "K9E��L����2m�CLcMTq�S#��et ��LM3!} �F�c��nspQ�c���c�_moq��� ��c1_e�����su��ޏ� �_ �@�5�G�join�i�j��oX��ł&cWv	 ���N�v9e��C�clm�&A�o# �|$finde��0STD �ter FiOLANG���R���
��n3��z0Cen���r,������ J����� ���K�〪Ú�=���_Ӛ��r~� "FNDR��� 3��f��tguid�䙃N�."��J�tq�� ��������� ����J����_������c��	m�Z��?\fndr.��n#�>
B2p��Z�CP� Ma�����38PA��� c��6� (�� �N�B�������H 2�$�81��m_���"ex�z5� .Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$�r*$ ��*$r*$%/s#C�d/�.,P�/0*ʲD�PN��$���$*�G}r�$k Exc�'{IF�$MASK�%�93 H5�%H5�58�$548 H��$4-1�$��#1(�$�0 E�$��$-b��$���!UPDT ��B�4�b�4�2�49�0`�4a�3�9j0"M�4<9�4  ��4��4tpsh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4���3adq\�5K�979":E�ajO l "DQ^E^�3�i�Dq ��4ҲO ?R�? ��q�5��T���3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F��t�4��.�5y N� >�2il(in�4��31 JH1�2Q4�2�51ݠ�4rmal� �3)�REo�Z_�� �Ox����4��^F�?onorTf��7_ja�UpZҒ4l�5rmsAU��Kkg���4�$HCd\��fͲ�eڱ�4�REM����4yݱ"u@�RERG5932fO��47Z�>�5lity,�U��8e"Dil\�5�r�o ��7987�?8�25 �3hk910�3 ��FE�0=0P_�Hl\mhm�5� �qe�=$�^�
E��u<�IAymptm�U��BU��vste�y\� 3��me�b�DvI�[�Qu �:F�Ub�*_�
E&,�su��_ E�r��ox���4hu#se�E-�?�sn��������FE��,�box�����c݌,"��� ����z��M��g��pdspw)�	�� 9���b���(��1���c��Y�R��  �>�P���W��������'�0ɵ�[���͂���  �w ,�@� �zA�bumpšuf��B*�Box%��7Aǰ60�BBw���MC� (6�,f�t{ I�s� ST���*��}B�����w��"BBF
�>�`����)��\bbk968 "�4��։�bb�9va69�����etbŠ��X�����ed	�F��1u�f� �sea"������'�\��,���b�ѽ�o6�H�
�	x�$�f���!y����Q[�! tpermr�fd� TPl0~o� Recov,���3D��R642� � 0��C@}s� tN@��(U�rro����yu2r��  ?�
  �����$$CLe� O�������������$z�_DIGsIT��������.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$j����+c:PRODU�CTM�0\PGSTKD��V&ohozf�99��D����$FEAT_I�NDEX��xd���  
��`ILECOMPW ;���#��`��cSETUP2� <�e�b��  N �a�c_�AP2BCK 1�=�i  �)�wh0?{%&c�� ��Q�xe%�I� m���8��\�n� ���!���ȏW��{� �"���F�Տj���w� ��/�ğS������� ��B�T��x������ =�үa������,��� P�߯t������9�ο �o�ϓ�(�:�ɿ^� ��Ϗϸ�G���k�  �ߡ�6���Z�l��� ��ߴ���U���y�� ���D���h��ߌ�� -���Q��������� @�R���v����)��� ��_�����*��N ��r��7�� m�&�3\�i�
pP 2#p�*.VRc�*��� /���PC/1/FR6:/].��/+T�`�/�/F%�/�,�`xr/?�*.F�D8?	H#&?e<�/<�?;STM �2�?н.K �?�=i�Pendant �Panel�?;H �?@O�7.O�?y?�O:GIF�O�O�5�OoO8�O_:JPG _J_��56_�O_�_�	P�ANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEINS.XML���0\���qC�ustom To�olbar	���PASSWORD�yFRS:\�L�� %Pas�sword Config���֏e� Ϗ�B0���T�f��� �������O��s�� ����>�͟b��[��� '���K��򯁯��� :�L�ۯp�����#�5� ʿY��}��$ϳ�H� ׿l�~�Ϣ�1����� g��ϋ� ߯���V��� z�	�s߰�?���c��� 
��.��R�d��߈� ��;�M���q���� ��<���`������%� ��I��������8 ����n���!�� W�{"�F� j|�/�Se ��/�/T/�x/ /�/�/=/�/a/�/? �/,?�/P?�/�/�?? �?9?�?�?o?O�?(O :O�?^O�?�O�O#O�O GO�OkO}O_�O6_�O /_l_�O�__�_�_U_ �_y_o o�_Do�_ho �_	o�o-o�oQo�o�o �o�o@R�ov ��;�_��� *��N��G������ 7�̏ޏm����&�8� Ǐ\�돀��!���E� ڟi�ӟ���4�ßX� j��������įS���w������B�#��$�FILE_DGB�CK 1=���/���� ( �)
SU�MMARY.DG<L���MD:������Diag Summary���Ϊ
CONSLO�G�������D�ӱ�Console �logE�ͫ��MEMCHECK:��!ϯ���X�Mem�ory Data|��ѧ�{)��HADOW�ϣϵ��J���Shado�w Change�sM�'�-��)	FTP7Ϥ�3ߨ����Z�mment� TBD��ѧ0=�4)ETHERNET�������T��ӱEthern�et \�figu?rationU�ؠ~��DCSVRF��p�߽�����%��� verify �all��'�1PY=���DIFF�����[���%��d�iff]������1pR�9�K��� ����X��CHGAD������c��r����2ZAS�� ��GD ���k��z��FY3bI[�� �/"GD ���s/����/�*&UPDATE�S.� �/��FR�S:\�/�-ԱU�pdates L�ist�/��PSRBWLD.CM(?����"<?�/Y�PS�_ROBOWEL ��̯�?�?��?&�O -O�?QO�?uOOnO�O :O�O^O�O_�O)_�O M___�O�__�_�_H_ �_l_o�_�_7o�_[o �_lo�o o�oDo�o�o zo�o3E�oi�o ���R�v� ��A��e�w���� *���я`�������� �O�ޏs������8� ͟\�����'���K� ]�쟁����4���ۯ j������5�įY�� }������B�׿�x� Ϝ�1���*�g����� Ϝ���P���t�	�� ��?���c�u�ߙ�(� ��L߶��߂���(� M���q� ���6��� Z������%���I��� B�����2�����h�����$FILE�_� PR� ���������MDONLY� 1=.�� 
 ���q����� �����~%� I�m�2� �h��!/�./W/ �{/
/�/�/@/�/d/ �/?�//?�/S?e?�/ �??�?<?�?�?r?O �?+O=O�?aO�?�O�O &O�OJO�O�O�O_�O�9_�OF_o_
VIS�BCKL6[*�.VDv_�_.PF�R:\�_�^.P�Vision V?D file�_�O 4oFo\_joT_�oo�o �oSo�owo�oB �of�o�+�� �����+�P�� t������9�Ώ]�� ����(���L�^���� ���5���ܟk� ��� $�6�şZ��~������
MR_GRPw 1>.L���C4  B���	� W������*u���R�HB ��2 ���� ��� ���B�����Z�l��� C���D�������Ŀ���K�
�J�}��I���T���EF�5UP���{���ֿ E��M.G�E$���;n߇:G���@O���@��@��Ef���2�@���@��p
*λ� F�@ �������J���NJk�H�9�Hu��F!��IP�s��?����(�9�<�9�89�6C'6<,6\b��+�&�(��a�L߅�p�A��A� �߲�v���r������ 
�C�.�@�y�d��� �����������?��Z�lϖ�BH�� A�Ζ�������
0��PS@�P�TR0��ܿ� �B���/ ���@�33:���.�gN�UUU�U���q	>u.�?!rX��	��-=[z�=��̽=V6<��=�=�=$�q�����@8��i7G��8��D�8@9!�7�:�����D�@ D�� �Cϥ��C������'/0-��P/��� �/N��/r��/���/� ??;?&?_?J?\?�? �?�?�?�?�?O�?O 7O"O[OFOOjO�O�O �O�O�гߵ��O$_�O H_3_l_W_�_{_�_�_ �_�_�_o�_2ooVo hoSo�owo�o�i��o �o�o��);�o_ J�j����� ��%��5�[�F�� j�����Ǐ���֏� !��E�0�i�{�B/�� f/�/�/�/���/��/ A�\�e�P���t����� ���ί��+��O� :�s�^�p�����Ϳ�� �ܿ� ��OH��o� 
ϓ�~ϷϢ������� ���5� �Y�D�}�h� �߳ߞ��������o� 1�C�U�y��߉�� �����������-�� Q�<�u�`��������� ������;&_ J\�������� ��ڟ�F�j4� �������� !//1/W/B/{/f/�/ �/�/�/�/�/�/?? A?,?e?,φ?P�q?�? �?�?�?O�?+OOOO :OLO�OpO�O�O�O�O �O�O_'__K_�o_ �_�_�_l��_0_�_�_ �_#o
oGo.okoVoho �o�o�o�o�o�o�o C.gR�v� ����	���<� `�*<��`��� ��ޏ��)��M�8� q�\�������˟��� ڟ���7�"�[�F�X� ��|���|?֯�?���� �3��W�B�{�f��� ��ÿ��������� A�,�e�P�uϛ�b_�� ���Ϫ_��߀�=�(� a�s�Zߗ�~߻ߦ��� ����� �9�$�]�H� ��l���������� ��#��G�Y� �B��� ����z�������
ԏ :�C.gRd�� ����	�? *cN�r��� ��/̯&/�M/� q/\/�/�/�/�/�/�/ �/?�/7?"?4?m?X? �?|?�?�?�?�?��O !O3O��WOiO�?�OxO �O�O�O�O�O_�O/_ _S_>_P_�_t_�_�_ �_�_�_�_o+ooOo :oso^o�o�op��o��  ��$��o �o�~����� ��5� �Y�D�}�h� ������׏���� 
�C�.�/v�<���8� �����П����?� *�c�N���r������� �̯��)��?9�_� q���JO�����ݿȿ ��%�7��[�F�� jϣώ��ϲ������� !��E�0�i�T�yߟ� ���߮��߮o�o��o >�t�>��b�� ���������+��O� :�L���p��������� ����'K6o Z�Z�|�~���� �5 YDi� z������/ 
//U/@/y/@��/�/ �/�/���/^/??? Q?8?u?\?�?�?�?�? �?�?�?OO;O&O8O qO\O�O�O�O�O�O�O��O_�O7_��$F�NO ����VQ��
F0fQ kP F�LAG8�(LRR�M_CHKTYP�  WP��^Pk�WP�{QOM�P�_MIN�P���}�P�  XNP�SSB_CFG �?VU ��_���S oo�IUTP_DEF__OW  ��R>&hIRCOM�P8o��$GENOVRoD_DO�V�6�nflTHR�V d�e�dkd_ENBWo �k`RAVC_G�RP 1@�WCa X"_�o_1 U<y�r��� ��	��-��=�c� J���n��������ȏ ����;�"�_�F�X�\��ibROU�`FVX.�P�&�<b>&�8�?������������  �D?�јs���@@g�B�7�p�)�ԙ����`SMT�cG�m�M���� �LQHOS�TC�R1H���Ps��at�SM���f�\���	_127.0��1��  e��ٿ��� ��ǿ@�R�d�vϙ��0�*�	anonymous�������ό���[�� � �����r����ߨ� ������-���&�8� [�I�π������ ���1�C��W�y��� `�r������ߺ����� ��%�c�u�J\n ��������� M�"4FX��i� �����7// 0/B/T/���m/� �/�/�/??,?�/ P?b?t?�?�/�?��? �?�?OOe/w/�/�/ �?�O�/�O�O�O�O�O =?_$_6_H_kOY_�? �_�_�_�_�_'O9OKO ]O__Do�Ohozo�o�o �o�O�o�o�o
?o }_Rdv���_�_ oo!�Uo*�<�N� `�r��o������̏ޏ �?Q&�8�J�\���~>�ENT 1I��� P!􏪟  ����՟ğ���� ���A��M�(�v��� ^�����㯦��ʯ+� � �a�$���H���l� Ϳ�����ƿ'��K� �o�2�hϥϔ��ό� �ϰ�������F�k� .ߏ�R߳�v��ߚ��� ����1���U��y�<�QUICC0��b�t����1�����%���2&���u�!ROUTERv��R�d���!PCJ�OG����!1�92.168.0�.10��w�NAM�E !��!R�OBOTp�S_�CFG 1H��� �Au�to-start{ed�tFTP�������  2D��hz�� ��U��
//./ �v���/���/ �/�/�/�/�!?3?E? W?i?�/?�?�?�?�? �?�?���AO�?eO �/�O�O�O�O�?�O�O __+_NO�OJ_s_�_ �_�_�_
OO.OoB_ 'ovOKo]ooo�oP_>o �o�o�o�oo�o5 GYk}�_�_�_� �8o��1�C�U� $y��������ӏf� ��	��-�?���� �Ə���ϟ��� ��;�M�_�q���.� (���˯ݯ��P�b� t�����m��������� ǿٿ�����!�3�E� h��{ύϟϱ���� $�6�H�J�/�~�S�e� w߉ߛ�jϿ������� �*߬�=�O�a�s���YT_ERR �J5
���PDUS_IZ  ��^J�����>��WRD� ?t�� � guest}��%�7�I�[�m��$SCDMNGR�P 2Kt������V$��K�� 	P01�.14 8�� �  y����B�    ;������ ���߇����
 �������������~����C.g�R|���  �i  �  
��������� +��������
����l .r���"�l��� �m
d������_�GROU��L��� �	����07�EQUPD  d	պ�J�TYa �����TTP_AUTH 1M��� <!iPeOndany��6��Y!KARE�L:*��
-K�C///A/ VI�SION SETT�/v/�"�/�/ �/#�/�/
??Q?(?�:?�?^?p>�CTRL N����5��
�FFF9�E3�?�FRS�:DEFAULT��<FANUC� Web Server�:
���� �<kO}O�O�O�O�O���WR_CONFI�G O�� ��?��IDL_CP�U_PC@�B���7P�BHUM�IN(\��<TGNR_IO������P�NPT_SIM_�DOmVw[TPM�ODNTOLmV >�]_PRTY�X7R�TOLNK 1P����_o!o3oEo�Woio�RMASTE�lP��R�O_CFG�o�iUO��o�bCYCLE�o�d@_ASG 1Q����
 ko,>P bt����������sk�bNUM�����K@�`IPC�H�o��`RTRY�_CN@oR��bSGCRN����Q���1 �b�`�bR����Տ��$J23_�DSP_EN	�����OBPROqC�U�iJOGP�1SY@��8G�?�!�T�!�?*��POSRE�zVKANJI_�`��o_H�� ��T�L�6͕<����CL_LGP<��_���EYLOGG+IN�`���LANGUAGE� YF7RD ,w���LG��U�?�+���x� ������=P��'0���$ NMC:\�RSCH\00\���LN_DISP V��
������f��OC�R.RDzVT�A{�OGBOOK W
{��i��ii��X�����ǿٿ�����"��6	h�����e�?��G_BUFF 1%X�]��2	ա� ������������ !�N�E�W߄�{ߍߺ� �����������J�����DCS Z>r� =����^π+�ZE��������a�I�O 1[
{ ُ!� �!�1�C�U� i�y������������� ��	-AQcu@�������EfP/TM  �d�2 /ASew��� ����//+/=/�O/a/s/�/�/��S�EV����TYP�/??y͆��RS@"��×�F�L 1\
���� ��?�?�?�?�?�?�?�/?TP6��">>�NGNAM�ե��U`�UPS��GI�}�𑪅mA_LO{AD�G %��%DF_MOT�N���O�@MAXUALRM<��J��@sA�Q����WS ��@C �]m�-_���MPt2�7�^
{ رƭ	�!P�+ʠ�;_/��Rr�W�_�WU�W�_��R	o�_ o?o"ocoNoso�o�o �o�o�o�o�o�o; &Kq\�x�� �����#�I�4� m�P���|���Ǐ��� ֏��!��E�(�i�T� f�����ß��ӟ��� � �A�,�>�w�Z��� ����ѯ����د�� �O�2�s�^��������Ϳ���ܿ�'��BD�_LDXDISA�X@	��MEMO_{APR@E ?�+
 � *�~ϐπ�ϴ����������@I�SC 1_�+ ��IߨT��Q�c�� �߇��ߧ�����w�� ��>�)�b�t�[��� ��{����������:� ��I�[�/�������� ����o�����6!Z lS��s�� ��2�AS' �w����g���.//R/d/�_M?STR `�-w%�SCD 1am͠ L/�/H/�/�/?�/2? ?/?h?S?�?w?�?�? �?�?�?
O�?.OORO =OvOaO�O�O�O�O�O �O�O__<_'_L_r_ ]_�_�_�_�_�_�_o �_�_8o#o\oGo�oko �o�o�o�o�o�o�o" F1jUg�� �������B� -�f�Q���u�����ҏ�h/MKCFG �b�-㏕"LTA�RM_��cL�� σQ�N�><�METPUI�ǂ����)NDSP_CMNTh����|�  d�.���ς�ҟܔ|�POS�CF����PST�OL 1e'�4@�<#�
5�́5� E�S�1�S�U�g����� ��߯��ӯ���	�K� -�?���c�u�����|��SING_CHK�  ��;�ODA�Q,�f��Ç��D�EV 	L�	�MC:!�HSIZ�Eh��-��TAS�K %6�%$1�23456789� �Ϡ��TRIGw 1g�+ l6�%���ǃ�����8��p�YP[� ��EM_INF 1h3�� `)�AT&FV0E�0"ߙ�)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ������H������A���AI�q�,���|���� ���� ������J���n���� ��W�����������" ����X��/���� e������0� T;x�=�as ��/�,/c=/b/ �/A/�/�/�/�/� �?���^?p?#/ �?�/�?s?}/�?�?O �?6OHO�/lO?1?C? U?�Oy?�O�O3O _�?�D_�OU_z_a_�_�O�NITOR��G �?5�   	�EXEC1Ƀ�R2*�X3�X4�X5�X����V7�X8�X9Ƀ �RhBLd�RLd�RLd�R Ld
bLdbLd"bLd.b�Ld:bLdFbLc2Sh2�_h2kh2wh2�h2��h2�h2�h2�h2*�h3Sh3_h3�R��R_GRP_SV� 1in���(�����C?BPP��A4�>%��gY�>r���x�_D=R^��PL�_NAME !�6��p�!De�fault Pe�rsonalit�y (from �FD) �RR2�eq 1j)TUX�)TX��q��X dϏ8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������2'�П�����*� <�N�`�r��<���� ����ү�����,��>�P�b� �Rdr 1�o�y �\�, Ӗ3���� @oD�  ��?���➱?䰺��A'��6����;�	l�ʲ	 �xoJ������ �<; �"�� �(p�K�K ���K=*�J���J���JV��0�Z�����rτ���p@j�@T;f���f��ұ]��l��I��������������b���3��´  ��`�>����bϸ�z��Ꜧ�Ͽ�Jm��
�  B�H�˱]���q�	�� p�  �P�pQ�p��p| � Ъ�g���c�	�'� � ���I� �  {����:�È
�?È=���"�n����	�ВI  �n @B�cΤ�\��ۤ��q�y�o�yN���  '�������@2��@�c����/�C��}C�C�@ C�������
�AT�W�@<�P�R�%
h�B�b�A��j������:��Dz ۩��߹�����j���( �� -��C���'�7L�����q�Y������ �?�ff ���gy ����o�:a��
�>+�  PƱj�( ����7	���^|�?����xZ��p<
6b<���;܍�<����<� <�&Jσ�AI�ɳ+�|���?fff?I��?&�k�@�.���J<?�` �q�.�˴fɺ�/ ��5/����j/U/�/ y/�/�/�/�/�/?�/0?q��F�?l? ?�?/�?+)�?�?ؿE�� E�I�G+� F��?)O �?9O_OJO�OnO�Of�BL޳B�?_h�.� �O�O��%_�OL_�?m_ �?�__�_�_�_�_�
��h�Îg>���_Co�_goRodo��o�GA�ds�q�C��o�o�o|���ؠ$]Hq���D���pC���pCHmZZ7t���6q�q���ܶN'�3A�A��AR1AO��^?�$�?��K/�±
=ç�>����3�W�
=�#�W��e��9�����{�����<���(�B�u���=B0��?����	L���H�F�G����G��H�U`�E���C�+����I#�I���HD�F���E��RC�j�=��
I���@H�!H�(� E<YD0 q�$��H�3�l�W� ��{��������՟� ��2��V�A�z���w� ����ԯ������� �R�=�v�a������� �����߿��<�'� `�Kτ�oρϺϥ��� �����&��J�\�G� ��kߤߏ��߳����� ��"��F�1�j�U�� y������������0��T�?�Q����(����3/E��<��u������q3�8�����q�4Mgs&I�B+2D�a���{�^^	�������uP2P7Q4_A��M0bt��R�������/   � /�b/P/�/t/�/ *�a)_3/�/�/�% 1a?�/?;?M?_?q?  �?�/�?�?�?��?O 2 F��$�vGb�/�A���@�a�`�qC��C@��o�Ot���KF�� DzH@�� F?�P D���O�O�ys<O!_3_E_W_�i_s?���@@*pZ�422!u2~
 p_ �_�_�_	oo-o?oQo couo�o�o�o�o��Q� ��+��1���$MSKCFM�AP  �5� �6�Q�Q�"~�cONREL  
q3�bEXCFENB?wq
s1uXqFNC_�QtJOGOVLI�M?wdIpMrd�bK�EY?w�u�bR�UN�|�u�bS?FSPDTY�av<Ju3sSIGN?Qt�T1MOT�Nq��b_CE_GRP� 1p�5s\ r���j�����T��� �������<��`�� U���M���̟��🧟 �&�ݟJ��C���7� ������گ��������4�V�`TCOM_�CFG 1q}иVp�����
P�_A�RC_\r
jyU?AP_CPL��nt�NOCHECK {?{ 	 r��1�C�U�g�y� �ϝϯ���������	���({NO_WAI�T_L�	uM�NT�X�r{�[m�_7ERRY�2sy3� &�������r��c� ��T_M�O��t��,  {�t$�k�3�PARAuM��u{�	�`[���u?�� =9@�345678901��&���E�W�3� c�����{������������=�U�M_RSPACE� �Vv��$OD�RDSP���jxO�FFSET_CAsRTܿ�DIS���PEN_FIL�E� �q��c֮�OPTION_IO���PWORK 5v_�ms �P�(�R�Q
�j.j	C ��Hj&6$� �RG_DSBL  �5Js�\��RIENTTO>p9!C��PqfA� �UT_SIM_D�
r�b� V� LCT ww�bc���U)+$_PEXE�d&RATp �vju��p��2X�j)TU�X)TX�##X d-�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O?O�H2�/oO�O�O�O��O�O�O�O�O_]�< ^O;_M___q_�_�_�_ �_�_�_�_o���X��OU[�o(�꘯(���$o��, ��IpB` �@D�  Ua?��[cAa?p]a]�D�WcUa쪋l;�	l�mb�`�xJ�`�p���a�< ��`�� ��b��H(���H3k7HSM�5G�22G���Gp
��
��c�'|��CR�	>�>q�GsuaT��3���  �4 spBpyr  ]o�*S�B_����j�]��t�q� ��rna �,����6  ��P�Q�|N��M�,k���	'� �� ��I� �  ��%�=��ͭ���ba�	���I  �n @��~���Dp�������N	 W�  '!o�:q�pC	 C�@@sBq�t|��� m�
�!*�h@ߐ�n����*�B	 �A���p�G �-�qbz��P��t�_�������( �� -��恊�n�ڥ[A"]Ѻ�b4�'!5�(p? �?�ff� ��
����OZ�R*��85�z���>΁  	Pia��(5���@����ک�a�c�dF#?��5�x��*�<
6�b<߈;܍��<�ê<� <�&�o&�)��A�lcΐI�*�?f7ff?�?&c����@�.uJ<?�`��Yђ^� nd��]e��[g��Gǡd <����1��U�@�y� dߝ߯ߚ����߼�	� ��-������&��"�E�� E��G+� Fþ����� �������&��J�5��bB��AT�8�ђ ��0�6���>���J� n�7��[m�0���h��1��>��M�I
��@��A�[��C�-�)��?�A��� /�YĒ�a�Jp��vav`CH/�������}!@I��Y�'�3A��A�AR1AO��^?�$�?�����±
=���>����3�?W
=�#����+�e��ܒ������{����<�����.(�B�u���=B0������	��*H�F�G����G��H�U�`E���C�+��-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�?O �?3OOWOBOTO�OxO �O�O�O�O�O�O_/_ _S_>_w_b_�_�_�_ �_�_�_�_oo=o(o aoLo�o�o�o�o�o�o �o�o'$]H �l������ �#��G�2�k�V��� z���ŏ���ԏ��� 1��U�g�R���v��� ��ӟ�������-���(�������y�a����Q�<c�,!3�8�}���,!4Mgs����ɢ�IB+կ篴a���{���A�@/�e�S���w��P!�	P�������7��0ӯ�ϑ�R9�K�`��oχϓϥ�  ���χ����)��M� �����z���{߉ߛ���ߒߤ�������  )�G�q�_����2 F;�$�&Gb���n�a�[ZjM!C�s��@j/�A�S�=�F�� Dz��� F�P D��W����)������������x?���@U@
9�=�=���=��
  v������ �*<N`�*�P ���˨�1���$PARAM�_MENU ?�-�� � DEFP�ULSEl	W�AITTMOUT��RCV� �SHELL_W�RK.$CUR_oSTYL�,�OPT�/PTB�./("C�R_DECSN���,y/�/ �/�/�/�/�/?	??�-?V?Q?c?u?�?�U�SE_PROG �%�%�?�?�3C�CR�����7_HOST !�#!�44O�:T̰�?�PCO)ARC�O�;_�TIME�XB� � �GDEBU�GV@��3GINP?_FLMSK�O�IqT`��O�EPGAPe �L��#[CH�O^�HTYPE����?�?�_�_�_�_�_ oo'o9obo]ooo�o �o�o�o�o�o�o�o :5GY�}�� �������1��Z��EWORD ?}	7]	RS`�_	PNS�$斂JOE!>�TE�s@WVTRACEC�TL 1x-��� ������ɆDT Qy�-���D � ��,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾��� ������*�<�N�`� r����������� ��&�8�J�T�(�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_j� �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �_����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/�/"#�$PGTR�ACELEN  �#!  ���" �8&_U�P z���2g!o S!h 8!_CFG {g%#Q#"!x!�$J ��#|"DEFSPD� |�,!!J ��8 IN TRLW }�-" 8�%��!PE_CONF�I� ~g%��g!�$�%�$LI�D�#�-74GR�P 1�7Q!��#!A ���&�ff"!A+33D��� D]� C�À A@+6�!��" d�$�9�9*1*0� 	 +9�(�&�"�? ´	C�?�;B@3AO�?OIO3O�mO"!>�T?��
5�O�O�N�O =��=#�
�O _�O_J_5_n_Y_�O�}_�_y_�_�_�_  #Dzco" 
oBo �_Roxoco�o�o�o�o �o�o�o>)b�M��;
V7.10beta1�$�  A�E}�rӻ�A " ޼p?!G��q>˙��r��0�q̽ͻqBQ��qAA\�p�q�4�q�p�"�BȔ2�D�V�h�Bw��p�?�?)2{ ȏw�׏���4�� 1�j�U���y�����֟ ������0��T�?� x�c�������ү���� !o�,�ۯP�;�M��� q�����ο���ݿ� (��L�7�p�+9��sF@ �ɣͷϥ� g%������+�!6I� [߆������ߵߠ��� ������!��E�0�B� {�f���������� ���A�,�e�P��� t���������� ��=(aL^�� �����'9 $]�Ϛ��ϖ��� ����/<�5/`�r� �ߖߏ/>�/�/�/�/ �/?�/1??U?@?R? �?v?�?�?�?�?�?�? O-OOQO<OuO`O�O �O�O�O���O_�O)_ _M_8_q_\_n_�_�_ �_�_�_�_o�_7oIo t���o�o���o �o�o(/!L/^/p/�/ {*o������ ���A�,�e�P�b� ���������Ώ�� +�=�(�a�L���p��� ���Oߟ񟠟� �9� $�]�H���l�~����� ۯƯ���#�No`oro �on��o�o�o�oԿ ���8J\ng�� ��vϯϚ�������	� ��-��Q�<�u�`�r� �ߖ��ߺ������� ;�M�8�q�\������ ��z������%��I� 4�m�X���|������� ����:�L�^���Z ����������� $�6�H�Swb �������/ /=/(/a/L/�/p/�/ �/�/�/�/?�/'?? K?]?H?�?��?�?f? �?�?�?O�?5O OYO DO}OhO�O�O�O�O�O �O&8J4_F_�� ��_�_��_�_" 4-o�O*ocoNo�oro �o�o�o�o�o�o) M8q\��� ������7�"� [�m��?����R�Ǐ�� �֏�!��E�0�i� T���x��������_ $_V_ �2�l_~_�_������R�$PLID�_KNOW_M � �T������SV �v�U͠�U��
��.�ǟR�=��O�����mӣM_G�RP 1��!`0*u��T@ٰo�ҵ�
���Pзj�� `���!�J�_�W�i� {ύϟϱ��������Ϭ߱�MR�����T��s�w� s��ߠ� �߯߅��ߩ߻����� A���'����� ����������=�� �#���������}���ء��S��ST��1 �1��U# ���0�_ A .��, >Pb����� ���3(iL ^p������2*���<-/3/)/;/M/A4f/x/�/�/5�/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?MA/D  d#`�PARNUM � w�%OS+CH?J ME
�G`A8�Iͣ�EUPD`OrE�
a�OT_CMPa_��B@�P@'˥~TER_CHK'U���˪?R$_6[RqSl�¯��_MOA@�_�U_�_RE_RES_G ��>� oo8o+o\oOo�oso �o�o�o�o�o�o�o�W �\�_%�Ue  Baf�S� ��� �S0����SR0� �#��S�0>�]�b��S��0}������RV 1񈟥��rB@c]���t�(@c\�����D@c[��$���RTHR_ICNRl�DA��˥d,�oMASS9� ZM��MN8�k�MON_�QUEUE ����˦��x� RDN�PUbQN{�P[��E�ND���_ڙEXE�ڕ�@BE�ʟ��OPTIOǗ�[���PROGRAM %��%��ۏ�O~��TASK_IAD�0�OCFG ��tO��ŠDATA����Ϋ@��2 7�>�P�b�t���,��� ��ɿۿ�����#�5ϼG���INFOUӌ�������ϭϿ��� ������+�=�O�a� s߅ߗߩ߻�������h�^�jč� y�ġ?PDIT ��ίc���WERFL�
��
RGADJ7 �n�A�����?����@���IOR�ITY{�QV���M�PDSPH�����U�z����OTOE�y�1�R� (!AF4�E�P]���?!tcph����!ud��!�icm��ݏ6�X�Y_ȡ�R��ۡ)� *+/ ۠�W:F� j�������%7[B�*���PORT#�BC�۠����_CARTREP
�R� �SKSTAz��ZS�SAV���n�	�2500H863����r�$!�R�
���q�n�}/�/��'� URGE�Bl��rYWF� DO{��rUVWV��$�A�W�RUP_DELA�Y �R��$R_'HOTk��%O]?��$R_NORMA�Lk�L?�?p6SEM�I?�?�?3AQSKkIP!�n�l#x 	1/+O+ ORO dOvO9Hn��O�G�O�O �O�O�O_�O_D_V_ h_._�_z_�_�_�_�_ �_
o�_.o@oRoovo do�o�o�o�o�o�o�o *<Lr`����n��$RCV�TM�����pDkCR!�LЈq�B��C*J��C$�>�$ �>5?-;��0�4M¹�O�������������~��9On�Y�<
6�b<߈;܍��>u.�?!<�&{�b�ˏ ݏ��8�����,�>� P�b�t���������Ο ���ݟ��:�%�7� p�S������ʯܯ�  ��$�6�H�Z�l�~� ������ƿ���տ� ��2�D�'�h�zϽ��� ����������
��.� @�R�d�Oψߚ߅߾� ����������<�N� ��r��������� ����&�8�#�\�G� ����}����������� S�4FXj|� �������� 0T?x�u� ���'//,/>/ P/b/t/�/�/�/�/�/ �/�?�/(??L?7? p?�?e?�?�?��?�?  OO$O6OHOZOlO~O �O�O�?�?�O�O�O�O  __D_V_9_z_�_�? �_�_�_�_�_
oo.o�@oRodovo�X�qGN_ATC 1��� AT&�FV0E/� �ATDP/6/9�/2/9�hAT�A�n,AT�%G1%B960�/�+++�o,��aH,�qIO_TYPE  �u��sn_�oREFP�OS1 1�P{O x�o�Xh_ �d_�����K� 6�o�
���.���R�����{{2 1�P{ ���؏V�ԏz����q3 1��$�6�p���ٟ���S4 1�����˟���n���>%�S5 1�<�N��`�����<���S6 1�ѯ���/������ѿO�S7 1� f�x���ĿB�-�f��S8 1������Y�������y�SMA�SK 1�P  q
9�G��XNOM����a~߈ӁqMO�TE  h�~t��_?CFG �������рrPL_RAN�G�ћQ��POWE/R ��e���SM_DRYPR/G %i�%��J���TART ��
�X�UME_PR�O'�9��~t_EX�EC_ENB  y�e��GSPD��p����c��TDB����RM��MT_�!�T���`OB�OT_NAME �i���iOB�_ORD_NUM� ?
�\q�H863  ��T��������bP�C_TIMEOU�T�� x�`S23�2��1��k L�TEACH ?PENDAN ��ƅ�}���`M�aintenance Cons�R�}�m
"{�dKC�L/Cg��Z ���n� No Use}�	��*�NPO��х����(CH_Lf�������	�~mMAVAIL���{��ՙ�SPA�CE1 2��| d��(>��&����p��M,8�?�ep/eT/�/ �/�/�/�W//,/>/ �/b/�/v?�?Z?�/�? �9�e�a�=??,?>? �?b?�?vO�OZO�?�OP�O�Os�2�/ O*O<O�O`O�O�_�_@u_�_�_�_�_[3_ #_5_G_Y_o}_�_�o��o�o�o�o[4 .o@oRodovo$�o�o ����"�	�7�[5K]o��A�� ��	�̏�?�&�T�[6h�z�������^� ԏ���&��;�\�C�q�[7��������͟ {���"�C��X�y�`���[8����Ưد ꯘ��0�?�`�#�u���}ϫ�[G �Ni� �ϋ
G� ����$�6�H� Z�l�~ߐ��8 ǳ�� ���߈��d(�� �M�_�q����� �������?���2�%� 7�e�w����������� ���������!�RE� W�����������?Q `�� @0��� �rz	�V_� ����
/L/^/|/ 2/d/�/�/�/�/�/�/ ?�/�/�/*?l?~?�? R?�?�?�?�?�?�?�?�2O�?
��O[_MODE  ��^�IS ���vO,*ϲ�O-_���	M_v_#dCWOR�K_AD�M-���%aR  ���ϰ�P{_�P_INT�VAL�@����JR_OPTION�V� �EBpVAT_GRP 2���w�(y_Ho �e_vo�o�oYo �o�o�o�o�o*< �bOoNDpw�� ����	���?� Q�c�u�����/���Ϗ Ꮳ����)�;���_� q���������O�ɟ� ��՟7�I�[�m�/� ������ǯٯ믁�� !�3���C�i�{���O� ��ÿտ���ϡ�/� A�S�e�'ωϛϭ�o� ��������+�=��� a�s߅�Gߕ߻����� ����'�9�K�]��� �����y�����������5�G�Y��E�$�SCAN_TIM�AYuew�R ��(�#((�<}0.aaP%aP
Tq>��Q��o�����O+O2/��:	d/JaR��WY��^���^R^	�r  P��w� �  8�P��	�D�� GYk}���������Qp/@/R//)P�;�o\T��Qp�g-�t�_D�iKT��[  � lv%������/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OWW�#�O�O �O�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_olO~Od+ No`oro�o�o�o�o�o �o�o&8J\ n������u�  0�"0g�/�-� ?�Q�c�u��������� Ϗ����)�;�M� _�q�����$o��˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�����Do�� ������ҿ����� ,�>�P�b�tφϘϪπ����������w
�  58�J�\�n߀ߒ� �կ���������	�� -�?�Q�c�u������ ��-���� � �2�D�V�h�z�����������������;�& ��%�	123456{78�" 	��/� `r�������� (:L^p���� ���� //$/6/ H/Z/l/~/��/�/�/ �/�/�/? ?2?D?V? h?�/�?�?�?�?�?�? �?
OO.O@Oo?dOvO �O�O�O�O�O�O�O_ _*_YON_`_r_�_�_ �_�_�_�_�_ooC_ 8oJo\ono�o�o�o�o �o�o�oo"4F Xj|���������	��s3��E�W�{�Cz  �Bp��   ���2���z�$SC�R_GRP 1��(�U8(�\x�^ @�  �	!�	 ׃���"�$�  ��-��+��R�w�7���D~������#����O����M-10iA 8909905 Ŗ5 ?M61C >4���Jׁ
� � ��0�����#�1�	"�z�������¯Ҭ ���c� ��O�8�J�������!�����ֿ��B�y���������9A��$�  @��<�D �R�?��d���Hy��u�O���F@ F�`�§�ʿ�϶��� ����%��I�4�m��<�l߃ߕߧ߹�B���\����1��U� @�R��v������ �����;���*<�=�
F���?�d�<�>g7�����@�:�n�� B���З�Й���EL_DE�FAULT  ~����B��MIPOWE?RFL  �$�1 WFDO� $��ERVENT 1������"�pL!DU�M_EIP��8���j!AF_IN�E �=�!FT$���!��4� ��[!RPC_MAIN\�>�J�nVIS�w=���!TMP�PU��	d��?/!
PMON_�PROXY@/�e ./�/"Y/�fz/�/�!RDM_SR�V�/�	g�/#?!�R C?�h?o?!%
pM�/�i^?�?�!RLSYNC̼?8�8�?O!gROS�.L�4�? SO"wO�#DOVO�O�O �O�O�O_�O1_�OU_ _._@_�_d_v_�_�_ �_�_o�_?oocoi�ICE_KL ?�%y (%S?VCPRG1ho8��e���o�m3�o�o�`4 �`5(-�`6PU�`7x}�`H���l9��{�d :?��a�o��a�oE� �a�om��a���aB ���aj叟a���a �5��a�]��a��� �a3����a[�՟�a�� ���a��%��aӏM��a ��u��a#����aK�ů �as���a��mob�` �o�`8�}�w������� ɿ���ؿ���5�G� 2�k�VϏ�zϳϞ��� �������1��U�@� y�dߝ߯ߚ��߾��� ����?�*�Q�u�`� ����������� �;�&�_�J���n������������sj_D�EV y	��MC:��_]OUT"�,REC 1��Z� d   � 	�     ��@���� ��A�����
 �PSD#6� r��O� �J� �� `�� �Z�T{� �� *N�  +X- � UI- �- !- � ��X�YZ�PSJU;4 �? � (�  �� ��R ��U� E- � �1/e/�l4�/���� X� (@,/>/P/�/�/�""4�� =�!� � ��  ?"S1��'!��/���("- � �\?�?$=�=�?�?�? "OOFO4OjO|O^O�O �O�O�O�O�O�O_ _ _T_B_x_f_�_�_�_ �_�_�_�_oooPo >oto�oho�o�o�o�o �o�o(
L:\@�p���w, ����4�"�X�F� |���p�����֏ď� ���0��@�f�T��� x�����ҟ�Ɵ��� ,��<�b�P���h�z� �����ί��(�:� �^�L�n�p������� ܿ�п� �6�$�Z� H�jϐ�rϴϢ����� �����2�D�&�h�V� ��z߰ߞ��������� ��
�@�.�d�R��Z�jV 1�w P����j 
ß� ����
T�YPEVFZN_CFG ��5�d�4�G�RP 1�A�c� ,B� A� D�;� B��� � B4RB{21HELL:��(
��?���<%RS'!�� H3lW�{�� ����2V�h������%@w����#!�1������7�2��0d����HK ;1��� �k/ f/x/�/�/�/�/�/�/ �/??C?>?P?b?�?��?�?�?��OMM �����?��FTOV_ENB ���+��HOW_REG_�UIO��IMWA�ITB�JKOU�T;F��LITIM�;E���OVAL|[OMC_UNITC��F+�MON_AL�IAS ?e�9 ( he��_&_ 8_J_\_B_�_�_�_ �_j_�_�_oo+o�_ Ooaoso�o�oBo�o�o �o�o�o'9K] n����t� ��#�5��Y�k�}� ����L�ŏ׏���� ��1�C�U�g������ ����ӟ~���	��-� ?��c�u�������V� ϯ������;�M� _�q��������˿ݿ ����%�7�I���m� ϑϣϵ�`������� ߺ�3�E�W�i�{�&� �߱������ߒ��� /�A�S���w���� X����������=� O�a�s���0������� ������'9K] ����b�� �#�GYk} �:������ /1/C/U/ /f/�/�/ �/�/l/�/�/	??-? �/Q?c?u?�?�?D?�? �?�?�?O�?)O;OMO _O
O�O�O�O�O�OvO��O__%_7_�C�$�SMON_DEF�PRO ����`Q �*SYSTEM*  d=OU�RECALL ?�}`Y ( �}�
xyzrate� 61 *.* �virt:\tm�pback\�P=�>192.168�.4�P46:1652 �Q�_�_�_�K�}�W�^5012� �_�_couo�ob9�copy frs�:orderfil.dat�\*o<a��o�o�ol0�bmdb:�_�o<a�obt�c6�o�hemp>:8188 W�t��.�v*.d� �~�`�r���e�Y+� =�O�����o)o҂ ��ҏc�u����o�o5 �wٟ���"���y`ҟc�u����4x��:�Q�_;�S�U����.
� }5��a���� �wׯh�z������:� կ���
����A�ӿ d�vψϛ�.�;�ѯ�� �����ϼ�O�`�r� �ߗ���2�Ϳ����� �'���K�\�n��� ��8����������#� ��G��j�|����_3��E�W��������Gg2244?o��bt� �߫�4�5���� "�5�bt��� ����:U��
/� ����h/z//�� 1/C/U/�/�/
?/j2T��/�/c?u?�?� �567�?�?�?" �?58�?bOtO�O��?��Nb60 WO�O�O �O��O�I�O`_r_�_ �/��;_M_�_�_o? '?�T�_�_couo�o�? �?5O�G�o�o�oO"O �o�H�obt���/ �/KtV���/� �>`�h�z���o�o :����
���A�ӏd�v������$S�NPX_ASG �1�������� P 0� '%R[?1]@1.1����?���%֟��&� 	��\�?�f���u��� �����ϯ��"��F� )�;�|�_�������ֿ ��˿���B�%�f� I�[Ϝ�Ϧ��ϵ��� ����,��6�b�E߆� i�{߼ߟ�������� ���L�/�V��e�� �����������6� �+�l�O�v������� ��������2V 9K�o���� ���&R5v Yk�����/ ��<//F/r/U/�/ y/�/�/�/�/?�/&? 	??\???f?�?u?�? �?�?�?�?�?"OOFO )O;O|O_O�O�O�O�O �O�O_�O_B_%_f_ I_[_�__�_�_�_�_ �_�_,oo6oboEo�o io{o�o�o�o�o�o �oL/V�e� �������6� �+�l�O�v��������PARAM ������ �	U��P�����OFT_KB_CFG  ⃱����PIN_SIM  ���C�U�g������RVQSTP/_DSB,�򂣟|����SR �/��� &  AR������TOP__ON_ERސ����PTN �/�@�A�	�RING_PR�M� ��VDT_GRP 1�ˉ�  	������ ������Я����� *�Q�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߣߠ߲������� ����0�B�i�f�x� ������������� /�,�>�P�b�t����� ����������( :L^p���� ��� $6H Z�~����� ��/ /G/D/V/h/ z/�/�/�/�/�/�/? 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�__\_��VPRG_�COUNT��8@���RENBU��U�M�S��__UPD� 1�/�8  
s_�oo*oSoNo `oro�o�o�o�o�o�o �o+&8Jsn �������� �"�K�F�X�j����� ����ۏ֏���#�� 0�B�k�f�x������� ��ҟ������C�>� P�b���������ӯί������UYSDOEBUG�P�P�)��d�YH�SP_PA�SS�UB?Z�L�OG ��U��S)�#�0�  ���Q)�
MC:�\��6���_MPC ���U���Qñ8�� �Q�SAV ������ǲ%��ηSV;�TEM_TIME 1��[W (�P"�T!y��ؿT1SVGUNYS�P�U'�U����ASK_OPTICON�P�U�Q�Q���BCCFG Ì�[u� n�X�G�`a�gZo��߃ߕ��� ��������:�%�^� p�[���������  �����6�!�Z�E�~�@i���������%��� ����&8��nY �}�?��ԫ � �(L:p^ �������/  /6/$/F/l/Z/�/~/ �/�/�/�/�/�/�/2? 8 F?X?v?�?�?? �?�?�?�?�?O*O<O 
O`ONO�OrO�O�O�O �O�O_�O&__J_8_ n_\_~_�_�_�_�_�_ �_o�_ o"o4ojoXo �oD?�o�o�o�o�oxo .TBx�� j������� �,�b�P���t����� Ώ��ޏ��(��L� :�p�^�������ʟ�� o��6�H�Z�؟ ~�l�������د��� ʯ ��D�2�h�V�x� z���¿���Կ
��� .��>�d�Rψ�vϬ� ���Ͼ�������*�� N��f�xߖߨߺ�8� ��������8�J�\� *��n�������� ����"��F�4�j�X� ��|����������� ��0@BT�x �d����� >,Ntb��� ���/�(//8/ :/L/�/p/�/�/�/�/ �/�/�/$??H?6?l? Z?�?~?�?�?�?�?�? O�&O8OVOhOzO�? �O�O�O�O�O�O
__ �O@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<o^o�oro�o�o�o �o�o�o J8 n$O�����X ���4�"�X�B�v���$TBCSG_�GRP 2�B���  ��v� 
 ?�  ������׏����叀��1��U�g�z����~��d, ����?v�	 HC���d�>����e�CL  B���Пܘ���\)>��Y  A�ܟ$�3B�g�B�Bl�i��X�ɼ���X��  �D	J���r�����C ����үܬ���D�@v�=�W�j�}�H�Z� ��ſ����������v�	V3.�00��	m61c�	*X�P�u�Lg�p�>���v�(:��� ��p͟�  O����p������z�JCFG ȖB��� ����������=��=�c�q�K�qߗ߂� �ߦ��������'�� $�]�H��l����� ��������#��G�2� k�V���z��������� �����p*<N ���l����� ��#5GY} h����v�b�� >�// /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?d?R?t?v?�? �?�?�?�?O�?*OO :O`ONO�OrO�O�O� �O�O�O_&__J_8_ n_\_�_�_�_�_�_�_ �_�_�_oFo4ojo|o �o�oZo�o�o�o�o�o �oB0fT�x �������,� �P�>�`�b�t����� Ώ�������&�L� �Od�v���2�����ȟ ʟܟ� �6�$�Z�l� ~���N�����دƯ� � �2��B�h�V��� z�����Կ¿���� .��R�@�v�dϚψ� ���Ͼ�������<� *�L�N�`ߖ߄ߺߨ� ���ߚ�������\� J��n������� ���"���2�X�F�|� j��������������� .TBxf� ������ >,bP�t�� ���/�(//8/ :/L/�/�ߚ/�/�/h/ �/�/�/$??H?6?l? Z?�?�?�?�?�?�?�? O�?ODOVOhO"O4O �O�O�O�O�O�O
_�O _@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<oro`o�o�o�o�o �o�o�o&�/>P �/������ ���4�F�X��(� ��|�����֏���� Ə0��@�B�T���x� ����ҟ������,� �P�>�t�b������� ��������:�(� ^�L�n�������2d �����̿�$�Z�H� ~�lϢϐ��������� �� ��0�2�D�zߌ� �߰�j���������� 
�,�.�@�v�d��� �����������<� *�`�N���r������� ������&J\ �t��B��� ���F4j| ��^����/��  2 6# �6&J/6"�$TB�JOP_GRP �2���?  ?�X,i#��p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�x�'�!�!>���
5�59>�0+1�33=�CL� �fff?+0?�ffB� J1�%Y?d7�.���/>��2�\)?0�5����;��hCY� ��  @� �!B� � A�P?�?�3EC�  D�!�,�0�*BOߦ?�3JB���
:���Bl�0��0�$�1�?O6!?Aə�AДC�1sD�G6�=q�E�6O0�p��B�Q�;�A�� �ٙ�@L3D	��@�@__�O�O>BÏ\JU�OHH�1ts}�A@33@?1� C�� �@�_�_&_8_>��D�UV_0��LP�Q30<{�zR� @�0�V�P!o3o �_<oRifoPo^o�o�o �oRo�o�o�o�oM (�ol�p~���p4�6&�q5	�V3.00�#m761c�$*(��$�1!6�A� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,IR�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^S@;Q��|8�E`rz@/&�8�6&�<��1�w�^$ES�TPARS  �*({ _#HR��AB_LE 1�p+Z�6#|�Q� � 1�|��|�|�5'=!|�	�|�
|�|�˕6!�|�|�|���RDI��z!ʟܟ� ��$���O������ ¯ԯ�����S��x# V���˿ݿ��� %�7�I�[�m�ϑϣ� �����������U-�� ��ĜP�9�K�]�o���-�?�Q�c�u���6�N�UM  �*z!� >  Ȑ�����_CFG ������!@b IMEBF_TT����x#��a�VER��b�w�a�R 1�p+
' (3�6"1 ��  6!����������  �9�$�:�H�Z�l�~� ���������������^$��_��@x�
�b MI_CHAN�m� x� kDBGLV;0o�x�a!n �ETHERAD �?�� �y��$"�\&n ROUmT��!p*!�*�SNMASK��x#�255.�h�fx^$OOL�OFS_DI���[ՠ	ORQCTRL �p+;/�� �/+/=/O/a/s/�/ �/�/�/�/��/�/�/�!?��PE_DET�AI��PON_�SVOFF�33P_MON �H��v�2-9STRTC_HK ����42VTCOMPA�Ta8�24:0FPR�OG %�%�CA)&O�3ISP�LAY��L:_IN�ST_MP GL�7YDUS���?�2L�CK�LPKQUIC�KMEt �O�2SC�RE�@�
tps��2�A�@�I���@_Y���9�	S�R_GRP 1Ҿ� ��� \�l_zZg_�_�_�_�_�_�^�^�oj�Q'O Do/ohoSe��oo�o �o�o�o�o�o! WE{i�������	1234�567��!���X��E1�V[
 �}�ipnl/a�g?en.htmno���������ȏ~�P�anel setup̌}�?��0�B�T�f� ��񏞟 ��ԟ���o���� @�R�d�v������#� Я�����*���ϯ ůr���������̿C� �g��&�8�J�\�n� ����϶��������� uϣϙ�F�X�j�|ߎ� �����;��������0�B��*NUALR�Mb@G ?�� [���������� �� ��%�C�I�z�m�������v�SEV � ����t�E?CFG Ձ=]�/BaA$   B�/D
 ��/C� Wi{�����@�� PRց;C �To\o�I�6?K0(%����0 �����//;/ &/L/q/\/�/�/�/lƇD �Q�/I_��@HIST 1׾�9  ( � ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1?v?�?�?ά?�� >?P=962c?�?
OO.O�?�?�136�?|O�O�O�O AOSOeO�O__0_�H M___q_�_�_�_�_H_ �_�_oo%o7o�_[o moo�o�o�oDo�o�o@�o!3E ��a 81�ou����� �o���)�;�M�� q���������ˏZ�l� ��%�7�I�[��� ������ǟٟh���� !�3�E�W�������� ��ïկ�v���/� A�S�e�Pb������ ѿ������+�=�O� a�s�ϗϩϻ����� ��ߒ�'�9�K�]�o� ��ߥ߷��������� ��#�5�G�Y�k�}�� ������������� 1�C�U�g�y���v��� ��������	�? Qcu��(�� ��)�M_ q���6��� //%/�I/[/m// �/�/�/D/�/�/�/? !?3?�/W?i?{?�?�? �?�����?�?OO/O AOD?eOwO�O�O�O�O NO`O�O__+_=_O_ �Os_�_�_�_�_�_\_ �_oo'o9oKo�_�_ �o�o�o�o�o�ojo�o #5GY�o}������?��$�UI_PANED�ATA 1������  	�}�0�B�0T�f�x��� )���� mt�ۏ����#�5� ��Y�@�}���v����� ן�������1��U�pg�N������ �1��Ïȯگ���� "�u�F���X�|����� ��Ŀֿ=������ 0�T�;�x�_ϜϮϕπ�Ϲ������,ߟ� M��j�o߁ߓߥ߷� �����`��#�5�G� Y�k��ߏ������ ��������C�*�g� y�`���������F�X� 	-?Qc��� �߫���� ~;"_F��| �����/�7/ I/0/m/�����/�/�/ �/�/�/P/!?3?�W? i?{?�?�?�??�?�? �?O�?/OOSOeOLO �OpO�O�O�O�O�O_ z/�/J?O_a_s_�_�_ �_�O�_@?�_oo'o 9oKo�_oo�oho�o�o �o�o�o�o�o#
G Y@}d��&_8_ ����1�C��g� �_��������ӏ��� ^���?�&�c�u�\� ������ϟ���ڟ� )��M��������� ��˯ݯ0�����7� I�[�m���������� ٿ�ҿ���3�E�,� i�Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#��� ���� ��$�6��Z� A�~�e�w������ �����2��V�h�O������v�p��$UI�_PANELIN�K 1�v��  � � ��}1234?567890���� 	-?G ���o �����a��@#5G�	����4p&���  R� ����Z��$/ 6/H/Z/l/~//�/�/ �/�/�/�/�/
?2?D? V?h?z??$?�?�?�? �?�?
O�?.O@OROdO vO�O O�O�O�O�O�O _�O�O<_N_`_r_�_�_�0,���_�X�_ �_�_ o2ooVohoKo �ooo�o�o�o�o�o�o ��,>r}��� �������� �/�A�S�e�w���� ����я���tv�z� ���=�O�a�s��� ����0S��ӟ���	� �-���Q�c�u����� ��:�ϯ����)� ��M�_�q��������� H�ݿ���%�7�ƿ [�m�ϑϣϵ�D��� �����!�3�Eߴ_i� {�
�߂����߸��� ���/��S�e�H�� ��~��R~'�'�a� �:�L�^�p������� �������� ��6 HZl~���#� 5��� 2D�� hz�����c �
//./@/R/�v/ �/�/�/�/�/_/�/? ?*?<?N?`?�/�?�? �?�?�?�?m?OO&O 8OJO\O�?�O�O�O�O �O�O�O[�_��4_F_ )_j_|___�_�_�_�_ �_�_o�_0ooTofo ��o��o��o�o�o ,>1bt� ���K���� (�:����{O���� ��ʏ܏�uO�$�6� H�Z�l���������Ɵ ؟����� �2�D�V� h�z�	�����¯ԯ� �����.�@�R�d�v� �������п���� ��*�<�N�`�rτ��O �Ϻ�Io��������� 8�J�-�n߀�cߤ߇� ���߽����o1�o X��o|�������� �����0�B�T�f� �������������S� e�w�,>Pbt� �'���� �:L^p��# ���� //$/� H/Z/l/~/�/�/1/�/ �/�/�/? ?�/D?V? h?z?�?�?�???�?�? �?
OO.O��ROdO�� �OkO�O�O�O�O�O�O _�O<_N_1_r_�_g_��_7OM�m�$�UI_QUICK�MEN  ���_AobR�ESTORE 1��  �|��Rto�o�im�o�o�o�o �o:L^p�%� �����o��� �Z�l�~�����E�Ə ؏���� �ÏD�V� h�z���7�������/� ��
��.�@��d�v� ������O�Я���� �ßͯ7�I���m��� ����̿޿����&� 8�J��nπϒϤ϶� a�������Y�"�4�F� X�j�ߎߠ߲����� �ߋ���0�B�T�goSCRE`?#mu1sco`Wu2��3��4��U5��6��7��8��bUSERq�v��Tp���ks����4���5��6��7��8���`NDO_CFoG �#k  n`� `PDATE� ���N�onebSEUFRAME  �T�A�n�RTOL_�ABRTy�l��E�NB����GRP �1�ci/aCz  A�����Q�� $6HRd���`U�����MSKG  �����Nv�%�U�%���b�VISCAND_wMAX�I���FAIL_IM)G� �PݗP#���IMREGNUMr�
,[SIZ��n`�A�,VO�NTMOU���@���2��a���a�����FR:\ �� MC:\ޚ\LOG�B@F� !�'/!+/�O/�Uz M�CV�8#UD1&r&EX{+�S�P�PO64_��0n'fn6PO��CLIb�*�#V����,f@�'�/� �=	�(SZV�.�;���'WAI�/STAT ���B�P@/�?�?�:$�?��?��2DWP  ��P G@+b=��� H�O�_JMPERRw 1�#k
  ��2345678901dF�ψO{O�O�O �O�O�O_�O*__N_�A_S_�_
� MLO�Wc>
 �_TI�=�'MPH?ASE  ��F���PSHIFT֗1 9�]@< �\�Do�U#oIo�oYo ko�o�o�o�o�o�o�o 6lCU�y ����� ��	��V�-�e2����	�VSFT1�2	uVM�� �5�1�G� ���%A� W B8̀̀�@ pكӁ˂�у��z�#ME@�?�{��!�c>&%�aM1��k�0�{ �$`0T?DINEND���\�O� �z����Sp��w��P���ϜRELE�Q��Y����\�_ACTIV���:�R�A �`�e���e�:�RD� ����YBOX ��9�د�6��02����190�.0.�83���254��QF�	 �X�j��1��robo�t���   �p�૿�5pc��̿�����7���x��-�f�ZABC�����,]@U��2ʿ� eϢωϛϭϿ�����  ���V�=�z�a�s�$��E�Z��1�Ѧ