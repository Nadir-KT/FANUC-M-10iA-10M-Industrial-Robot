��   I�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��ETH_FLT�R.� $� �  �FT�P_CTRL.� @ $LOG�_8	�CMO>�$DNLD_FI�LTE� � SUB�DIRCAP��� HO��NT.� 4� H_NAM�E !AD�DRTYPA H_LENGTH'� �z +LS� D $R�OBOTIG P�EER^� MAS�KMRU~OM�GDEV#� R�DM*�DIS�ABL&� T�CPIG/ 3 $ARPSIZ&�_IPF'W_�MC��F_IN�� FA~LASS�s�HO_� IN{FO��TELKG PV�b�	 WORD  �$ACCESS�_LVL?TIM�EOUTuORT� � �ICEUS�=    �$�#  �����!�� � � VIRTUAL�/�!'0 ��%
���F����� �"�%�v��+ ��F���$�� �-2%;��SHARED �1�)  P!!�!�?���!|?�? �?�?�?O�?%O�?1O OZOOBO�OfO�O�O �O�O_�O�OE__i_ ,_�_P_�_t_�_�_�_ o�_/o�_SooLo�o xo�opo�o�o�o�o �o*Os6�Z �~�����9� �]� ���D�V���z� ۏ����#���Y��H�}�@���)7z _L�IST 1=x/!1.ܒ0��d��ە1�d�2551.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I����o�������O�6���8�`����� �$� ��-� ���-� �&P�%��&!Ò�)�0�H!� ���rj3_tpd����! � �!!K�C� e�0ٙ��&W�!Cm ��w߉�S�?!CON� ��z1�=�smon��W�