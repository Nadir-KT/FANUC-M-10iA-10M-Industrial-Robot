��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �
  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�H UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2F�G1_�3�B�2iG�XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1G ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�0@� �zsa�!ip;G0� � 
$WARNM�0f�!,P� ܁s�pNST� CO�RN�"a1FLTR^�uTRAT� T�p; H0ACCa1�p��{�ORI
`l"S={RT0_S�BְqHG,I1 E[ Tp�"3I9�CTY�D,P*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7ʳ�8��94���CO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS���}Aw��"�@&�wCP_*0OFSzRw @� RO_K8̨��aIT�3��NO�M_�0�1ĥ3u�qPT �� �$���AxP��K}EX �� �0g0I01��p��
$TFa��C$M�D3��TO�3�0U�� �� �H�w2�C1|�EΡg0�wE{vF�vF�40C�Pp@�a2 
P$�A`PU�3N1)#�dR*�AX�!sD�ETAI�3BUFpV�p@1 |�p�۶�pPIdT� PP[�MZ�Mg�Ͱj�}F[�SIMQSI �"0��A.���nQ��lw' Tp|zM��P��B�FACTrbHPEW7�P1Ӡ��vv��MCd� ��$*1JB�p<�*1DECHښ�H��(�c�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF4P��� &k�Bv�u�cu� �aE�� !2��+�MQ��E�SIZ�3�����T��P�����aRSINF�����kq�� ������LX������F�CRCMu�3CClpG��p���O}�� �b�1�������2�V�DxIC��C���r��`��P��{� EV ��zF_��F�pNB0�?������A�! �r�Rx�� ��V�lp�2��aR�t��,�g�rRTx #�5�5"2��uA�R���`CX�$LG�p��B�1 `s�P�tB�aA�0{�У+0R���tME�`!BupCfrRA 3tAZ��h��pc�OT�FC�b�`�`FNp���1��ADI+�a%��b �{��p$�pSp�c�`aS�P��a,QMP6䒁`Y�3��M'�pUt��aU  $>�TITO1�S�S�!���$�"0�DBPX�WO��!��$cSK��2p�DB��"�"@�PR8�� 
� ���# �>�q1$��$��+�L9$?(�V�R%@?R4C&_?�R4ENE��'4~?�A
�!RE�pY2�(H �OSn��#$L�3$$3�R��;3�MVOk_9D@!V�ROScrr��w�S���CRIGGER2FPA�S��7�ETURN0B�cM[R_��TUː[��0EWM%���G1N>`��RLA���E�ݡ�P�&$PD�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWAY�RMO#�aw!��DCS_)  `IS#� ��� �s3S�AQ汯  4Rx�ZSW�AQ�p�@1U9W��cTNTV)�5RV
a���|c�éWƃ¤�JB��x0��SAsFEۥ�V_SV�b�EXCLUU�;�N�ONL��cYg��~az�OT�a{�HI�_V? ��R, M�_G *�0� ��_z��2� �qQSGO  +�rƐm@�A@�c~b���w@��V�i|�b�fANNUNx0,�$�dIDY�UABc�@Sp�i�a+ �j�f��!�pOGIx2,���$F�b�$ѐO�T�@A $DUMMY��Ft��Ft�±� 6U- ` !�HE�|s���~bc�B@ SUFFmI��4PCA��Gs5Cw6dr�!M�SWU. 8!�KgEYI��5�TM�10�s�qoA�vINޱ��D, / D��H7OST�P!4����<���<�°<��p<�E�M'���Z�� SBL�� UL��0  ��	����DT��01 � $|��9USAMPL�@��/���決�$ I@|갯 $SUBӄ���w0QS�����#��SAV�����c�S< X9�`�fP$�0E!�� YN_B�#2 M0�`DI�d�pO|��m��#$F�R_I�C� �ENC2s_Sd3  ��< 3�9���� cgp����4�"��2�A9��ޖ5���`ǻ�@Q@K&D-!�a�AVER�q��λ�DSP
���PC�_�q��"�|�ܣ�V7ALU3�HE�(��M�IP)���OP5Pm �TH�*�D�S" T�/�Fb�B;�d����d ��g����16 H(rLL_DUǀ�a�@��0k���֠OT�"U��/���R_N_OAUTO70�C$}�x�~�@s��*|�C� ��C� 2��w�L�� 8/H *��L� � ��Բ@sv��`� �� � ����Xq��cq���q��T�q��7��8��9���0���1�1 �1�-�1:�1G�1T�1*a�1n�2|�2��U2 �2-�2:�2G�U2T�2a�2n�3|ʥ3�3� �3-�3�:�3G�3T�3a�3�n�4|����9� <���z�ΓKI`����H硵BaFEq@�{@: ,��&a?g P_P?��>�����E�@��v��QQ��;fp$T�P�$VARI�����,�UP2Q`< W�߃TD��g�����`��������BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P�"�Fl@``>Gt ;��6����ST����T��M ����0	��i���F� ��������kRt ����FORCEUP�b^܂FLUS
pH(�N��� ��6bD_CM�@E�7N� (��v�P��REM� F a��@j���
�K�	N���EFF�/���@IN�QO�V��OVA�	TgROV DT)��DTMX:e � P:/��Pq�vXpCLN _�p��@d ��	_|��_T: T�|�&PA�QDI���1��0�&Y0RQm�_+qH�2��M���CL�d#��RIV{�ϓN"EAmR/�IO�PCPd��BR��CM�@�N 1b 3GCLF��!DY�(��a6�#5T�DG���8� �%�FSS� )��? P(q1�1��`_1"811�E�C13D;5D6�GSRA���@�����PW�ON2EBUG�S�2���g�ϐ_E A ���@a �TER�M�5B�5��'ORIw�0C�5 ��SM_-`���0D��6�0A�9E�5�߹�UP��Fg� -QϒA�P|�3�@B$SEGGJv� EL�UUSEPNFI��pBx��1x@��4>DC$UF�P��$���Q�@C���G�0T�����SwNSTj�PATۡ<g��APTHJ�A�E*�Z%qB\`F�{E���F�q�pARxPY�aS�HFT͢qA�AX_�SHOR$�>��6 �@$GqPE���O#VR���aZPI@P@$�U?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi� [Y)��G�@R��i�e԰�i�R�!P�uAScYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C�%UaP���P���WOR�@�M��k0SMT��G��GR��3�a�PA�@��5�'�H� � j�A�T�OCjA7pP]Pp$OPd�O��C�%��p�O!��RE.pR�C�AO�?��Be5pR�EruIx'Q�G�e$PWR) IMdu�RR_$s��5�.�B Iz2H8�=��_ADDRH�H_LENG�B�q�q:��x�R��So�J.�SS��SK������ ��-�SE*���rmSN�MN1K	��j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ���p�Q� ��OUPW3��b_>�I��!q�a1 ��������|��� �����-���:���i+IOX2S=�D�e�x�]���L $��<p�!_OFF[r_��PRM_��bT�TP_�H��M (�pOBJ�"�pG�[$H�LE�C��>ٰN � 9�*��AB_�T��
�S��`�S��LV��KR�W"duHITCOU�?BGi�LO�q ����d� Fpk�GpsSS� ���HWh��wA��O.��`IN�CPUX2VISIO��!��¢.�á<��á-� �IOLN.)�P 87�R'�[p�$SL�bd P7UT_��$dp��Pz �� F_AuS2Q/�$LD���D�aQT U�0]P�Aa������PHYG�0��Z���5�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp����x��ٶ��-@J���S����NE�WJsOG�G �DIS��b&�KĠ��3T |���AV��`_�CTR<!S^�FLAGf2&�;LG�dU �n�:���3LG_SIZ���ň��=���FD��I����Z �ǳ� �0�Ʋ�@s��-ֈ�-ր=�-���-��0-�ISGCH_��Dq��N?�*��V��EE!2��C��n�U�����`LܞӔ�DAU��EA`��Ġt����GHr��I�BOO)�WgL ?`�� ITV���0\�REC�S#CRf 0�a�D^�����MARG��`!P�@)�T�/ty�?I�S��H�WW�I���T�JG=M��MNCH��I�_FNKEY��K��7PRG��UF��Pn��FWD��HL�STP��V��@��,���RSS�H�` �Q�C�T1�ZbT�R ����U�����|R��t�di���G��8PPO���6�F�1�M��FOC�U��RGEXP�TKUI��IЈ�c ��n��n����ePf� ��!p6�eP7�N���C�ANAI�jB��VA�IL��CLt!;eDCS_HI�4�.�"�O�|!�S �Sn�e��_BWUFF1XY��PT�$�� �v���f��� �A�rYY���P �����pOS1
�2�3���� >0Z �  ��apiE�*��IDX�d	P�RhrO�+��A&+ST��R��Yz�<!� Y$EK&C K+���Z&m&�5�0[ L��o�0�� ]PL�6pwq�t^����w���7�_ \ ��`��瀰�7��#�0C��] ��CLD�P��;eTRQLI��jd.�094FLG z�0r1R3�DM�R7Ɩ�LDR5<4R5ORG.���e2(`���V�8�.��T<�4�d^ ��q�<4��-4R5S�`T�00m��0DFRCLMC!D�?�?3I@��&�MIC��d_� d���RQm��q�DSTB	�  ��Fg�HAX;b ��H�LEXCESHZr�rBMup�a`렁�B;d��rB`��`a��F_A�J��$[�O�H0K�db \���ӂS�$MB��L�IБ}SREQUI�R�R>q�\Á�XDESBU���AL� MPŁc�ba��P؃ӂ!BF�AND���`�`d�Ҙ��c�cDC1��I�N�����`@�(h?Npz�@q��o�_N�SwPST8� e�r7LOC�RI�p�EX�fA�p��A�A�ODAQP�f Xf��ON��[rMF�� ���f)�"I��%�e���T��FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y��RFЭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?
�uD�)�b�	@Ð�i �@CU��V��T0�eRR2�j� Dɐ�Qނ�Bd$OCALI�@F�G�:s�2�RIN��v��<��NTE���k�E���,��b����_Nl��ڂ��~�ՆR�m�DIV�DH��@ـn�$V؀�'c!$��$AZ�����~�[���oH �$B�ELTb��!ACC�EL+��ҡ��ICRC�t����T/!���$PS�@#2LPq�Ɣ83������<� ��PATH����D����3̒Vp�A_� Q�.�4�B�Cᐈ��_MGh�$DDxQ���G�$FWh���p��m�����b�DE���PPABNԗR?OTSPEED����00J�Я8��@��~P$USE_�2�P��s�SY��c�ZA kqYNu@Ag���OFF�q�MO�UN�NGg�K�OL�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I(���4�\B�ݠVEO�w�Ͳ23�_UPE�߳LOWL���00����D���Bp��� �1RyCʀƶMOSIV��JRMO���@GPE�RCH  �OV ��^��i�<!�ZD <!�c��d@�P��!V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�(��<�1Ӣ`0 ��RTI$Qx�0 MO���МB@ R�0J��D��s�H�x���b�DUM2(��S_BCKLSH_C(���>�=�q�#��U��ԑ���2�t�$ACLALvŲ�1n�PN�CHK00'%SD�RTY4�k��y�1r�q_6#2�_UM$Prj�Cw�_�SCL���ƠLMT_J1_�LO��@���q��E������๕�幘S�PC��7������P	Co���H� �PU�m�C/@�"XT_�c�C�N_��N��e���S	Fu���V�&#�����9�(���=�C�u�SH6#��c����1�Ѩ��o�0�͑
��_�PALt�h�_Ps�W�_10���4�R�01D�VG�Jb� L�@J�OGW����TORQU��ON*�Mٙ�sRHљ�&�_W��-�_=��PC��I��I�I�%II�F�`�JLA.,�1[�VC��0�D�B�O1U�@i�B\J�RKU��	@DBOL_SMd�BM%`�_DLC�BGRV���C��I��H_p� �*COS+\�(LN�7+X>$ C�9)I�9)u*c,)b�Z2 HƺMY@!̳( "TH&-�)TH�ET0�NK23�I��"=�A CB6CB=�C�A�B(261C�616SBC�T25'GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t���B�6���AQ|r�f$NE�DpIB U�\B$5��$!��!A�%Ep(G%(!LPH$U�2׵�2SXpCc%pC�r%�2�&�C�J�&!�V�AHV6H3�YLVhJV�uKV�KV�KV�KV
�KV�IHAHZF`RXM���wXuKH�KH�KH��KH�KH�IO2LORAHO�YWNOhJOuKUO�KO�KO�KO�KO�&F�2#1ic%�d�4GSPBALANgCE_�!�cLEk0H_�%SP��T&�b�c&�br&PFULC��hr�grr%Ċ1k�y�UTO_?�jTg1T2Cy��2N&� v�ϰctw�g�p�0Ӓ~���T��O���� �INSEGv�!�R�EV�v!���DIF���1l�w�1m�
�OB�q
����M�Iϰ1��LCHW3AR����AB&u�?$MECH,1� X:�@�U�AX:�P��pY�G$�8pn 
Z���|���ROBR�C�R��N�c��MS�K_�`f�p P Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�MTCOM_C@>j�q  L��p~��$NORE³�5���$�r 8f� GR�E�SD�0�ABF�$XYZ�_DA5A���DE�BU�qI��Q�s ��`$�COD��� ��k�F�f��$BUFINDXrР����MOR��/t $-�U��)��r�B��������G�ؒu � $SIMULT ��~��< ���OBJE�` ��ADJUS>�1�A'Y_Ik��D_�����C�_FIF�=�T� ��Ұ��{��p@� �����p�@��D��FRI��ӥT��RIO� ��E������OPWO�ŀv}0��SYSBU�@ʐ$SOP�����#�U"��pPRUN,�I�PA�DH�D�\���_OU�=���qn�$}�IMA�G��ˀ�0P�qIM����IN�q���?RGOVRDȡ:����|�P~���Р�0L�_6p���i��RB����0��M���E�DѐF� ��N`Md*�����̰SL�`�ŀw x $OwVSL�vSDI��DEXm�g�e�9w�$����V� ~�N���@w����Ûǖȳ�M�����q<��� �x HˁE�F�AT+US���C�0à�ǒ��BTM����I
f���4����(�ŀy DˀEz�g���PE�r�����
���EXE��V��E�Y�8$Ժ ŀz @ˁ��3UP{�h�$�p��XN���9�H�� �PG"�{ h? $SUB��c��@_��01\�MPW�AI��P����LO��<�F�p�$R�CVFAIL_C�f�BWD"�F����DEFSPup | Lˀ`�D�� U�UNI��S�b��R`���_L�pAP��̐���ā}���� B�~���|��`ҲNN�`KET��y���P� $�~���0SIZE�ଠ{����S<�OR��FORMAT/p � F��ᖫrEMR��y�U�X��³&�P�LI7�ā  �$�P_SWIp�����_PL7�?AL_ �ސR�A��B�(0C��Dnf�$Eh�����C_=�U� �� � ���~�J�3�0����TIA4���5��6��MOM������� �B�AD��*��* PU70NRW���W ��U����� A$PI�6���	 ��)�4l�}6�9��Q���c�SPEED�PGq�7�D� >D����>tMpt[��SAM�`�痰>��MOV ���$��p�5��5�D�1�$2��������{�Hip�IN?,{�F(b+=$��H*�(_$�+�+GAM�M�f�1{�$GE�T��ĐH�D����
�^pLIBR�ѝI.��$HI��_��Ȑ$*B6E��*8A$>G086LW=e6\<G9�6�86��R��ٰV��$PDCK�DQ�H�_����;" ��z�.%�7�4*�9�� �$IM_SRO�D�s"���LH�"�LE�O�0�\H��6@�� �ŀ��P�qUR_SC�R�ӚAZ��S_SAVE_D�E��NO��CgA�Ҷ��@ �$����I��	�I�  %Z[� ��RX" �� m���"�q�'"� 8�Hӱt�W�UpS(��рM��O㵐 .'}q��Cg���@ʣȳ��тM�AÂ� ?� $PY��g$WH`'�NGp� ��H`��Fb��Fb��Fb��PLM���	� 0h�H�{�X��O��z�Zp�eT�M���� pS��C��O__0_�B_�a��_%�� | S����@	�v��v  �@���w�v��EM��%� =�es�B�ːt��ftP��PM���QU� �U�Q���Af�QTH=�H{OL��QHYS�3ES�,�UE��B���O#��  -�P�0�|�gAQ���ʠu���O��ŀ�ɂv�-�8�A;ӝROG��a2D�E�Âv�_�Ā^Z�INFO&��+�h���bȜ�OI��� ((@SLEQ /�#������o���S`c0O�0�051EZ0NUe�_��AUT�Ab�COPAY��Ѓ�{��@M���N�����1�P�
� ���RGI�����X_�Pl�$�����`
�W��P��j@�G����EXT_CY�Ctb���p�����h�_NA�!�$�\�<�RO�`]��� � m��P�OR�ㅣ���SReVt�)����DI �T_l���Ѥ{�ۧ�Шۧ �ۧ5٩6٩7�٩8����S�B쐒���$�F6���PL�A�A^�TAR ��@E `�Z������<��d� ,(@FL�q`h��@YNL���Mz�C���PWR���쐔e�DELA4Ѱ�Y�pAD#qX� �QSKIP��� ĕ�x�O�`NeT!� ��P_x� ��ǚ@�b�p1�1� 1Ǹ�?� �?��>�@�>�&�>�3�>�9��J2R;쐖 m4��EX� TQ�� ��ށ�Q���[�KF�ܴ�w�RDCIf� )�U`�X}�R�#%�M!*�0�)��$RGE7AR_0IO�TJB�FLG�igpER�a��TC݃������2�TH2N��� S1�b��Gq T�0' ����M���`�Ib���R�REF:�1�� l�h���ENAB��lcTPE?@���!(ᭀ�� ��Q�#�~�+2 H�W���2�Қ���"�P4�F�X�j�3�қ{�@��������j�4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:Lj�7�ҟo@�����j�8�ҁ���"4F ���SMSK��R���a��E�A���REMOTE������@ "1��Q��IO�5"%I��P���POWi@쐣  �����X�gpi������Y"$DSB_SIGN4A�Qi�̰�C�ШP�S232�%�Sb�iDEVI�CEUS#�R�RP�ARIT�!OP�BIT�Q��OWCONTR��Q�Ѭ��RCU� M�SU_XTASK�3NB���0�$TATU�P#�"@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�UKPDl�ARB�#P%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG�G|�.2���F��1�!d�9Z�8+5K��+5��E�y�L0�4��X �0m�LN�T�3Hz��89��%�4�3%G��W�0�W�RdD�Z��Tܳ��K�a�3d��$cV 2!���1��I1H�0U2K2sk3K3J ci�aI�i�a�L��SLL��R$Vؠ�BV�E�Vk��A bQ*R��� �,6Lc���9V2�F{/P:B��PS_�E���$rr�C�ѳ3$A0��wPR���v�U�cSk�� {��8��G� 0���VX`�!�tX`��0P�Ё��
�Љ2SK!� E�-qR��!0����z�NJ AX�!h�A�@LlA��A�THI�C�1�������1T�FE���q>�IF_CH�3A�I0�����G1�x������9º��Ɇ_JF҇P�R(���RVAT�� �-p��7@̦���DO�E��CO9U(��AXIg���OFFSE+�TRIG�SK��c���Ѽe�[�K�Hk���8�IGGMAo0�A-������ORG_UNE9V��� �S��?�d �$����=��GROU��ݓ�TO2��!ݓDSP���JOG'��#	�_	P'�2OR���>Pn6KEPl�IR�d0�PM�RQ�AP�Q²�E�0q�e���SY�SG��"��PG��B�RK*Rd�r�3�-�`������ߒ<pAD��<ݓJ�BSOC� �N�DUMMY1�4�p\@SV�PDE�_OP3SFSP_D_OVR��ٰ1CO��"�OR-���N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA�"�LCHDL�REGCOV��0�W�@1M�յ�RO3�r�_�0� @���@VERE�$O�FS�@CV� 0BWDG�ѴC��2j�
��TR�!��E_�FDOj�MB_CiM��U�B �BL=r0�w�=q�tVfQ��x0�sp��_�Gxǋ�AM���k�J0������_M���2{�#�8$C�A�{Й���8$HcBK|1c��IO��q.�:!aPPA"ڀN�3�^�F���:"�DVC_DB�C��d� w"����!��1������3����ATIO"� �q0�UC�&CAB�BS�P ⳍP�Ȗ��_0c�?SUBCPUq��S�Pa aá�}0�Sb���c��r"ơ$HW�_C��� :c��IcA��A-�l$UNIT��l��ATN�f�����CYCLųNE�CA��[�FLTR_2_FI���(�ӌ}&��LP&�����_�SCT@SF_��F0����G���FS|!����CHAA/����2��RSD�x"ѡ�b�r�: _T��PR�O��O�� EM�_���8u�q �u�q��DI�0e�R�AILAC��}RM�ƐLOԠdC��:a`nq��wq����PR��%SLQ�pfC�ѷ =	��FUNCŢ�rRINkP+a�0 �f�!RA� >R 
�p��ԯWARF�BLFQ��A�����DA�����LDm0�aBd9��nqBTIvrpbؑ���PRIAQ1�"AFS�P�!���@��`%b���M�9I1U�DF_j@��ly1°LME�FA�@OHRDY�4��Pn@�RS@Q�0"�MU�LSEj@f�b�qG �X��ȑ����$.A$�1$�c1Ó���� x~�EG�0ݓ��q!AR����09p>B�%��AXE���ROB��W�A4�_�-֣SY���!6��&MS�'WR���-1���STR��5�9�E�� 	5B��=QB90�@6������kOT�0o 	$�ARY8�w20����	%�FI��;�$�LINK�H��1��a_63�5�q�2XYZ"��;�q�3�@��1�2�8{0B�{D��� CFI��6G��
�{�_J��6��3a'OP_O4Y;5�Q#TBmA"�BC
�z��DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ ��@�5<:7�� +1�?0K�Mc�6�8Cb�vrb�4�ORQ��X�>8�#op�� ����wq�Uf�����T'OVE�Q��M;�@E#�UK#�UQ"�VW�Z Q�W���Tυ� ;� ���QH�!`�ҽ��U�Q��WkeK#kecXER��	GE	0��S�dAWaǢ:D���7!�!AX�rB! {q��1uy-!y �pz�@z�@z6Pz \Pz� z1v�y �y�+y�;y�Ky �[y�ky�{y��y��q�yDEBU��$����L�!º2WG`  AB!�,��S9V���� 
w��� m���w����1���1�� �A���A��6Q��\Q����!�m@��2CLAB3B�U�����S{ R �SER��>�� � $�@� mAؑ!p�PO���Z�q0w�^�_MR}Aȑ� d  9T�ĴERR��TYz�B�I�V83@�cΑTOQ�d:`!L� �d2�]�X�}C[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	V FZN_wCFG_!� 4�� ?º�|�ų����@�Ȳ�W �]���\$� �n���Ѵ��9c�Q��(�FA�He�,�XEDM�(�����!�s�Q�g�P{RV H�ELLĥ� }56�B_BAS!�GRSR��ԣo �#QS��[��1r�%��U2ݺ3ݺ4ݺ5ݺ�6ݺ7ݺ8ݷ��R�OOI䰝0�0NL�K!�CAB� ��A[CK��IN��T:��1�@�@ z�m�_P�U!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KcARӑ��RE~���P��(��QUE������P
��CST?OPI_AL������0&���㰑�0SE�Ml�b�|�M��d�T�Y|�SOK�}�DI������(���_T}M\�MANRQ���0E+�|�$KEYSWITCH&�	���HE
�BE�AT����E� LE(Ғ���U��FO���|��O_HOM��O�REF�PPR�z��!&0��C+�OA�ECO��B�rIOCM�D8׵��\���8�` � DH�1����U��&�MHx�»P�CFORC��n� ��OM�  � @V��|�U,3P� 1-�`� �3-�4�p �SN�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��0�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fi�7s��VP�U�PD��  ���|�԰��YSLO>Ǣ� � z��� ����o�E��`>�^t���АALUץ����C�U���wFOqID_YL�ӿuHI�zI�?$FILE_���tf��$`�JvSA���� h���E_B�LCK�#�C,�D_CPU<�{�<�o�����tJr��R ;��
PW O�[ ��LA��S��8������RUNF�Ɂ ��Ɂ����F�ꁡ�ꁾ�� �TBCu�C�� �X -$�LENi��v������I��G�LOWo_AXI�F1�
�t2X�M����D�
 ���I�� ��}�T#OR����Dh��� L=��⇒�s���#�_MA`�ޕ���ޑTCV����T ���&��ݡ����J�$����J����Mo����J�Ǜ �������2�Ѓ v�����F�JK��VKi�ΡvњΡ3��J0�ңJ�JڣJJ�AAL�ң�ڣ��4�5z�&�N1-�9����ʅ�L~�_Vj��&y���� ` ��GROU�pD��B>�NFLIC��REQUIREa�EBUA��p����2¯�����c��� \��APP�R��C���
�E�N�CLOe��SC_M v�,ɣ�
�ޣ�� ���MCp�&���g�_MG�q�C� �{�9���|�wBRKz�NOL��t|ĉ R��_LI|�H�Ǫ�k�J����P
� ��ڣ�����&���/����6��6��8��������� ���8�%�W�2�e�PATHa�z�p�z�=�hvӥ�ϰ�x�CN=��CA�����p�INF�UC��bq��CO�UM��YZ������q�E%���2������P�AYLOA��J2=L3pR_AN��<�L��F�B�6�R�{�R_F2LSHR��|�LOG��р��ӎ�>��ACRL_u��Ր����.���H�p��$H{���FLEX�
�s�J�� :�/����6�2�`����;�M�_�F16� ����n���������ȟ��Eҟ�����,� >�P�b���d�{�������������5�T��X��v���E ťmFѯ����� ��&�/�A�S�e�D�}Jx�� � ��0����j�4pAT����6n�EL  �%ø�J���ʰJE��C�TR�Ѭ�TN��F�&��HAND_V�B[
�pK�� $F2{�6� �r�SW$#�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�(#�� &0�_�ERx!V9�SQASYM��] �����x��ݑ���_SHl������̀sT�(����(�:�J�A���S�cir��_�VI�#Oh9�``V_UNI��td�~�J���b�E�b��d�� �d�f��n���������$uN����D�찙H������"CqE�N� a�DI��>�Opbt2Dpx�� �
�2IxQA����q���-��s �� �����{ ��OMME���rr/�TVpP�T�P ���qe�i� ���P�x ��yT�Pj�� $DUMM�Y9�$PS_f��RFq�0$:�� ���!~q�c X����K�STs��ʰSBR��M2�1_Vt�8$SV_ERt�O��z���WCLRx�A  O�r�?p? Oր � �D $GLOB���#LO��Յ$�po��P�!SYS�ADR�!?p�pTC}HM0 � ,�����W_NA���/�e�$%SR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T>D�XSCRE�ƀ5�� ��STF���#}�pТ6�1] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��t<qUE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SSx�!&; SHIF��|s�P�p�6�s����R���OSURzW�pRADIz��2�_�q�h�g! ؎q)�LUza$�OUTPUT_BM��IML�oR6�(`)�@TIL<SCO�@Ce�;�� 9��F��T��a�� o�>�3�����w�E2u�ӝ�P{t���%�DJU��|#�/WAIT����ک�%ONE��Y�BOư ��� $@p%�C�SB�n)TPE��NEC���x"�$t$���*B_T��R��%�qR� $���sB�%�tM�+Z��t�.�F�R!݀��O�Pm�MAS�_DUOG�OaT	�D�����C3S�	�O2DELcAY���e2JO�� n8E��Ss4'#J�aP60%�����Y_��O2�� �2���5��`?� ;��ZABC~S��  $�2��J�
���$$C�LAS����i�A���� @�VIRT��O.@A�BS�$�1 <E�� < *AtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v���8��M@[�AXLր��&A�dC  ���IqN��ā��PRE������LAR�MRECOV �<I䂥�NG�� �\K	 A  � J�\�M@PPLIMC�?<E�E��Handl�ingTool ��� 
V7.5�0P/28[�  o��o��
�w_SW�� UP*A7� ��F0ڑ���AG@�� S20��*A���:�ާ�X{FB �7DA5�� �'@�oy@����None������� ��T��*A4yn+xl�_��V����:g�UTOB���������HGAPO�N8@��LA��U��D� 1<EfA����������� Q 1שI Ԁ��Ԑ�:�i�n��܍�#BGB �3��\�HE�Z��r�HTTHKY ��$BI�[�m����� 	�c�-�?�Q�o�uχ� �ϫϽ��������_� )�;�M�k�q߃ߕߧ� ���������[�%�7� I�g�m������� ������W�!�3�E�c� i�{������������� ��S/A_ew �������O +=[as�� �����K//'/ 9/W/]/o/�/�/�/�/ �/�/�/G??#?5?S? Y?k?}?�?�?�?�?�? �?COOO1OOOUOgO yO�O�O�O�O�O�O?_�	__-_K_Q_��(�T�O4�s���DO_C�LEAN��e��SN�M  9� ��9oKo]ooo�o�D?SPDRYR�_%�HI��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ|��g�PLUGGҠ��Wߣ��PRC�`B�`9��o�=�OxB��oe�SEGF��K������o%o�����#�5�m���LAP �oݎ����������џ �����+�=�O�a�>��TOTAL�.����USENUʀ�׫ �X���R(�RG�_STRING �1��
��M��Sc�
��_�ITEM1 �  nc��.�@�R�d�v� ��������п������*�<�N�`�r��I/O SIGN�AL��Try�out Mode��Inp��Simulated��Out��O�VERR�` = �100�In �cycl���P�rog Abor������Stat�us�	Hear�tbeat��M?H FaulB�K�AlerUم�s߅� �ߩ߻��������� �S���Q�� f�x���������� ����,�>�P�b�t�p������,�WOR�� ����V��
.@ Rdv����� ��*<N`PO��6ц��o �����//'/ 9/K/]/o/�/�/�/�/��/�/�/�/�DEV �*0�?Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�OPALTB��A�� �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_�oo(o:o�OGRI �p��ra�OLo�o�o�o �o�o�o*<N `r������`o��RB���o�>� P�b�t���������Ώ �����(�:�L�^�xp����PREG�N ��.��������*� <�N�`�r����������̯ޯ���&�����$ARG_��D �?	���i���  w	$��	[}��]}���Ǟ�\�SB�N_CONFIG� i��������CII_SAV/E  ��۱Ҳ�\�TCELLSE�TUP i�%�HOME_IO��͈�%MOV_8�2�8�REP����V�UTOBACK�
�ƽF�RA:\�� X�Ϩ���'`!���x������ �� ��$�6�c�Z�lߙ���������������� �!凞��M�_�q�� ���2��������� %�7���[�m������ ��@�������!3E$���Jo��p�����INI�@���ε��MESSAG����q�>�ODE_D$��ĳ�O,0.��PA�US�!�i� ((Ol���� ���� /�// $/Z/H/~/l/�/�'a~kTSK  qx�����UPDT%��d0;WSM�_CF°i��еU�'1GRP 2�h�93 |�B��A|�/S�XSCRD+1;1
1; ����/�?�?�? OO$O ��߳?lO~O�O�O�O �O1O�OUO_ _2_D_�V_h_�O	_X���GR�OUN0O�SUP�_NAL�h�	ܢĠV_ED� 1�1;
 �%-B?CKEDT-�_`�!oEo%���a�o�����ߨ���e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[8�5GED4�n�#�� ~�j���ED5Z��Ǐ6� ~��8�}���ED6�����k�ڏ ~G���!�3�ED7��Z��~� ~�8V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W�Ư�
}3�����CR o�����3�տ@ϯ�����P�PNO_DE�L�_�RGE_UN�USE�_�TLAL_OUT q��c�QWD_ABO�R� �΢Q��ITR�_RTN����N'ONSe����CAM_PARA�M 1�U3
 �8
SONY �XC-56 234567890�H� � @����?���( Щ�V�|[r؀~�X�HR5k�|U�Q��ο�R57����A�ff��KOWA SC310M|[�r�̀�d @6�|V��_�Xϸ� ��V��� ���$�6���Z�l��CE_RIWA_I857ЍF�1��R|].��_LIO4W=� ���P<~�F<�GwP 1�,����_GYk*C*�  ��C1� 9J� @� G� �CL�C]� d� l� s��R� ��[�m�� v� � �� ��� C�� �"��|W��7�HEӰON�FI� ��<G_P_RI 1�+P� m®/���������'CHKPAU�S�  1E� ,�>/P/:/t/^/�/ �/�/�/�/�/�/?(?@?L?6?\?�?"O������H�1_MO�R�� �XaB�iq-���5 	 �9 O�?$OOHOZK��2	���=9"�Q?$55��C�PK�D3�P������aÃ-4�O__|Z
 �OG_�7�PO�� ��6_���,xV�ADB����='�)
mc:c?pmidbg�_`ϖ�S:�)����Yp0�_)o�S`�BBia�P�_mo8j�)�aKoo�o9i�)Ѕ�og�o�o�oLnf��oGq:I�ZDEFg f8��)�R�6pbuf.txt m�]n�@����# �	`)Ж�A=L�m��zMC�21�=���9���4�=��n׾�Cz  BH�BCCPUeB��_B�y;���>C���Cn�SZE@E?{hD�]^Dْ?�r����D��^���G	��F���F��Cm	�fF�O�F��I�SY���vqG����Em�)�.����1)��<�q�G�x�2��Ң �� a�D��j���E�e��X��EQ�EJP� F�E�F�� G���F^�F E�� FB�� H,- Ge���H3Y����  >�33 s���xV  n2xQ@��5Y��8B� yA�AST<#�
�� �_'�%��wRS/MOFS���~2��yT1�0DE ��O c
�(�;��"�  <�6�z�Rb���?�j�C4�)�SZm� W��{�Jm�C��B-G�C�`�@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"��_ , 
�^����o xvf`MT�I�^�rl@�:sONT�IM�������Zv�i
õ�cMOT�NEND���dRECORD 1(R�qa��ua�O��q ��sb�.�@�R��x Z�������ɏۏ� ����#���G���k�}� ����<�ş4��X�� �1�C���g�֟���� ����ӯ�T�	�x�-� ��Q�c�u�������� ��>����)Ϙ�M� ��F�࿕ϧϹ���:� ������%�s`Pn&�]� o��ϓ�~ߌ���8�J� ����5� ��k��� �ߡ��J�����X�� |��C�U�������� ���0�����	��db�TOLERENC�qdBȺb`L����PCS_CFG �)�k)wdM�C:\O L%04�d.CSV
�`cl�)sA �CH� z�`)~���h�MRC_OUT �*�[�nSG�N +�e�r���#�10-MAY�-20 10:3�7*V15-JAN�j51�k P/Vt��)~�`�pa�m��P�JPѬVE�RSION �SV2.0.�8.|EFLOGI�C 1,�[ 	DX�P7)�PF."�PROG_ENB��o�rj ULSew ��T�"_WRST�JNEp�V�r`dEM�O_OPT_SL� ?	�es
 ?	R575)s7)��/??*?<?'�$TO  �-��?&[V_@pEX�Wd�u��3PATH ASA\�?�?O�/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C��SqqF�PMAU�� t/XrMSWR.D�i�a.|S/�Z!D_N�O0__T_C_�x_g_�_�tSBL_/FAUL"0�[3w/TDIAU 16M�a�p�A12�34567890gFP?BoTofo xo�o�o�o�o�o�o�o ,>Pb�S�p-P�_ ���_s �� 0`����� )�;�M�_�q����������ˏݏ��|)UM�P�!� �^�T�R�B�#+�=�PME�fEI�Y_TEMP9 È�3@�3A �v�UNI�.(YN_BRK 2Y�)EMGDI_S�TA�%WЕNC2_SCR 3��1o"�4�F�X�fv����������#��ޑ14����)�;���t��ݤ5��� ��x�f	u�ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /߭P�b�t�� ��x� �߰���������
�� .�@�R�d�v���� ����������*�<� N���r����������� ����&8J\ n������� �"`�FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/4?,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O? �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �o�O�O�o�o�o
 .@Rdv��� ������*�<� N�`�r����o����̏ ޏ����&�8�J�\� n���������ȟڟ�����H�ETMODoE 16���W ��ƨ
R��d�v�נRROR_PROG %A��%�:߽�  ��TABLE  A�������#�L�RR�SEV_NUM � ��Q���K�S���_AUTO_ENB  ���I�Ϥ_NOh� �7A�{�R�  �*������������^�+��Ŀֿ迄��HISO���I�}�_�ALM 18A�� �;�����+ �e�wωϛϭϿ��_H���  A��|��4�TCP_�VER !A�!�����$EXTLO�G_REQ��{�V�SIZ_�Q�T�OL  ��Dz���A Q�_B�WD����r���n�_�DI�� 9���}�z���m���ST�EP����4��OP�_DO���ѠF�ACTORY_T�UN�dG�EAT?URE :�����l�Han�dlingToo�l ��  - C�Englis�h Dictio�nary��ORD�EAA Vi�s�� Masteyr���96 H���nalog I/yO���H551���uto Soft�ware Upd_ate  ��J���matic Ba�ckup��Par�t&�ground Edit���  8\ap�Camera��F���t\j6R�elyl���LOADR�7omm��shq��oTI" ��co��
! o���p�ane�� 
!���tyle s�elect��H5�9��nD���oni7tor��48�����tr��Relia�b���adin�Diagnos�"����2�2 ual� Check S�afety UI�F lg\a��h�anced Ro�b Serv q� ct\��lUs�er FrU��D�IF��Ext. oDIO ��fiAs d��endr �Err L@��I%F�r��  �П��90��FCTN /MenuZ v'���74� TP In���fac  S�U (G=�p���k Excn g��3��High-wSper Ski+�  sO�H9 � m�munic!�on5sg�teur� �����V����c�onn��2��ENމ�Incrst�ru���5.fd�KAREL �Cmd. L?u�aA� O�Runw-Ti� Env��R��K� ��+%�s#�S/W��74��L?icenseT��  (Au* ogBook(Sy���m)��"
MACROs,V�/Offse��a�p��MH� ����p�fa5�MechS�top ProtL��� d�b i��Shif���j545�!xr ��#���,�}b ode Switch��m\e�!o4.�& pro�4���g��Multi�-T7G��net�.Pos RGegi��z�P���t Fun���3s Rz1��Numx ������9m�1�  �Adjuj��1 J7�7�* ����6�tatuq1EIK�RDMtot���scove�� ���@By- }uest1�$Go� � U5�\SNPX �b"���YA�"Li�br����#�� �$~@h�pd]0�J�ts in VCCCM�����0�  �u!��2 R�0�/�I�08��TMI�LIB�M J92:�@P�Acc>�F�{97�TPTX�+6�BRSQelZ0�M�8 Rm��q%��6�92��Unexc�eptr motn>T  CVV�P���KC����+-��~K  II)�VS�P CSXC�&.ac�� e�"�� t�@�Wew�AD� Q�8bvr nm�en�@�iP� a�0y�0�pfGri�dAplay !�� nh�@*�3R�1M-�10iA(B20k1 �`2V"  F����scii�lo{ad��83 M��yl����Guar�dO J85�0�mP'��L`���stuaPa9t�&]$Cyc����|0ori_ x%Da�ta'Pqu���cAh�1��g`� j� RLJam�5���IMI De-B(�\A�cP" #^0C~  etkc^0�asswo%q�)6�50�ApU�Xn�t��Pven�CT�qH�5�0YELLOW BO?Y���� Arc�0vi�s��Ch�Wel=dQcial4Izt�Op� ��gs�`k 2@�a��poG3 yRjT1 NEf�#HT� xyWbF��! �p�`gd`����p\� =P��JP�N ARCP*P�R�A�� OL��pSup̂fil��p��J�� ��cro�670�1C~E�d���SS�pe�tex��$ �P� So7 t^� ssagN5 <Q"�BP:� �9 "0�Q#rtQC��P�l0dpn�笔�rpf�q��e�ppmas�cbin4psy=n�' ptx]08��HELNCL �VIS PKGS9 �Z@MB &���B J8@IPE� GET_VAR� FI?S (Un�i� LU�OOL:� ADD�@29.KFD�TCm���E�@�DVp���`A�ТN�O WTWTEST �� ��!��c��FOR ��ECT� �a!� ALSE� ALA`�CPMO-130��� b �D: HANG FROMg��2���R709 DRA�M AVAILC�HECKS 54�9��m�VPCS �SU֐LIMCH�K��P�0x�FF WPOS� F�� q�8-12 C�HARS�ER6�O�GRA ��Z@AV�EH�AME��.SV��Вאn$��9�wm "y�TRCv�� SHADP�UP�DAT k�0��S�TATI��� M�UCH ���TI�MQ MOTN-�003��@OB�OGUIDE DAUGH���b��@�$tou� �@C� <�0��PATH�_��MOVET�� R�64��VMXPA�CK MAY A�SSERTjS��C�YCL`�TA��B�E COR 71��1-�AN��RC �OPTIONS � �`��APSH-�1�`fix��2�S�O��B��XO򝡞�_�T��	�i��0j��d�u�byz p wa��y�٠HI�������U�pb XSPD �TB/�F� \hcehΤB0���END�[CE�06\Q�p{ }smay n@��pk��L ��tr'aff#�	� ���~1from sy�svar scr��0R� ��d�DJUD���H�!A��/��SET ERR��D�P7����NDA�NT SCREE�N UNREA �VM �PD�D��P�A���R�IO gJNN�0�FI��}B��GROUNנD Y�Т٠�h�SVIP 53 Q�S��DIGIT �VERS��ká�N{EW�� P06�@=C�1IMAG�ͱ4���8� DI`����pSSUE�5��EPLAN JON�� DEL���157�QאD��CALL�I���Q��m���IP�ND}�IMG N�9 PZ�19��MwNT/��ES ���`LocR Hol�߀=��2�Pn� PG�:��=�M��can�����С: 3D� mE2view gd X��ea1 ��0b�pof Ǡ"�HCɰ�ANNO�T ACCESS? M cpie$E�t.Qs a� lo^MdFlex)a:���w$qmo G�sA�9�-'p~0��h0pa���eJ AUTO1-�0��!ipu@Т|<ᡠIABLE+�� 7�a FPLN:9 L�pl m� �MD<�VI�и�W�IT HOC�Jo~1Qui��"���N��USB�@�Pt� & remov����D�vAxis �FT_7�PGɰC�P:�OS-14�4 � h s 2968QՐOST�p � CRASH D�U��$P��WOR�D.$�LOGI�N�P��P:	�0�0�46 issue�E�H�: Slo[w st�c�`�6����໰IF�I�MPR��SPOT�:Wh4���N1STyY��0VMGR�\b�N�CAT��4oR�RE�� � 5�8�1��:%�RTU�!Pe -M a�SE:B�@pp���AGpL��r�m@all���*0a�OCB WA����"3 CNT0� T9DWroO0a�larm�ˀm0d� t�M�"0�2|� 9o�Z@OME<�� ���E%  #1-�S�RE��M�st}0g�     5K�ANJI5no �MNS@�INISITALIZ'�3 E�f�we��6@�� dr�@ fp �"��SCII L��afails w|��SYSTE[��i��  � Mq��1QGro8�m �n�@vA����&��nx�0q��RWRI �OF Lk��� \gref"�
�up� de-rela�Q_d 03.�0SS�chőbetwe�4�IND ex 6ɰTPa�DO� �l� �ɰGigE��soperabi]l`p l,��Hc�B��@]�le�Q0c�flxz�Ð���O�S {����v4pfigi GLA�$�c2z�7H� lap�0�ASB� If��g�2 l\c�0��/�E�� EXCE	 㰁�P���i��� o0��Gd`]Ц�f<q�l lxt��EFal��#0�i�O�Y�n�CLOS��S[RNq1NT^�F��U��FqKP�ANIO' V7/ॠ1�{����DB �0���v��ED��DET|��'� �bF�NLI;NEb�BUG�T�:��C"RLIB��A���ABC JAR�KY@��� rkeMy�`IL���PR���N��ITGAR� D$�R �Er *�T��a�U�0��h�[��ZE V� TASK p.vr��P2" .�XfJ�srqn�S谥dIBP	c����B/��BUS.��UNN� j0-��{��cR'���LO�E�DIVS�CUL`s$cb����BW!���R~�W`P�����I�T(঱tʠ�OF��UNEXڠ+����p�FtE��SVE�MG3`NML 5�05� D*�CC_SAFE�P*� ���� PET��'P�`��F  !���IR(����c i S>� �K��K�H GU�NCHG��S�M�ECH��M��T�*�%p6u��tPOR�Y LEAK�J���SPEgD��2�V 74\GRI���Q�g��CTLN��TRe @�_�p ��6�EN'�IN���`���$���r��T3)�.i�STO�A�s�	L��͐X	���q��1Y� ��TO2�J �m��0F<�K����D)U�S��O��3	 9�J F�&���S?SVGN-1#I�N��RSRwQDAU�C@ޱ� �T6�g��� 3��]���BRKCTR8/"� �q\j5��_��Q�S�qINVJ0D ZO�Pݲ���s���г�Ui ɰ̒�a�D�UAL� J50�e�x�RVO117 AW�TH!Hr%�nN�247%�52��|�&aol ���R��(�at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���M�d�Rǰt� \fosB�A�0Np�c�����{�U��ROP �2�b�pB��ITP�4M��b !AU�t c0< � plet9e�N@� z1^q�R635 (Ac�cuCal2kA���I) "�ǰ�1
a\�Ps��ǐ� b���0P򶲊���ig�\cbacul "A3p_ �1��ն����etaca��AT���PC�`�����;_p�.pc!Ɗ�<�:�circB����5�tl��Bɵ�:�f!m+�Ί�V�b�ɦ�~r�upfrm.����ⴊ�xed��Ί�N~�pedA�D �}b>�ptlibB�� �_�rt��	Ċ�a_\׊ۊ�6�fm�� ��oޢ�e��̆Ϙ���c�Ӳ�5�j>�����#tcȐ��	�r���ʸ�mm 1��T�sl�^0��T�mѡ�#�r�m3��ub Y�q�s3td}��pl;�&�cckv�=�r�vf������9�vi����Cul�`�0fp�q ��.f��� daq�; i Data A�cquisi��nB�
��T`��1��89��22 D�MCM RRS2�Z�75��9 3 �R710�o59�p5\?��T "��1 (D�T� nk@��������E Ƒ�ȵ��Ӹ�etdm�m ��ER����gxE��1�q\mo? ۳�=(G���[0(

�2�` ! �@�JMACRO��S�kip/Offs�e:�a��V�4o9<� &qR662����s�H�
 6Bq8�����9Z�43 �J77� 6�J783�o ��n�"vv�R5IKCBq?2 PTLC�Z�g R�3 (�s�, �������0�3�	зJԷ\sf�mnmc "MN�MC����ҹ�%mnf�FMC"Ѻ0�>� etmcr� ��8���� ,��}D�} �  874\p'rdq>,jF0�ޢ�axisHPr�ocess Axwes e�rol^�PRA
�Dp� 56o J81j�59� 56o6� ���0w��690 98� [!I#DV�1��2(x2��2ont�0�
�����m2���?C��e�tis "ISD���9�� Fprax�RAM�P� D��d�efB�,�G�is_basicHB�@p޲{6�� 708�6��(�Acw:�������D
�/,��AMOX �� ��DvE��?;T��2>Pi� RAFM';�]�!PAM�V�W�Ee`�U�Q'
bU�75��.�ceNe� nt?erface^�1' 5&!54�K��b(Devam±�/�#����/<�Tane`"�DNEWE���btp_dnui �AI�_�s2�d_rsono���bAsfjN��bdv_arFvf�x0hpz�}w��hkH9x�stc��gApon1lGzv{�ff� �r���z�3{q'�Td>pchamp�r;e�p� ^597@7��	܀�4}0��mɁ��/�����lf�!�pcochmp]aMP&xB�� �mpev��8����pcs��Ye�S�� Macro�OD��16Q!)*��:$�2U"_,��Y�(PC ��$_;�������o��J�gegemQ@GEMSW�~ZG�gesndy��OD��ndda��S��s1yT�Kɓ�su^Ҋ�ĩ�n�m���L��  ���9:p'ѳ޲���spotplusp���`-�W�l�J��s��t[�׷p�key�ɰ�$��s�-Ѩ��m���\featu� 0FEAWD�o;olo�srn'!�2 p���a�As3��t�T.� (N. A.)��!e!�J#
 (j�,��oBIB��oD -�.�n��k9�"K��u[-�_����p� "PSE�qW����wop "sEЅ�&�:�J��� ���y�|��O8��5� �Rɺ���ɰ[��X� ������%�(
ҭ�q HL�0k�
�z�@a!�B�Q�"(g� Q�����]�'�.��� ��&���<�!ҝ_�#��tpJ�H�~Z��j��� ��y������2��e� �����Z����V��! %���=�]�͂��^2�@�iRV� on�Q$Yq͋JF0� 8ހ�`�	(^�dQueue���X\1�ʖ`�+~F1tpvtsn��YN&��ftpJ0v �RDV�	f��J1 iQ���v�en�^�kvstk��mp���btkclrq8���get�����r��`kacqk�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�m	c�N+v3�_� �����.v�/\jF��� �`Q�΋�ܒ�N50 (FR�A��+��͢fraparm��Ҁ�} =6�J643p:V��ELSE
#�V�AR $SGSY�SCFG.$�`_UNITS 2�D`G~°@�4Jgfr��4A�@FRL-��0ͅ �3ې���L�0NE�: �=�?@�8�v�9~Q�x304��;�BPR�SM~QA�5TX.�$VNUM_OLp��5��DJ507��~l� Functʂ�"qwAP��琉�3 �H�ƞ�kP9jQ�Q5 ձ� ��@jLJzBJ[ �6N�kAP����S>��"TPPR��\�QA�prnaSV��ZS��AS8Dj510U�-�`cr�`8 ���ʇ�DJR`jYȑH_  �Q �P�J6�a21��48�AAVM 5̕Q�b0 lB�`TU�P xbJ54s5 `b�`616����0VCAM ~9�CLIO b71�5 ���`gMSC8�
rP R`�\sSTYL� MNIN�`J6�28Q  �`NR�Ed�;@�`SCH ���9pDCSU M�ete�`ORSR� Ԃ�a04 kR�EIOC �a5.�`542�b9vpP@<�nP�a�`�R�`7�`��MASK 3Ho�.r7 �2�`OOCO :��r3� �p�b�p���r0X��a��`13\mn�a3?9 HRM"�q�q~��LCHK�u�OPLG B��a0�3 �q.�pHCR� Ob�pCpPosyi�`fP6 is[r�J554�òpDS�W�bM�D�pqR�a337 }Rjr0 �1�s�4 �R6�7��52�r5 �2�r7 1� P6���Regi��@T�uFRD�M�uSaq%�4�`9{30�uSNBA�u�SHLB̀\sf�"pM�NPI�S�PVC�J520v��TC�`"MNрoTMIL�IFV��PAC W�pTP�TXp6.%�TELN N Me��09m3UEC9K�b�`UFR�`���VCOR��VIPuLpq89qSXC�S��`VVF�J�TPy �q��R626l��u S�`Gސ�2�IGUI�C��P�GSt�\ŀH86�3�S�q�����q34:sŁ684���a��@b>�3 :B��1� T��96 .�+�E�51 y�q53̀3�b1 ���b1 �n�jr9 ���`VAsT ߲�q75 s�xF��`�sAWSMӞ�`TOP u�ŀRq52p���a80 
��ށXY q���0 \,b�`885�QXр�OLp}�"pE࠱t�p�`LCMD��EgTSS���6 �>V�CPE oZ1�gVRCd3
�NLH�h��001m2Ep���3 f��p��4 //165C��6l����7PR��008 �tB��9 -200��`U0�pF�1޲1	 ��޲2L"���p���޲4��5 \h�mp޲6 RBCF`�`ళ�fs�8 ������~�J�7 rbcfA�L�8\PC����"�32m0u�n�K��Rٰn�5 5EW�
n�9 z��4�0 kB��3 ��6|ݲ�`00iB/��I6�u��7�u��8 �0�������sU0�`�t� �1 05\rb��2 E���K���dj���5˰��60��a�HУ`:�63�jAF�_���F�7 ڱ݀H�a8�eHЋ��cU0���7�p��1u��8<u��9 73����&��D7� ��5t�W97 ��8U�1���2��1�1:���h���1np�"��8(�U=1��\pyl��,�p��v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6C B���цp��1��r��1�`͵155ض�157 �2��62 �S����1b��2$����1Π"�2����B6`�1<c�4� 7B�5 DR��8�_�B/��187 �uJ�8 06�9s0 rBn�1 (���202 0EW,�ѱ2^��2��90�U12�p�2��2 b��u4��2�a"RB����9\�U2�`w�l����4 60Mp��7�������b�s
5 ¿�3����pB"9 �3 ����`ڰR,:7 �2��V�2���5���2^��a^9����qr����n�5 ����5᥁"�8a�Ɂ}�5B���5����`!UA���� ��86 �+6 S�0��5�p�2<�#�529 �2^��b1P�5~�2�`���&P5��8"��5��u�!�5��ٵW544��5��R��P nB^z�c (4�����U5J�V�5��1�1^���%�����5 b2a1��gA��58W[82� rb��5N��E�5890r� 1�95 �"������ c8"a��|�L ���!�J"5|6��^!�6��B�"8�`#��+�58%�6B�AME�"�1 iC��622D�Bu�6V��d� 4��{84�`ANRSP�e/S� C�5 � �6� ��� \� �6�� �V� 3t��� �T20CA�R��8�� Hf� 1DH�� A�OE� �� ,�|�� �0\�� �!64K��ԓrA� ��1 (M-7�!/50T�[PM��P�Th:1�C�#Pe� ��3�0� 5`M75cT"� �D8p� �0�Gc� u�4��i1-7'10i�1� Skd�7�j�?6�:-HS, � �RN�@�UB�f<�X�=m75sA*A�6an���!/CB�B2.6A �0;A�CIB�A��2�QF1�UB2�21� /70�S� �4��A��Aj1�3p���8r#0 B2\m*A@�C��;bi"i1K�u"A�~AAU� imm7c�7��ZA@I�@�Df��A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5�*A�EA�5B�4>\77
B7=Q�D�2�Q$BR�E7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E
"l7�@7�A
1�E�V$~`�W2%Q�R9ї@0L_�#����"Aȉ��b��H3s=rA/2�R5nR4�74rNUpQ1ZU�A�s\m9
1M92L2�!F!^Y�ps� 2ci��-?�qhimQ�t  w043�C��p2�mQ�r�H_ �H2�0�Evr�QHsXBSt62�q`s����� �<�Pxq350_*A3#I)�2�d�u0�@� �'4TX�0�pa3i1A3sQ25�c��st�r�VR1%e�q0
��j1��O2  �A�UEiy�.�‐ �0dCh20$CXB79#A��ᓄM Q1]�~�� 9�Q��?PQ��qA!P vs� 5	15aU����?PŅ���ဝQ9A6�zS*�7�qb5�1p����Q��00P(��V7]u�aitE1���À�p?7� !?�z��r=bUQRB1PM=�Q�a9��H��QQ�25L��������Q��@L���8ܰ��y00\}ry�"R2BL�t�N  ��� �1D�}�2�qeR�5���_b�3�X^]1m1lcqP1�a��E�Q� 5F����!5<���@M-16Q��  f���r��Q�e� ��8� PN�LT_�1��i1��9453��@�e�|�b1l>F1u *AY2�
��R8�Q����RJ�J3�D}T� 85
Qg�/0��*A!P@�*A�Ð𫿽�2ǿپ6t�6=Q���P�ȓ��� AQ�  g�*ASt]1^u�ajrI� B����~�|I�b��y&I�\m�Qb�I�uz��A�c3Apa9q� B6�S��S��m���}�8�5`N�N�  �(M���f1���6�����161��5�s`�SC��U��A�����5\set06c�����10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��� �5�B��B��h`�F� ��X0���A:���C�M�B��AZ��@��4�6i� ���� e�O�-	�� �f1��F �ᱦ�1pF�Y	���T6HL3���U66~`���U�dU�9D20Lf0��Qv � ��fjq��N���� ��0v
� ��i	�	.��72lqQ2�������� \chng�move.V��d����@2l_ar f	�f~��6��� ���9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�A]�,�V�1\�Qn�BJ�2W�EM!5�0��)�#:�64��F��e50S�\��0� =�PV���e�������E�����m7;shqQSH"U��)@��9�!A��(����� ,�}�ॲTR1!��,�60e=�4F�����2��	 R-����� ������Ж��4���LSR�)"�!l�OA��Q�) %!� 16�
U/��2�"2��E�9p���2X� SA�/i��'�
7F�H �@!B�0��D���5V ��@2cVE��p��T�2�pt갖�1L~E�#ȚF�Q��9E�#De/��RT��59���	�A��EiR������9\7m20�20��+�-u�19r4�`�E1�= `O9`�1"ae��O2��_$W}am4�1�4�3�/d1c_std��1)�!�`_T��r�_ 4\jdg�a�q�PJ%! ~`-�r�+bgB��#Nc300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W�"Ps A��e���� t�i�P�W.��c�@FX.�e�kE14��44�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2a���2A;_2��QW2��bF�(�V11�23`�`��X5�Ra21�!J*9�a:88J99X�l5�m1a첚��*���(85�&��� ����P6���R,!52&A����,fA9INfI50\u�z�OV
 �v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&� �P1��vB)e�m������1p� �1D˖}�27�F�KA�REL Use =S��FCTN��� J97�FA+�� (�Q޵�p%�)?�V�j9F?(�j�Rtk?208 "Km�6Q��y�j��iæPr�9��s#��v�krcfp�RCFt3���Q�¿kcctme�!M�E�g����6�mai�n�dV�� ��ru��kDº�c���o��L��J�dt�F ����.vrT�f������E%�!��5�FRj7%3B�K���UER�H�J�O  J�� (ڳF���F�q�Y�&T���p�F�z��19�tk vBr���V�h�9p�E�y�<�k������;�v���"CT��f�� ��)�
І��)�V	� 6���!��qFF��1 q���=�����O�?�$"����$��je���T?CP Aut�r�<�520 H5�J[53E193��9��+96�!8��9��	 n�B574��52�uJe�(�� Se%!�Y�����u��ma�Pqtool�ԕ��������conrel��Ftrol Re?liable�Rmv9CU!��H51���p�� a551e"<�CNRE¹�I�c�&��it�l\�sfutst "�UTա��"X�\u@��g@�i�6Q]V0�B$,Eѝ6A� �Q� )C���X��Yf�I�1�|6s@6i��T6AIU��vR�d�
$e%1��2�C58�E6���8�Pv�iV4OFH58�SOeJ� mvBM6E~O58�I�0�E�#+@ �&�F�0���F�P6a����)/++�</N)0�\tr1�����P �,�}ɶ�rmaski�msk�aA���Iky'd�h	A	�P�s�DisplayI�m�`v����J88G7 ("A��+Heůצprds��IϩǪ��h�0pl�2�R2Ƚ�:�Gt�@��PRD�TɈ�r�C�@Fm�8�D�Q�AscaҦ�� V<Q&��bVvbrl�eې@��^S��&5�Uf�j8710�yAl	��Uq���7�&��p�p��P^@�P�firmQ����Pp�2�=bk�6�r�3��6��otppl��PL���O�p<b�ac�q	��g 1J�U�d�J��gait_9e��Y�&��Qx���	�Shap��eration�0<��R67451j9:(`sGen�ms�42-f��r�p�5����2�rsgl�E��pp�G���qF�205p��5S���Ձ�retsdap�BP�O�\s�� "GCR�ö? ^�qngda�G��V��st2axU��A1a]��bad�_�>btputl/�&�|e���tplibB_��=�2.����5���gcird�v�slp���x�hex��v�rqe?�Ɵx�key��v�pm��x�us$�6�gcr��F���p���[�q27j92��v�ollismqS�k�9O�ݝ� (p#l.���t��p!o��A29$Fo8��cg7no~@�tptcls` �CLS�o�b�\�km�ai_
�s>�v�o�	�t�b���ӿ�E��H��6�1enu�501�[m��ut�ia|$calma�UR��CalMat�eT;R51%�i=1 ]@-��/V� ��Z��� �fq1�9 "K9�E�L����2m�C�LMTq�S#��et �LM3!} �F�c�nspQ�c���Oc_moq��� ��cc_e�����su���ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ���N�sve��C�clm��&Ao# �|$find�e�0STD� ter Fi�LANG���R���
��n3��z0C3en���r,���� ��J����� ���K ��Ú�=���_Ӛ���r� "FNDRК� 3��f��tguid�䙃N�."��J�tq�� �������@������J����_�� ����c��	m�Z�~�\fndr.��n#>
B2p��Z�C�P Ma�����3�8A��� c��6� ( ���N�B�������� 2�$�81��m_���"ex�z5 �.Ӛ��c��bS���efQ��	���RBT;�OPTN �+#Q�*$�r *$��*$r*$%/s#C��d/.,P�/0*ʲDPN��$���$*��Gr�$k Exc��'IF�$MASK��%93 H5�%H�558�$548 H�$4-1�$��#1(�$�0 E�$��$�-b�$���!UPDT �B�4�b�4�2�49��0�4a�3�9j0"Mx�49�4  ��4<�4tpsh���4<�P�4- DQ� �3 �Q�4�R�4�pR%0�2�r�4.b
E\���5�Ax�4��3adq\�5K979":E�ajO? l "DQ^E^�3i�Dq ��4ҲO) ?R�? ��q�5��T��3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F蠠�4��.�5y N|� �2il(in�4��31 JH1�2Q4�251ݠ�4rma	l� �3)�REo�Z_ �æOx����4��^F�?onorTf��7_ja��UZҒ4l�5rms�AU�Kkg���4�$HCd\�fͲ�eڱ�4�RE	M���4yݱ"u@�RE�R5932fO��47|Z��5lity,�Up��e"Dil\�5���o ��7987p�?�25 �3hk910 �3��FE�0=0P_>�Hl\mhm�5 ��qe�=$�^�
E�x�u�IAymptm�U0��BU��vste�y\ �3��me�b�DvI�[� Qu�:F�Ub�*_�
EL,�su��_ �Er��ox���4hGuse�E-�?�sn��������FE��,�box�����c݌,"� ������z��M��<g��pdspw)�	� �9���b���(��1���c��Y�R� � �>�P���W��������'�0ɵ�[���͂���  �� ,�@� ��A�bump�šf��B*�Box%��7Aǰ60�BBw�\��MC� (6�,f��t I�s� ST ��*��}B�����=w��"BBF
�>��`���)��\bb?k968 "�4��ω�bb�9va699����etbŠ��1X�����ed	�F�b�u�f� �sea""������'�\��,� ���b�ѽ�o6�H�
�x�$�f���!y�����Q[�! tpe�rr�fd� TP�l0o� Recov�,��3D��R64�2 � 0��C@}s�� N@��(U�rroč��yu2r��  �
  �����$$CLe� ��������������$z�_DI�GIT��������.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$j���+c:PROD�UCTM�0\PG/STKD��V&oho�zf99��D����$FEAT_�INDEX��xd���  �
�`ILECOM�P ;���#���`�cSETUPo2 <�e�b?�  N �a�c�_AP2BCK �1=�i  �)wh0?{%&c����Q�xe%�I �m���8��\� n����!���ȏW�� {��"���F�Տj��� w���/�ğS������ ���B�T��x���� ��=�үa������,� ��P�߯t������9� ο�o�ϓ�(�:�ɿ ^���Ϗϸ�G��� k� �ߡ�6���Z�l� �ϐ�ߴ���U���y� ���D���h��ߌ� ��-���Q������� ��@�R���v����)� ����_�����*�� N��r��7� �m�&�3\t�i
pP 2#p*.VRc�*��� /�ƗPC/1/F'R6:/].��/+T�`�/�/F%�/�,�`r/?�*.F��8?	H#&?e<x�/�?;STM �2��?�.K �?�=�iPendant? Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OpoO�O_:JPG _�J_�56_�O_�_�	�PANEL1.D	T�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�W�I��
TP�EINS.XML��0\���q�Custom T?oolbar	���PASSWOR�DyFRS:�\L�� %Pa�ssword Config���֏ e�Ϗ�B0���T�f� ���������O��s� �����>�͟b��[� ��'���K��򯁯� ��:�L�ۯp�����#� 5�ʿY��}��$ϳ� H�׿l�~�Ϣ�1��� ��g��ϋ� ߯���V� ��z�	�s߰�?���c� ��
��.��R�d��� ����;�M���q�� ����<���`������ %���I�������� 8����n���!� �W�{"�F �j|�/�S e��/�/T/� x//�/�/=/�/a/�/ ?�/,?�/P?�/�/�? ?�?9?�?�?o?O�? (O:O�?^O�?�O�O#O �OGO�OkO}O_�O6_ �O/_l_�O�__�_�_ U_�_y_o o�_Do�_ ho�_	o�o-o�oQo�o �o�o�o@R�ov ��;�_�� �*��N��G���� ��7�̏ޏm����&� 8�Ǐ\�돀��!��� E�ڟi�ӟ���4�ß X�j��������įS���w������B�#���$FILE_DG�BCK 1=���/���� ( �)
S�UMMARY.DyGL���MD:������Diag� Summary���Ϊ
CONSLOG�������D�ӱ�ConsoleO logE�ͫ���MEMCHECK�:�!ϯ���X�Me�mory Dat�a��ѧ�{)>��HADOW�ϣ����J���Shad�ow Chang�esM�'�-��)	FTP7Ϥ�3������Z�mmen�t TBD��ѧ0�=4)ETHERNET��������T�ӱEther�net \�figurationU��ؠ��DCSVRF��߽߫�����%��� verify� all��'�1P{Y���DIFF��p����[���%��diff]�������1R�9�K��� ����X��CH�GD������c��r����2ZAS�� ��GAD���k��z��FY3bI[�� �/"GAD���s/�����/*&UPDAT�ES.� �/��FORS:\�/�-Ա�Updates �List�/��PS�RBWLD.CM�(?���"<?�/Y�P�S_ROBOWEL��̯�?�?��?&� O-O�?QO�?uOOnO �O:O�O^O�O_�O)_ �OM___�O�__�_�_ H_�_l_o�_�_7o�_ [o�_lo�o o�oDo�o �ozo�o3E�oi �o���R�v ���A��e�w�� ��*���я`������ ���O�ޏs������ 8�͟\�����'��� K�]�쟁����4��� ۯj������5�įY� �}������B�׿� x�Ϝ�1���*�g��� ��Ϝ���P���t�	� ߪ�?���c�u�ߙ� (߽�L߶��߂��� (�M���q� ���6� ��Z������%���I� ��B�����2������h����$FIL�E_� PR� ���������MDONL�Y 1=.�� 
 ���q��� �������~% �I�m�2 ��h��!/�./ W/�{/
/�/�/@/�/ d/�/?�//?�/S?e? �/�??�?<?�?�?r? O�?+O=O�?aO�?�O �O&O�OJO�O�O�O_��O9_�OF_o_
VI�SBCKL6[�*.VDv_�_.POFR:\�_�^.P�Vision VD file�_ �O4oFo\_joT_�oo �o�oSo�owo�o B�of�o�+� ������+�P� �t������9�Ώ]� 򏁏��(���L�^�� �����5���ܟk� � ��$�6�şZ��~������
MR_GR�P 1>.L~��C4  B����	 W������*u����RHB ��2 ���� ��� ���B�����Z�l� ��C���D�������Ŀ���K��L6�mJ�p3F��5UT\Q�����ֿ G�,�FI�/E����.��9:�]�@�'��A&�#A�+�f�?�f�A���r��E�� F�@ �������J���NJk�H�9�Hu��F!��IP�s��?����(�9�<�9�89�6C'6<,6\b��+�&�(�`a�L߅�XȞ�A��� ��v���r������
� C�.�@�y�d����� ����������?�Z��lϖ�BH�� ��Ζ�������
0�P=��P�T���ܿ� �B���/ ��O@�33:��.��g&�@UUU�U���q	>u.�?!rX��	��-=[z�=��̽=V6<��=�=�=$�q�����@8��i7G��8��D�8@9!�7�:�����D�@ D�� �Cϥ��C���� ��Q�,/������/ M��/q��/�/�/�? ?:?%?^?p?[?�?? �?�?�?�? O�?�?6O !OZOEO~OiO�O�O�O �OW�ߵ��O$_�OH_ 3_l_W_�_{_�_�_�_ �_�_o�_2ooVoho So�owo�o�i��o�o �o��);�o_J �j������ �%��5�[�F��j� ����Ǐ���֏�!� �E�0�i�{�B/��f/ �/�/�/���/��/A� \�e�P���t������� �ί��+��O�:� s�^�p�����Ϳ��� ܿ� ��OH��o�
� ��~ϷϢ�������� ��5� �Y�D�}�hߍ� �ߞ��������o�1� C�U�y��߉��� ���������-��Q� <�u�`����������� ����;&_J \���������� ڟ�F�j4�� �������!/ /1/W/B/{/f/�/�/ �/�/�/�/�/??A? ,?e?,φ?P�q?�?�? �?�?O�?+OOOO:O LO�OpO�O�O�O�O�O �O_'__K_�o_�_ �_�_l��_0_�_�_�_ #o
oGo.okoVoho�o �o�o�o�o�o�o C.gR�v�� ���	���<� `�*<��`���� �ޏ��)��M�8�q� \�������˟���ڟ ���7�"�[�F�X��� |���|?֯�?����� 3��W�B�{�f����� ÿ���������A� ,�e�P�uϛ�b_���� �Ϫ_��߀�=�(�a� s�Zߗ�~߻ߦ����� ��� �9�$�]�H�� l������������ #��G�Y� �B����� ��z�������
ԏ:� C.gRd��� ���	�?* cN�r���� �/̯&/�M/�q/ \/�/�/�/�/�/�/�/ ?�/7?"?4?m?X?�? |?�?�?�?�?��O!O 3O��WOiO�?�OxO�O �O�O�O�O_�O/__ S_>_P_�_t_�_�_�_ �_�_�_o+ooOo:o so^o�o�op��o��  ��$��o�o �~������ �5� �Y�D�}�h��� ����׏����
� C�.�/v�<���8��� ���П����?�*� c�N���r�������� ̯��)��?9�_�q� ��JO�����ݿȿ� �%�7��[�F��j� �ώ��ϲ�������!� �E�0�i�T�yߟߊ� �߮��߮o�o��o>� t�>��b���� �������+��O�:� L���p����������� ��'K6oZ �Z�|�~���� �5 YDi�z ������/
/ /U/@/y/@��/�/�/ �/���/^/???Q? 8?u?\?�?�?�?�?�? �?�?OO;O&O8OqO \O�O�O�O�O�O�O�O�_�O7_��$FN�O ����VQ�
�F0fQ kP FL�AG8�(LRRM�_CHKTYP � WP��^P��WP�{QOM�P_�MIN�P�����P�  XNPS�SB_CFG �?VU ��_���S ooIU�TP_DEF_O/W  ��R&h�IRCOM�P8o��$GENOVRD7_DO�V�6�fl�THR�V d�ed�kd_ENBWo �k`RAVC_GR�P 1@�WCa X"_�o_1U <y�r���� �	��-��=�c�J� ��n��������ȏ� ���;�"�_�F�X���.ibROU�`FVX�P�&�<b&�8�?��埘��������  Da?�јs���@@g�B�7�p�)�ԙ���`WSMT�cG�mM����� �LQHOST�C�R1H���PĹ�at�SM���f�\���	1�27.0��1��  e��ٿ���� �ǿ@�R�d�vϙ�0��*�	anonymous���������F��X[�� � �����r����ߨߺ� ����-���&�8�[� I�π����� �1�C��W�y���`� r������ߺ������� %�c�u�J\n� ��������M� "4FX��i�� ����7//0/ B/T/���m/��/ �/�/??,?�/P? b?t?�?�/�?��?�? �?OOe/w/�/�/�? �O�/�O�O�O�O�O=? _$_6_H_kOY_�?�_ �_�_�_�_'O9OKO]O __Do�Ohozo�o�o�o �O�o�o�o
?o}_ Rdv���_�_o o!�Uo*�<�N�`� r��o������̏ޏ� ?Q&�8�J�\���>��ENT 1I��� P!􏪟  ����՟ğ����� ��A��M�(�v���^� ����㯦��ʯ+��  �a�$���H���l�Ϳ �����ƿ'��K�� o�2�hϥϔ��ό��� ��������F�k�.� ��R߳�v��ߚ��߾߀��1���U��y�<�?QUICC0��b�t����1�����%��2&���u�!?ROUTERv�R��d���!PCJO�G����!19�2.168.0.�10��w�NAME� !��!RO�BOTp�S_C�FG 1H�� ��Aut�o-starte�d�tFTP� ������  2D��hz��� �U��
//./�v ���/���/�/ �/�/�/�!?3?E?W? i?�/?�?�?�?�?�? �?���AO�?eO�/ �O�O�O�O�?�O�O_ _+_NO�OJ_s_�_�_ �_�_
OO.OoB_'o vOKo]ooo�oP_>o�o �o�o�oo�o5G Yk}�_�_�_� �8o��1�C�U�$ y��������ӏf��� 	��-�?����� Ə���ϟ���� �;�M�_�q���.�(� ��˯ݯ��P�b�t� ����m���������ǿ ٿ�����!�3�E�h� �{ύϟϱ����$� 6�H�J�/�~�S�e�w� �ߛ�jϿ�������� *߬�=�O�a�s��Y�T_ERR J�5
���PDUSI�Z  ��^J�����>��WRD �?t��  �guest }��%�7�I�[�m�$�SCDMNGRPw 2Kt�������V$�K��� 	P01.�14 8��  � y����B    ;������ ���������
 �������������~����C.gR�|���  i�  �  
��������� +��������
����l .r�
��"�l��� m
�d������_G�ROU��L�� e�	����07EQUPD  	ղ��J�TYa �����TTP_A�UTH 1M��� <!iPen'dany��6�Y�!KAREL�:*��
-KC�///A/ VISION SETT�/v/�"�/�/�/ #�/�/
??Q?(?:?��?^?p>�CTRL� N����5�
��.FFF9�E3�?�FRS�:DEFAULT��<FANUC� Web Server�:
���� �<kO}O�O�O�O�O���WR_CONFI�G O�� ��?��IDL_CP�U_PC@�B���7P�BHUM�IN(\��<TGNR_IO������P�NPT_SIM_�DOmVw[TPM�ODNTOLmV >�]_PRTY�X7R�TOLNK 1P����_o!o3oEo�Woio�RMASTE�lP��R�O_CFG�o�iUO��o�bCYCLE�o�d@_ASG 1Q����
 ko,>P bt����������sk�bNUM�����K@�`IPC�H�o��`RTRY�_CN@oR��bSGCRN����Q���1 �b�`�bR����Տ��$J23_�DSP_EN	�����OBPROqC�U�iJOGP�1SY@��8G�?�!�T�!�?*��POSRE�zVKANJI_�`��o_H�� ��T�L�6͕<����CL_LGP<��_���EYLOGG+IN�`���LANGUAGE� YF7RD ,w���LG��U�?�+���x� ������=P��'0���$ NMC:\�RSCH\00\���LN_DISP V��
������f��OC�R.RDzVT�A{�OGBOOK W
{��i��ii��X�����ǿٿ�����"��6	h�����e�?��G_BUFF 1%X�]��2	ա� ������������ !�N�E�W߄�{ߍߺ� �����������J�����DCS Z>r� =����^π+�ZE��������a�I�O 1[
{ ُ!� �!�1�C�U� i�y������������� ��	-AQcu@�������EfP/TM  �d�2 /ASew��� ����//+/=/�O/a/s/�/�/��S�EV����TYP�/??y͆��RS@"��×�F�L 1\
���� ��?�?�?�?�?�?�?�/?TP6��">>�NGNAM�ե��U`�UPS��GI�}�𑪅mA_LO{AD�G %��%DF_MOT�N���O�@MAXUALRM<��J��@sA�Q����WS ��@C �]m�-_���MPt2�7�^
{ رƭ	�!P�+ʠ�;_/��Rr�W�_�WU�W�_��R	o�_ o?o"ocoNoso�o�o �o�o�o�o�o�o; &Kq\�x�� �����#�I�4� m�P���|���Ǐ��� ֏��!��E�(�i�T� f�����ß��ӟ��� � �A�,�>�w�Z��� ����ѯ����د�� �O�2�s�^��������Ϳ���ܿ�'��BD�_LDXDISA�X@	��MEMO_{APR@E ?�+
 � *�~ϐπ�ϴ����������@I�SC 1_�+ ��IߨT��Q�c�� �߇��ߧ�����w�� ��>�)�b�t�[��� ��{����������:� ��I�[�/�������� ����o�����6!Z lS��s�� ��2�AS' �w����g���.//R/d/�_M?STR `�-w%�SCD 1am͠ L/�/H/�/�/?�/2? ?/?h?S?�?w?�?�? �?�?�?
O�?.OORO =OvOaO�O�O�O�O�O �O�O__<_'_L_r_ ]_�_�_�_�_�_�_o �_�_8o#o\oGo�oko �o�o�o�o�o�o�o" F1jUg�� �������B� -�f�Q���u�����ҏ�h/MKCFG �b�-㏕"LTA�RM_��cL�� σQ�N�><�METPUI�ǂ����)NDSP_CMNTh����|�  d�.���ς�ҟܔ|�POS�CF����PST�OL 1e'�4@�<#�
5�́5� E�S�1�S�U�g����� ��߯��ӯ���	�K� -�?���c�u�����|��SING_CHK�  ��;�ODA�Q,�f��Ç��D�EV 	L�	�MC:!�HSIZ�Eh��-��TAS�K %6�%$1�23456789� �Ϡ��TRIGw 1g�+ l6�%���ǃ�����8��p�YP[� ��EM_INF 1h3�� `)�AT&FV0E�0"ߙ�)��E0�V1&A3&B1�&D2&S0&C�1S0=��)A#TZ������H������A���AI�q�,���|���� ���� ������J���n���� ��W�����������" ����X��/���� e������0� T;x�=�as ��/�,/c=/b/ �/A/�/�/�/�/� �?���^?p?#/ �?�/�?s?}/�?�?O �?6OHO�/lO?1?C? U?�Oy?�O�O3O _�?�D_�OU_z_a_�_�O�NITOR��G �?5�   	�EXEC1Ƀ�R2*�X3�X4�X5�X����V7�X8�X9Ƀ �RhBLd�RLd�RLd�R Ld
bLdbLd"bLd.b�Ld:bLdFbLc2Sh2�_h2kh2wh2�h2��h2�h2�h2�h2*�h3Sh3_h3�R��R_GRP_SV� 1in���(ͅ�
�3�8��r��ۯ_MOx�_�D=R^��PL_N�AME !6���p�!Defa�ult Pers�onality �(from FD�) �RR2eq �1j)TUX)TsX��q��X dϏ 8�J�\�n��������� ȏڏ����"�4�F�@X�j�|������2'� П�����*�<�N�`�r��<�������� ү�����,�>�P�tb� �Rdr 1o�y� �\�, ��3���� @D��  ��?�����?x䰺��A'�6�����;�	lʲ	� �xJ������ �< ��"�� �(pK��K ��K=�*�J���J���JV���Zό����rτ́p@j�@T;f��f��ұ]�l���I��p�����������b��3���´  �
`�>�����bϸ�z��w꜐r�Jm��
� B�H�˱]Ӂt��q�	� p��  P�pQ�p�>�p|  Ъ�g����c�	'� �� ��I� ��  ����:��È
�È=����"�s��	�ВI�  �n @@B�cΤ�\��ۤ��t�q�y߁rN���  �'�����@2��@�����/��C��C�C�@� C������
��A�W�@<�*P�R�
h�B�b�A��j�����:����Dz۩��߹������j��( ?�� -��C�`��'�7�����q��Y����� �?�ff ��gy �����q�+q��
>+�  PƱj�(����7	����|�?���xZ�p<
6b�<߈;܍��<�ê<� �<�&Jσ�A�I�ɳ+���?ff�f?I�?&�k�@��.��J<?�`�q�.�˴ fɺ�/��5/���� j/U/�/y/�/�/�/�/��/?�/0?q��F �?l??�?/�?+)��?�?�E�� E��I�G+� F� �?)O�?9O_OJO�OXnO�Of�BL޳B� ?_h�.��O�O��%_�O L_�?m_�?�__�_�_x�_�_�
�h�Îg>��_Co�_`goRodo�o�GA�ds�q�C�o�o�o|����$]Hq�m��D��pC����pCHmZZ7t����6q�q��ܶN'�3�A�A�AR1�AO�^?�$��?�K�0±
�=ç>�����3�W
=�#�\W��e��9������{����<���(�B��u��=B�0�������	L��H�F�G����G��H��U`E���C��+���I#��I��HD��F��E��R�C�j=��
�I��@H�!�H�( E<YD0q�$��H� 3�l�W���{������� �՟���2��V�A� z���w�����ԯ���� ����R�=�v�a� �����������߿� �<�'�`�Kτ�oρ� �ϥ��������&�� J�\�G߀�kߤߏ��� ��������"��F�1� j�U��y������� �����0��T�?�Q�t���(�1��3/�E�����5�������q3�8�x����q4Mgs�&IB+2D�a���{�^ ^	������u%P2P7Q4_A���M0bt��R�������/   �/�b/P/�/ t/�/ *a)_3/�/�/�%1a?�/?;?8M?_?q?  �?�/��?�?�?�?O 2 �F�$�vGb��/�A��@�a�`�qC��C@�o�O2���O�F� DzH@��� F�P D�!��O�O�ys<O!_�3_E_W_i_s?��W�@@pZ.t2�2!2~
 p_�_�_�_	oo -o?oQocouo�o�o�o��o��Q ��+���1��$MSK�CFMAP  ��5� ��6�Q�Q"~�cONR�EL  
�q3�bEXCFE�NB?w
s1uXqF�NC_QtJOGO/VLIM?wdIpMr]d�bKEY?w�u]�bRUN�|�u��bSFSPDT�Y�avJu3sSIG�N?QtT1MOT��Nq�b_CE_�GRP 1p�5s\r���j����� T��⏙������<� �`��U���M���̟ ��🧟�&�ݟJ�� C���7�������گ��������4�V�`TC�OM_CFG 1�q}�Vp�����
�P�_ARC_\r�
jyUAP_CP�L��ntNOCHE�CK ?{ 	r��1�C� U�g�yϋϝϯ����������	��({NO_?WAIT_L�	u6M�NTX�r{�[�m�_ERRY�29sy3� &�������r�c� �촯T_MO��t��,�  �$�k�3�P�ARAM��u{��V[��!�u?��� =9@345678901��&��� E�W�3�c�����{������� �����=�UM_RSP�ACE �Vv��$ODRDSP����jxOFFSET�_CARTܿ�D�IS��PEN_FILE� �q��c����OPTION_�IO��PWOR�K v_�ms �P(�R�Q
�j.j	 ��Hj&�6$� RG_DS�BL  �5Js��\��RIENTkTO>p9!C��P�qfA� UT_SIM_D
r�b� �V� LCT w�w�bc��U)+$_P�EXE�d&RAT�p �vju�p��2X�j�)TUX)TX�>##X d-�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?O�H2�/oO �O�O�O�O�O�O�O�O_]�<^O;_M___q_ �_�_�_�_�_�_�_o����X�OU[�o(��(���$}o�, ���IpB` @D�  &Ua?�[cAa?��]a�]�DWcUa쪋l;��	lmb�`��xJ�`������a�<; ��`� ��b, �H(��H3k7�HSM5G�22�G���Gp
��
�!��'|, KCR�>�>q�Gs�uaT�3���  �4spBpyr  ]�o�*SB_�����j]��t�q� ��rna ��,���6  U��PQ��|N�M�,k�!�	�'� � ���I� �  {��%�=��ͭ�迋ba	���I  �n @� �~���p�����r �N	 W�  '!�o�:q�pC	 C�@�@sBq�|��� m�
S�!�h@ߐ�n�����Z�B	 �A8���p� �-�qbz�P��t�_�������( �� -��恊�n�ڥ[A]Ѻ�b4�'!���(p �?�fAf� ��
����O�Z�R��8��z���>N΁  Pia��(�� ��@���ک�a�c�dF#/?����x�����<
6b<߈�;܍�<�ê�<� <�&�o&�)�A�lcΐIƾ*�?fff?�?y&c���@�.u��J<?�`�� Yђ^�nd��]e��[g ��Gǡd<����1�� U�@�y�dߝ߯ߚ��� �߼�	���-�������&��"�E�� E���G+� F� ������������&���J�5��bB��A T�8�ђ��0�6���>� ��J�n�7��[mx�0��h��1��>�M�I`
�@��A�[��C-�)��?���� /�
YĒ��Jp��vav`#CH/�������}!@I�Y�'��3A�A�AR�1AO�^?�$��?����±�
=ç>�����3�W
=�#�����+e��ܒ������{�����<��.(��B�u��=�B0�������	�*H�F��G���G���H�U`E����C�+�-I#��I��HD��F��E���RC�j=U>
�I��@H��!H�( E<YD0/�?�?�? �?�?O�?3OOWOBO TO�OxO�O�O�O�O�O �O_/__S_>_w_b_ �_�_�_�_�_�_�_o o=o(oaoLo�o�o�o �o�o�o�o�o' $]H�l��� ����#��G�2� k�V���z���ŏ��� ԏ���1��U�g�R� ��v�����ӟ��������-��(���������a�����Q�c�,!3�8��}���,!4Mgs8����ɢIB+կ���a���{� ��A�/�e�S���w�J�P!�P��������7��ӯ�ϑ�R9�Kτ�oχϓϥ�  ���χ���� )��M����������{߉ߛ���ߒߤ�p������  )�G�q�_���2� F�$�&Gb	���n�[ZjM!C�s�@j/�A�S�~��F� Dz����� F�P DC��W����)������������x?̯��@@
9�RE�E��E��
 v��� ����*<pN`�*P �������1��$PA�RAM_MENU� ?-���  DEFPULSEl�	WAITTM�OUT�RCV�� SHEL�L_WRK.$CUR_STYL�;,OPT�/�PTB./("C�R?_DECSN��� ,y/�/�/�/�/�/�/ ?	??-?V?Q?c?u?��?�USE_PR_OG %�%�?\�?�3CCR������7_HOST !�!�44O�:AT̰�?PCO)ARC|�O�;_TIME��XB�  �GD�EBUGV@��3G�INP_FLMS�K�O�IT`��O�EP+GAP �L��#[�CH�O�HTYPE
����?�?�_�_ �_�_�_oo'o9obo ]ooo�o�o�o�o�o�o �o�o:5GY� }����������1�Z��EWOR�D ?	7]	�RS`�	PNS2�$��JOE!>��TEs@WVTRA�CECTL 1xv-�� ���Ӱ��ɆDT� Qy-����D � �� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� T�(�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_j��_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�_����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv��������//"#�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �" |"DEFSPD |�,�!!J �8 IN~ TRL }�-�" 8�(IPE__CONFI� ~g%��g!�$��$�"8 LID�#��-74GRP 1��7Q!�#!A ���&ff"!�A+33D�� �D]� CÀ SA@+6�!�" d�$�9�9*1*0� 	� +9�-+6�? ��	C�?�;B@3AO��?OIO3OmO"!>�?T?�
5�O�O��N�O =��=#�
�O_�O_J_ 5_n_Y_�O}_�_y_�_<�_�_  Dzco" 
oBo�_Roxoco �o�o�o�o�o�o�o�>)bM��;�
V7.10be�ta1�$  �A�E�rӻ�A " �p?!G���q>���r�܁0�q�ͻqBQ��qA\�p�q�4T�q�p�"�BȔ 2�D�V�h�w��p�?�?)2{ȏw�׏ ���4��1�j�U��� y�����֟������ 0��T�?�x�c����� ��ү����!o�,�ۯ P�;�M���q�����ο ���ݿ�(��L�7��p�+9��sF@  �ɣͷϥ�g%����� �+�!6I�[߆����� �ߵߠ���������!� �E�0�B�{�f��� ����������A� ,�e�P���t������� �����=(a L^������ �'9$]�Ϛ� �ϖ�������/ <�5/`�r߄ߖߏ/> �/�/�/�/�/?�/1? ?U?@?R?�?v?�?�? �?�?�?�?O-OOQO <OuO`O�O�O�O�O�� �O_�O)__M_8_q_ \_n_�_�_�_�_�_�_ o�_7oIot���o �o���o�o�o(/! L/^/p/�/{*o�� �������A� ,�e�P�b��������� �Ώ��+�=�(�a� L���p������Oߟ� ��� �9�$�]�H��� l�~�����ۯƯ��� #�No`oro�on��o�o �o�oԿ���8J \ng����vϯϚ� ������	���-��Q� <�u�`�r߫ߖ��ߺ� ������;�M�8�q� \��������z���� ��%��I�4�m�X��� |�����������:� L�^���Z������� ����$�6�H� Swb���� ���//=/(/a/ L/�/p/�/�/�/�/�/ ?�/'??K?]?H?�? ��?�?f?�?�?�?O �?5O OYODO}OhO�O �O�O�O�O�O&8J 4_F_����_�_� �_�_"4-o�O*o coNo�oro�o�o�o�o �o�o)M8q \������� ��7�"�[�m��?�� ��R�Ǐ���֏�!� �E�0�i�T���x��� �����_$_V_ �2��l_~_�_�����R�$�PLID_KNO�W_M  �T������SoV ��U͠�U��
�� .�ǟR�=�O�����m�ӣM_GRP 1���!`0u��T@Rٰo�ҵ�
�� �Pзj��`���!� J�_�W�i�{ύϟϱ����������߱�MR������T��s�w� s��ߠ޴߯߅��� �߻�����A���'� ���������� ����=���#����������}������S��S�T��1 1��U�# ���0�_ A .��,>Pb� �������3 (iL^p��P���2*N���<-/3/)/;/M/4f/x/�/�/5�/�/�/�/A6??(?:?7S?e?w?�?8�?�?�?��?MAD  �d#`PAR�NUM  �w�%OSCH?J �ME
�G`A�Iͣ�EUPD`OrE
a�OT_CMP_��B@�P�@'˥TER_wCHK'U��˪?R$_6[RSl�¯��G_MOA@�_�U_�_~RE_RES_G ��>�oo8o+o \oOo�oso�o�o�o�o��o�o�o�W �\ �_%�Ue Baf�S � ����S0�� ��SR0��#��S�0 >�]�b��S�0}������RV 1�����rB�@c]��t�(�@c\����D�@c[�$���RT?HR_INRl�DA���˥d,�MASS69� ZM�MN8�k��MON_QUEUE ���˦��x�� RDNPUbQN8{�P[��END���_�ڙEXE�ڕ�@B�E�ʟ��OPTI�OǗ�[��PROG�RAM %��%���ۏ�O��TAS�K_IAD0�OCFG ���tO��Š�DATA���Ϋ@��27�>�P�b� t���,�����ɿۿ������#�5�G���IN+FOUӌ������ �ϭϿ��������� +�=�O�a�s߅ߗߩ߀���������^�jč�� yġ?PDI�T �ίc���W�ERFL
��
RGADJ �n�A����?����@�~��IORITY{��QV���MPDSP(H�����Uz����oOTOEy�1�R� (!AF4��E�P]���!t�cph���!u�d��!icm���ݏ6�XY_ȡ�R��ۡ)� a*+/ ۠� W:F�j��� ���%7[�B�*��POR�T#�BC۠�����_CARTRE�P
�R� SKSTyAz��ZSSAV����n�	2500H863���r�$�!�R�����q�n�}/�/�'� UR�GE�B��rYWFF� DO{�rUVWV���$�A�WRUP_�DELAY �|R��$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?�3AQSKIP!�vn�l#x 	1/ +O+ OROdOvO9Hn� �O�G�O�O�O�O�O_ �O_D_V_h_._�_z_ �_�_�_�_�_
o�_.o @oRoovodo�o�o�o �o�o�o�o*<�Lr`���n��?$RCVTM������pDCR!��LЈqCl�f�C��C��>�?�A�>:���<l��4M�b�����O�
�n�������{�4Oi��O� <
6b<�߈;܍�>u�.�?!<�&{�b�ˏݏ��8� ����,�>�P�b�t� ��������Ο���ݟ ��:�%�7�p�S��� ���ʯܯ� ��$� 6�H�Z�l�~������� ƿ���տ���2�D� '�h�zϽ��ϰ����� ����
��.�@�R�d� Oψߚ߅߾ߩ����� ����<�N��r�� ������������ &�8�#�\�G�����}� ����������S�4 FXj|���� �����0T ?x�u���� '//,/>/P/b/t/ �/�/�/�/�/�/�? �/(??L?7?p?�?e? �?�?��?�? OO$O 6OHOZOlO~O�O�O�? �?�O�O�O�O __D_ V_9_z_�_�?�_�_�_ �_�_
oo.o@oRodo�vo�X�qGN_AT�C 1�� �AT&FV0�E0�kATD�P/6/9/2/�9�hATA�n�,AT%G1�%B960�iW+++�o,�aH�,�qIO_TYPOE  �u�sn_��oREFPOS1� 1�P{ x	�o�Xh_�d_� ����K�6�o�
����.���R����{{2 1�P{���؏�V�ԏz����q3 1��$�6�p��ٟ�>��S4 1������˟���n���%�S5 1�<�N�`������<���S6 1� ѯ���/�����ѿO�S7 1�f�x����ĿB�-�f��S8 1�����Y��������y�SMASK ;1�P  
9�G�N�XNOM���a�~߈ӁqMOTE � h�~t��_CFG� ������рrP?L_RANG�ћQ���POWER 壡e��SM_�DRYPRG �%i�%��J��TA�RT �
�X�U?ME_PRO'�9����~t_EXEC_?ENB  �e��GSPD������c���TDB���RM\��MT_!�T�����`OBOT_NAME i����iOB_OR�D_NUM ?�
�\qH863  �T���������bPC_T�IMEOUT�� �x�`S232��1���k LT�EACH PEN�DAN �ǅ��}���`Main�tenance �Cons�R}�m
"�{�dKCL/C�g��Z ��n� �No Use�}�	��*NPO���х����(CH_L���̥���	�mMA�VAIL��{����ՙ�SPACE1w 2��| d@��(>��&���p���M,8�?� ep/eT/�/�/�/�/ �W//,/>/�/b/�/ v?�?Z?�/�?�9�e�a �=??,?>?�?b?�? vO�OZO�?�O�O�Os
�2�/O*O<O �O`O�O�_�_u_�_�_�_�_[3_#_5_G_ Y_o}_�_�o�o�o�o�o[4.o@oRo dovo$�o�o��� �"�	�7�[5K] o��A����	�@̏�?�&�T�[6h� z�������^�ԏ����&��;�\�C�q�[7 ��������͟{��� "�C��X�y�`���[8����Ưدꯘ�� 0�?�`�#�uϖ�}ϫ��[G �i�� �ϋ
G�  ����$�6�H�Z�l�~� ���8 ǳ�����߈��d(���M�_� q���������� �?���2�%�7�e�w� ���������������� ���!�RE�W��� ��������?Q `�� @0��ߖrz	�V_���� �
/L/^/|/2/d/�/ �/�/�/�/�/?�/�/ �/*?l?~?�?R?�?�? �?�?�?�?�?2O�?�
��O[_MOD�E  �˝IS ����vO,* ϲ�O-_��	M_v_�#dCWORK_A�D�M9�P%aR  ��ϰ�P{_��P_INTVAL��@����JR_OPoTION�V �E�BpVAT_GR�P 2�����(y_Ho � e_vo�o�oYo�o�o�o �o�o*<�bOo NDpw����� �	���?�Q�c�u� ����/���ϏᏣ��� �)�;���_�q����� ����O�ɟ���՟ 7�I�[�m�/������� ǯٯ믁��!�3��� C�i�{���O���ÿտ ���ϡ�/�A�S�e� 'ωϛϭ�oρ����� ��+�=���a�s߅� Gߕ߻����ߡ��� '�9�K�]��߁��� ��y����������5��G�Y��E�$SCAN_TIM�AYue�w�R �(ӿ#((�<0.a�aPaP
Tq>��Q��oa�����OOE2/��:	d/"JaR��WY��^����^R^	r  �P��� �  8�P�	�D��GY k}������p��Qp/�@/R//)P;��o\T��Qpg-�?t�_DiKT��>[  � lv% ������/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OWW�#�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_olO~Od+No`oro �o�o�o�o�o�o�o &8J\n������u�  0 �"0g�/�-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ��$o��˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�����Do�������� ҿ�����,�>�P� b�tφϘϪϼ�����0����w
�  58� J�\�n߀ߒߜկ��� ������	��-�?�Q��c�u����� ��-����� �2� D�V�h�z���������a���������&� ��%	12345678�"� 	��/�� `r���� ����(:L ^p������ � //$/6/H/Z/l/ ~/��/�/�/�/�/�/ ? ?2?D?V?h?�/�? �?�?�?�?�?�?
OO .O@Oo?dOvO�O�O�O �O�O�O�O__*_YO N_`_r_�_�_�_�_�_ �_�_ooC_8oJo\o no�o�o�o�o�o�o�o o"4FXj|@�������� �	��s3�E�W�{�Cz  Bp��_   ��2����z�$SCR_G�RP 1�(�U�8(�\x}^ @ � 	!�	 ׃ ���"�$� ��-���+��R�w�����D~�����#�����O���M-10iA 8909�905 Ŗ5 M61C >4��Jׁ
� ���0�@����#�1�	"�@z�������¯Ҭ ���c���O� 8�J�������!�p����ֿ��B�y�!��������A��$χ  @��<� �R�?��d���Hy�u�O���F@ F�`�� ��ʿ�϶�������%� �I�4�m��<�l�0�ߕߧ߹�B���\� ���1��U�@�R�� v���������@��;���*<=�
F����?�d�<�>m�̎��@�:��� B���ЗЙ����EL_DEFAU�LT  �����B�M�IPOWERFL�  �$1 W7FDO $���ERVENT 1O�����"�p�L!DUM_E�IP��8��j!?AF_INE ��=�!FT���!��4 ���[!RPC_OMAIN\>�J��nVISw=����!TP�P�U��	d�?/!
�PMON_PROXY@/�e./�/"�Y/�fz/�/!R?DM_SRV�/�	9g�/#?!R C?��h?o?!
pM�/�i^?�?!R�LSYNC�?8��8�?O!ROS�.L�4�?SO"wO �#DOVO�O�O�O�O�O _�O1_�OU__._@_ �_d_v_�_�_�_�_o��_?oocoiICE�_KL ?%y� (%SVCPRG1ho8��e���o"�m3�o�o�`4 "�`5(-�`6PU�`7x}�`���l	9��{�d:?��a �o��a�oE��a�om� �a���aB���aj 叟a���a�5��a �]��a����a3��� �a[�՟�a�����a�� %��aӏM��a��u��a #����aK�ů�as�� �a��mob�`�o�`8� }�w�������ɿ��� ؿ���5�G�2�k�V� ��zϳϞ�������� ��1��U�@�y�dߝ� �ߚ��߾������� ?�*�Q�u�`���� ���������;�&� _�J���n������������sj_DEV �y	�MC�:P�_O�UT",REC 1�Z� d �  	 	�������
 �PJ��%6 (�&a�[w�,ݚ*  T J- �- �A�- c| �P�����/ /B/0/f/x/Z/�/�/ �/�/�/�/�/?�/? P?>?t?b?�?�?�?�? �?�?�?OOOLO:O pO�OdO�O�O�O�O�O �O�O$__H_6_X_~_ l_�_�_�_�_�_�_�_  ooDo2oTozo\o�o �o�o�o�o�o�o. R@vd��� �},����4� "�X�F�|���p����� ֏ď����0��@� f�T���x�����ҟ� Ɵ���,��<�b�P� ��h�z������ί� �(�:��^�L�n�p� ������ܿ�п� � 6�$�Z�H�jϐ�rϴ� �����������2�D� &�h�Vߌ�z߰ߞ��� ��������
�@�.�d��R��ZjV 1��w P�m��	�>   y��
TYPEV�FZN_CFGw ��d�7�GRP �1�A�c ,B� A� D;� �B���  B4~RB21/HELL:�(
�� X����%RSR����E 0iT�x��� ���/Se~w�  ��%w�����b#������犍2#�d����H�K 1���  �k/f/x/�/�/�/�/ �/�/�/??C?>?P?�b?�?�?�?�?��OM�M ����?��FTOV_ENB ����+�HOW_RE�G_UIO��IM/WAITB�JK�OUT;F��LIT�IM;E���OV�AL[OMC_UNI�TC�F+�MON_�ALIAS ?e~�9 ( he�� _&_8_J_\_��_�_ �_�_�_j_�_�_oo +o�_Ooaoso�o�oBo �o�o�o�o�o'9 K]n���� t���#�5��Y� k�}�����L�ŏ׏� �����1�C�U�g�� ��������ӟ~���	� �-�?��c�u����� ��V�ϯ������ ;�M�_�q�������� ˿ݿ����%�7�I� ��m�ϑϣϵ�`��� ����ߺ�3�E�W�i� {�&ߟ߱������ߒ� ��/�A�S���w�� ���X�������� ��=�O�a�s���0��� ����������'9 K]����b ���#�GY k}�:���� ��/1/C/U/ /f/ �/�/�/�/l/�/�/	? ?-?�/Q?c?u?�?�? D?�?�?�?�?O�?)O ;OMO_O
O�O�O�O�O �OvO�O__%_7_�C��$SMON_D�EFPRO ����`Q� *SYS�TEM*  d=�OURECALL� ?}`Y ( ��}4xcopy� fr:\*.*� virt:\t�mpback�Q=�>192.168�.4�P46:8144 �R�_�_�_�K}5�Ua�_�_�V�_�goyo�o}9�Ts:�orderfil.dat.l@oVo�o��o}0�Rmdb:+o�oRc�odv� a�_2o?U��
� o��Sod�v����o �o6Q���+ ƏO`�r����*�<� �ޟ���'���K��\�n����
xyz�rate 61 �+�=�O�����|����6788 �� үc�u�������5�6� ٿ����"���5�ѿ�b�tφ��6����e�mp:�6976 �W����ύ�.��*.d������`�r߄ߗ�1 +�=�O������ �)�������c�u�� ����5���������� "Ͻ�����b�t����� ����:�V����������6 ��gy� ���9�T���	� �@��cu���- ?����/�� N_/q/�/��1� �/�/?&�/J[? m??��7/��?�? �?/"/�?F/�?iO{O �ߠ�2ODOVO�O�O_�Ř284>��Oa_ s_�_�/�/3?4Y�_�_ �_?"?�_5X�_boto��o�ϫ_��8Q392 Wo�o�o�o߹o�j �oas��O��<N ���_(_�s�� c�u����_�_5o�gُ ���o"o���hяb��t������$SNP�X_ASG 1��������� P 0 �'%R[1]�@1.1����?���%֟��&�	�� \�?�f���u������� �ϯ��"��F�)�;� |�_�������ֿ��˿ ���B�%�f�I�[� ��Ϧ��ϵ������� ,��6�b�E߆�i�{� �ߟ����������� L�/�V��e���� ��������6��+� l�O�v����������� ����2V9K �o������ �&R5vYk �����/�� <//F/r/U/�/y/�/ �/�/�/?�/&?	?? \???f?�?u?�?�?�? �?�?�?"OOFO)O;O |O_O�O�O�O�O�O�O _�O_B_%_f_I_[_ �__�_�_�_�_�_�_ ,oo6oboEo�oio{o �o�o�o�o�o�o L/V�e��� �����6��+��l�O�v�������PA�RAM ���}�� �	���P����OF�T_KB_CFG�  ヱ���PI�N_SIM  ���C�U�g������RVQSTP_DSB,�򂣟�����SR �/�� �&  ULTI�ROBOTTAS�K�����TOP�_ON_ERR � ���PT�N /�@��A	�RINGo_PRM� ���VDT_GRP �1�ˉ�  	 ������������Я� ����*�Q�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߣߠ߲� ����������0�B� i�f�x�������� �����/�,�>�P�b� t��������������� (:L^p� ������  $6HZ�~�� �����/ /G/ D/V/h/z/�/�/�/�/ �/�/?
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8___\_��VP�RG_COUNT���@���REN�BU��UM�S��__�UPD 1�/�8  
s_�oo *oSoNo`oro�o�o�o �o�o�o�o+&8 Jsn����� ����"�K�F�X� j���������ۏ֏� ��#��0�B�k�f�x� ��������ҟ����� �C�>�P�b������� ��ӯί�����UYSDEBUG�P��P�)�d�YH�SP�_PASS�UB�?Z�LOG �V�U�S)�#��0�  ��Q)�
�MC:\��6���_MPC���U���Q�ñ8� �Q�SA/V �����ǲ�&�ηSV;�T�EM_TIME �1��[ (m�7�&�4:�}YT1S�VGUNS�P�U'��U���ASK_?OPTION�P�U��Q�Q��BCCF�G ��[u� 8n�A�a�`a�gZ o��߃ߕ��߹����� ��:�%�^�p�[�� ������� ����� 6�!�Z�E�~�i���������&�������& 8��nY�}� ?��ԫ ��( L:p^��� ����/ /6/$/ F/l/Z/�/~/�/�/�/ �/�/�/�/2?8 F? X?v?�?�??�?�?�? �?�?O*O<O
O`ONO �OrO�O�O�O�O�O_ �O&__J_8_n_\_~_ �_�_�_�_�_�_o�_  o"o4ojoXo�oD?�o �o�o�o�oxo. TBx��j�� ������,�b� P���t�����Ώ��ޏ ��(��L�:�p�^� ������ʟ��o� �6�H�Z�؟~�l��� ����د���ʯ �� D�2�h�V�x�z���¿ ���Կ
���.��>� d�Rψ�vϬϚ��Ͼ� ������*��N��f� xߖߨߺ�8������� ��8�J�\�*��n� ������������"� �F�4�j�X���|��� ����������0 @BT�x�d�� ���>,N tb������ /�(//8/:/L/�/ p/�/�/�/�/�/�/�/ $??H?6?l?Z?�?~? �?�?�?�?�?O�&O 8OVOhOzO�?�O�O�O �O�O�O
__�O@_._ d_R_�_v_�_�_�_�_ �_o�_*ooNo<o^o �oro�o�o�o�o�o�o  J8n$O� ����X����4�"�X�B�v��$T�BCSG_GRP� 2�B���  �v� 
? ?�  ���� ��׏�������1���U�g�z���ƈ�d�, ���?v�	� HC��d�>󙚲�e�CL  �B���Пܘ��ݸ��\)��Y g A�ܟ$�B�g�FB�Bl�i�X�ɼ�|��X��  D	J���r�����C����$үܬ���D�@v�=� W�j�}�H�Z���ſ���������v�	V3.00���	m61c�	�*X�P�u�g�p�>ə��v�(:�� ���p͟�  O�����p�����z�JC�FG �B���� ������r����=��=� c�q�K�qߗ߂߻ߦ� �������'��$�]� H��l�������� ����#��G�2�k�V� ��z����������� ���p*<N��� l������� #5GY}h� ���v�b��>�/ / /V/D/z/h/�/�/ �/�/�/�/�/?
?@? .?d?R?t?v?�?�?�? �?�?O�?*OO:O`O NO�OrO�O�O��O�O �O_&__J_8_n_\_ �_�_�_�_�_�_�_�_ �_oFo4ojo|o�o�o Zo�o�o�o�o�o�o B0fT�x�� �����,��P� >�`�b�t�����Ώ�� �����&�L��Od� v���2�����ȟʟܟ � �6�$�Z�l�~��� N�����دƯ�� � 2��B�h�V���z��� ��Կ¿����.�� R�@�v�dϚψϪ��� ��������<�*�L� N�`ߖ߄ߺߨ����� ��������\�J�� n���������� "���2�X�F�|�j��� ������������ .TBxf��� ����>, bP�t���� �/�(//8/:/L/ �/�ߚ/�/�/h/�/�/ �/$??H?6?l?Z?�? �?�?�?�?�?�?O�? ODOVOhO"O4O�O�O �O�O�O�O
_�O_@_ ._d_R_�_v_�_�_�_ �_�_o�_*ooNo<o ro`o�o�o�o�o�o�o �o&�/>P�/ �������� �4�F�X��(���|� ����֏����Ə0� �@�B�T���x����� ҟ������,��P� >�t�b����������� ����:�(�^�L� n�������2d��� ��̿�$�Z�H�~�l� �ϐ��������Ϻ� � �0�2�D�zߌߞ߰� j����������
�,� .�@�v�d����� ��������<�*�`� N���r����������� ��&J\�t ��B����� �F4j|���^����/� s 2 6# 6&�J/6"�$TBJO�P_GRP 2���� O ?�X,i#�p,�� �x/J� �6$� � �< �z� �6$ @2 ��"	 �C�� >�&b  Cق'�!�!>���
559�>�0+1�33=��CL� ff�f?+0?�ffB@� J1�%Y?d7�.��/�>��2\)�?0�5���;���hCY� �  �@� �!B�  A��P?�?�3EC� � D�!�,�0*B�Oߦ?�3JB��
�:���Bl�0���0�$�1�?O6!A�ϙ�AДC�1D�G6�=q�E6O0��p��B�Q�;��A�� ٙ7�@L3D	�@�@�__�O�O>B�\pJU�OHH�1ts�A�@33@?1� C��� �@�_�_&_8_>G��D�UV_0�LP<�Q30<{�zR� @�0�V�P!o3o�_<o RifoPo^o�o�o�oRo �o�o�o�oM(�o�l�p~��p4��6&�q5	V3�.00�#m61c�$*(��$1!6��A� Eo��E��E���E�F���F!�F8���FT�Fqe\�F�NaF����F�^lF����F�:
F�)�F��3G��G��G���G,IR�CH`��C�dTDU��?D��D���DE(!/E\��E��E�h��E�ME���sF`F+'�\FD��F`�=F}'�F���F�[
F����F��M;S@;WQ��|8�`rzQ@/&�8�6&<���1�w�^$ESTP?ARS  *({ �_#HR��ABLE� 1�p+Z�6#D|�Q� � 1�|�|��|�5'=!|�	|�
�|�|�˕6!|��|�|���RDI��z!ʟܟ� ��$���O������¯ԯH�����S��x# V� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������U-����Ĝ P�9�K�]�o��-�?��Q�c�u���6�NUM�  �z!�� >  Ȑ����_?CFG ������!@b IMEBF_TT����x#��a�GVER��b�w�a��R 1�p+
 (I3�6"1 ��   6!���������� �9� $�:�H�Z�l�~����� ����������^$��_��@x�
b M�I_CHANm� �x� kDBGLV�;0o�x�a!n ET�HERAD ?*�� �y�$"x�\&n ROUT��!p*!*�?SNMASK�x#>�255.h��fx^$OOLOF/S_DI��[ՠ	�ORQCTRL �p+;/���/ +/=/O/a/s/�/�/�/ �/�/��/�/�/!?���PE_DETAI���PON_SV�OFF�33P_M�ON �H�v�2�-9STRTCHK� ���42VTCOMPATa8��24:0FPROG� %�%MU�LTIROBOT�TO!O06�PLA�Y��L:_INST+_MP GL7YD�US���?�2LCK��LPKQUICKM�Et �O�2SCRE��@�
tps��2�A�@�I��@�_Y���9�	SR_�GRP 1��/ ���\�l_ zZg_�_�_�_�_�_�^�^�oj�Q'ODo/o hoSe��oo�o�o�o �o�o�o!WE {i�������	123456�7��!���X�E1��V[
 �}i�pnl/a�gen.htmno���������ȏ~�Pan�el setup̌}�?��0�B�T�f� ��񏞟�� ԟ���o����@�R� d�v������#�Я� ����*���ϯůr� ��������̿C��g� �&�8�J�\�n���� �϶���������uϣ� ��F�X�j�|ߎߠ�� ��;�������0�B�|��*NUALRMb@oG ?�� [� ������������ � �%�C�I�z�m��������v�SEV  ����t�ECFG Ձ=]/Ba}A$   B�/D
 ��/C�Wi {�������� PRց; P�To\o�I�6?K0(%����0�� ���//;/&/L/�q/\/�/�/�/l�D ��Q�/I_�@H�IST 1ׁ9 � (  ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153,1 Ec0p?�?�?��?/C�� >?P=962n?�?
OO.O�?�?�136c?|O�O�O �OAOSO�?�O__0_ �O�O_Lu_�_�_�_:_ �/�_�_oo)o;o�_ _oqo�o�o�o�oHo�o@�o%7I~��a 81�ou����� �o���)�;�M�� q���������ˏZ�l� ��%�7�I�[��� ������ǟٟh���� !�3�E�W�������� ��ïկ�v���/� A�S�e�Pb������ ѿ������+�=�O� a�s�ϗϩϻ����� ��ߒ�'�9�K�]�o� ��ߥ߷��������� ��#�5�G�Y�k�}�� ������������� 1�C�U�g�y���v��� ��������	�? Qcu��(�� ��)�M_ q���6��� //%/�I/[/m// �/�/�/D/�/�/�/? !?3?�/W?i?{?�?�? �?�����?�?OO/O AOD?eOwO�O�O�O�O NO`O�O__+_=_O_ �Os_�_�_�_�_�_\_ �_oo'o9oKo�_�_ �o�o�o�o�o�ojo�o #5GY�o}������?��$�UI_PANED�ATA 1������  	�}�0�B�0T�f�x��� )���� mt�ۏ����#�5� ��Y�@�}���v����� ן�������1��U�pg�N������ �1��Ïȯگ���� "�u�F���X�|����� ��Ŀֿ=������ 0�T�;�x�_ϜϮϕπ�Ϲ������,ߟ� M��j�o߁ߓߥ߷� �����`��#�5�G� Y�k��ߏ������ ��������C�*�g� y�`���������F�X� 	-?Qc��� �߫���� ~;"_F��| �����/�7/ I/0/m/�����/�/�/ �/�/�/P/!?3?�W? i?{?�?�?�??�?�? �?O�?/OOSOeOLO �OpO�O�O�O�O�O_ z/�/J?O_a_s_�_�_ �_�O�_@?�_oo'o 9oKo�_oo�oho�o�o �o�o�o�o�o#
G Y@}d��&_8_ ����1�C��g� �_��������ӏ��� ^���?�&�c�u�\� ������ϟ���ڟ� )��M��������� ��˯ݯ0�����7� I�[�m���������� ٿ�ҿ���3�E�,� i�Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#��� ���� ��$�6��Z� A�~�e�w������ �����2��V�h�O������v�p��$UI�_PANELIN�K 1�v��  � � ��}1234?567890���� 	-?G ���o �����a��@#5G�	����4p&���  R� ����Z��$/ 6/H/Z/l/~//�/�/ �/�/�/�/�/
?2?D? V?h?z??$?�?�?�? �?�?
O�?.O@OROdO vO�O O�O�O�O�O�O _�O�O<_N_`_r_�_�_�0,���_�X�_ �_�_ o2ooVohoKo �ooo�o�o�o�o�o�o ��,>r}��� �������� �/�A�S�e�w���� ����я���tv�z� ���=�O�a�s��� ����0S��ӟ���	� �-���Q�c�u����� ��:�ϯ����)� ��M�_�q��������� H�ݿ���%�7�ƿ [�m�ϑϣϵ�D��� �����!�3�Eߴ_i� {�
�߂����߸��� ���/��S�e�H�� ��~��R~'�'�a� �:�L�^�p������� �������� ��6 HZl~���#� 5��� 2D�� hz�����c �
//./@/R/�v/ �/�/�/�/�/_/�/? ?*?<?N?`?�/�?�? �?�?�?�?m?OO&O 8OJO\O�?�O�O�O�O �O�O�O[�_��4_F_ )_j_|___�_�_�_�_ �_�_o�_0ooTofo ��o��o��o�o�o ,>1bt� ���K���� (�:����{O���� ��ʏ܏�uO�$�6� H�Z�l���������Ɵ ؟����� �2�D�V� h�z�	�����¯ԯ� �����.�@�R�d�v� �������п���� ��*�<�N�`�rτ��O �Ϻ�Io��������� 8�J�-�n߀�cߤ߇� ���߽����o1�o X��o|�������� �����0�B�T�f� �������������S� e�w�,>Pbt� �'���� �:L^p��# ���� //$/� H/Z/l/~/�/�/1/�/ �/�/�/? ?�/D?V? h?z?�?�?�???�?�? �?
OO.O��ROdO�� �OkO�O�O�O�O�O�O _�O<_N_1_r_�_g_��_7OM�m�$�UI_QUICK�MEN  ���_AobR�ESTORE 1��  �|��Rto�o�im�o�o�o�o �o:L^p�%� �����o��� �Z�l�~�����E�Ə ؏���� �ÏD�V� h�z���7�������/� ��
��.�@��d�v� ������O�Я���� �ßͯ7�I���m��� ����̿޿����&� 8�J��nπϒϤ϶� a�������Y�"�4�F� X�j�ߎߠ߲����� �ߋ���0�B�T�goSCRE`?#mu1sco`Wu2��3��4��U5��6��7��8��bUSERq�v��Tp���ks����4���5��6��7��8���`NDO_CFoG �#k  n`� `PDATE� ���N�onebSEUFRAME  �T�A�n�RTOL_�ABRTy�l��E�NB����GRP �1�ci/aCz  A�����Q�� $6HRd���`U�����MSKG  �����Nv�%�U�%���b�VISCAND_wMAX�I���FAIL_IM)G� �PݗP#���IMREGNUMr�
,[SIZ��n`�A�,VO�NTMOU���@���2��a���a�����FR:\ �� MC:\ޚ\LOG�B@F� !�'/!+/�O/�Uz M�CV�8#UD1&r&EX{+�S�P�PO64_��0n'fn6PO��CLIb�*�#V����,f@�'�/� �=	�(SZV�.�;���'WAI�/STAT ���B�P@/�?�?�:$�?��?��2DWP  ��P G@+b=��� H�O�_JMPERRw 1�#k
  ��2345678901dF�ψO{O�O�O �O�O�O_�O*__N_�A_S_�_
� MLO�Wc>
 �_TI�=�'MPH?ASE  ��F���PSHIFT֗1 9�]@< �\�Do�U#oIo�oYo ko�o�o�o�o�o�o�o 6lCU�y ����� ��	��V�-�e2����	�VSFT1�2	uVM�� �5�1�G� ���%A� W B8̀̀�@ pكӁ˂�у��z�#ME@�?�{��!�c>&%�aM1��k�0�{ �$`0T?DINEND���\�O� �z����Sp��w��P���ϜRELE�Q��Y����\�_ACTIV���:�R�A �`�e���e�:�RD� ����YBOX ��9�د�6��02����190�.0.�83���254��QF�	 �X�j��1��robo�t���   �p�૿�5pc��̿�����7���x��-�f�ZABC�����,]@U��2ʿ� eϢωϛϭϿ�����  ���V�=�z�a�s�$��E�Z��1�Ѧ