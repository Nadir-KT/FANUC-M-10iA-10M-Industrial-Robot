��   �A��*SYST�EM*��V7.5�0122 8/�1/2   A ����$$CLA�SS  ����(��D��D V?IRTUAL%7�MNUFRAME� AFD�� � 	 88�?��� }��y����� �1=gQs ������	/��/?/��WNUM � ��>lq on�tWTOOLa4 
wY/�/5/�/ �/�/?5??A?k?U? w?�?�?�?�?�?�?O �?	OCO-O?OaOcOuO��O�Om&�!{&���'�