��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  ��'�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"�SBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�� W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2F�G1_�3�B�2	��XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1� ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�0@� �zsa�!ip;G0� � 
$WARNM�0f�!,P� ܁s�pNST� CO�RN�"a1FLTR^�uTRAT� T�p; H0ACCa1�p��{�ORI
`l"S={RT0_S�BְqHG,I1 E[ Tp�"3I9�CTY�D,P*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7���8��94�qO�$ <� $6x8K3 1w`O_M�@�C_ t � E#f6NGP�ABA�  �c��ZQ���`���@n!r��� ��P�0��,��x�p�PzP�b26����"J�_)R��BC�J��3�JVP��tBS��}�Aw��"�tP_*0O�FSzR @� RcO_K8���aIT�3���NOM_�0�1�ĥ3�ACPTC �� $���AxP��K}EX�� �0g0I0x1��p�
$TFa�ކC$MD3��TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF�vF��40CPp@�a2 6
P$A`PU�3N�)#�dR*�AqX�!sDETAI�3�BUFV��p@1c |�p۶�pPIdT�� PP[�MZ�M�g�Ͱj�F[�SIMQSI�"0��A.���9
��lw Tp|z�M��P�B�FAC5TrbHPEW7�P1�Ӡ��v��MCd�k �$*1JB�p<�*1DECHښ�H���(�c� � ~+PNS_EMP��G$GP���,P_���3�p�@Pܤ��TC ��|r��0�s��b�0��� �B���!
���JR|� ��SEGFR���Iv �aR�TkpN&S,�PVF4��� &k�Bv�u �cu��aE�� !2��+�8MQ��E�SIZ�3�����T��P�����aRSINF����Ӏkq��������LpX�����F�CRCMu�3CClpG��p��� O}���b�1�������T2�V�DxIC��C����r����P��{� E�V �zF_��FR�pNB0�?���8���A�! �r� Rx����V�lp�2��a�R�t�,�g�RTx #�5�5"2���uAR���`CX�$LG�p��B�1 `s�P�t�aA�0{�У+01R���tME�`!B�upCrRA 3tA�Z�л�pc�OT�FC�b�`�`FNp���1��ADI+�a% ��b�{��p$�pSp��c�`S�P��a,QMIP6�`Y�3��M'ұpU��aU  ]$>�TITO1�S��S�!��$�"0�DBOPXWO��!��$SK��2�P� d�"�"@�PR8� 
� ���#� >�q1$��)$��+�L9$?(ӤV�%@?R4C&�_?R4ENE��1'~?(�� RE�pY2�(H �OSn��#$L�3$$3�R��;3�MVOk_9D@!V�ROScrr��w�S���CRIGGER2FPA�S��7�ETURN0B�cM[R_��TUː[��0EWM%���G1N>`��RLA���E�ݡ�P�&$PD�t�'�@4a��C�DϣV�DXQ��4�1���MVGO_AWAY�RMO#�aw!��DCS_)  `IS#� ��� �s3S�AQ汯  4Rx�ZSW�AQ�p�@1U9W��cTNTV)�5RV
a���|c�éWƃ¤�JB��x0��SAsFEۥ�V_SV�b�EXCLUU�;�N�ONL��cYg��~az�OT�a{�HI�_V? ��R, M�_G *�0� ��_z��2� CdSGO  +�rƐm@�A@�c~b���w@��V�i|�b�fANNUNx0,�$�dIDY�UABc�@Sp�i�a+ �j�f��!�pOGIx2,���$F�b�$ѐO�T�@A $DUMMY��Ft��Ft�±� 6U- ` !�HE�|s���~bc�B@ SUFFmI��4PCA�UGs5Cw6CrZ� wMSWU. 8!��KEYI��5�TM`�1�s�qoA�vINޱpE��!, / D��oHOST�P!4� ��<���<�°<��p<��EM'���Z�� SB�L� UL��0 � �	����D�T�01 � �$��9USAMPL�о�/���決�$ I�@갯 $SUB ӄ��w0QS�����#��SAV�����c�S�< 9�`�fP$�0E�!� YN_B�#2� 0�`DI�d�pO�|�m��#$F�R_�IC� �ENC�2_Sd3  ��< 3�9���� cgp����4�"��2�rA��ޖ5�� �`ǻ�@Q@K&D-!<�a�AVER�q�����DSP
���PC_�q��"�|�ܣ�oVALU3�HE��(�M�IP)���OkPPm �THЈ*��S" T�/�F�b�;�d����d D���'��ET6� H(rLL_DU ǀ�a�@��k���֠OT�"U�/��o�@@�NOAUTO7�0�$}�x�~�@sT��|�C� ��C� �2iaz�L�� _8H *��L�  ���Բ@sv��`� ��  ÿ���Xq��cq���q����q��7��8��9R��0���1�1 �U1-�1:�1G�1T�U1a�1n�2|�2˪�2 �2-�2:�2�G�2T�2a�2n�3J|�3�3� �3-�U3:�3G�3T�3a�3n�4|�w�����9 <���z�Γ�KI����H硵BaFqEq@{@: ,���&a? P_P?Q��>�����E�@���iaQQ��;fp�$TP�$VA�RI����,�UP2fQ`< W�߃TD�� g���`������q��wBAC�"= T2����$)�,+r³�p IFI��p�� q M�P"�Fl@``>t ;��6����ST����T ��M ����0	��i� ��F���������kRt �����FORCEUyP�b܂FLUS
p�H(N��� ��6bD_CM�@E�7N�� (�v�P��REM� Fa��@j����
K�	N���EcFF/���@IN�Q�OV��OVA��	TROV DyT)��DTMX: e �P:/��Pq�XvXpCLN _�p���@ ��	_|��_QT: �|�&PA�Q	DI���1���0�Y0RQm�_�+qH���M���CL�d#�RIV{�ϓN"�EAR/�IO�P�CP��BR��C�M�@N 1b 3GgCLF��!DY�(ء�a�#5T�DG����� �%��FS9S� )�? P(q1�1�`_1"81�1�EC13D;5�D6�GRA���@������PW�ON<2EBUG�S�2�C`gϐ_E �A ��o� ��TERM�5B�6� �ORIw�0C>�7 �SM_-`����0D�5�qTA�9E~�5�J�UP���F� -Qϒ�A�P�3�@B$SE�GGJ� EL�UUS]EPNFI��pB�x��1@��4>DC$U9F�P��$���QD�@C���G�0T��ܘ��SNSTj�PA�Tۡg��APTHJ�A�E*�Z%qB\`F� {E��F�q�pARxPY�aSHFT͢qA�A>X_SHOR$�>�J�6 @$GqPE���OVR���aZPI�@P@$U?r *aAY#LO���j�I�"�p�Aؠ��ؠERV� �Qi�[Y)��G�@R��Pi�e��i�R�!P�u�ASYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U���C�%UP���P���WO�R�@M��k0SkMT��G��GR��3�aPA�@��p5��'�H � j�NA�TOCjA7pP]Pp$OPd�O��(C�%�p�O!��KRE.pR�C�AO�,?��Be5pR�Eru�Ix'QG�e$PWRf) IMdu�RR_$s���5��B Iz2H|8�=�_ADDRH�?H_LENG�B�q��q:�x�R��So�J6.�SS��SK���`��� ��-�SE*ڕ��0HSN�MN1K	�j�5�@r�֣OL��\�WpW�<Q�>pACRO�p�� �@H ����Q� ��OUPW3�b_>�I��!q�a1������ ��|��������-����:���iIOX2S�=�D�e��]����L $��p�!_O�FF[r_�PRM_����HTTP_��H��M (�pOcBJ�"�pG�$H��LE�C��ٰN � 9�*�AB_�T��
�S�`�S��LV��KRW"duH�ITCOU?BGi�LO�q����`d� Fpk�GpSS� ����HWh�wA��O�.��`INCPU>X2VISIO��!���¢.�á<�á-� ��IOLN)�P �87�R'�[p$S�L�bd PUT_&��$dp�Pz ��� F_AS2Q/�$LD���D�aQ"T U�0]P�A�������PHYG灱Z��Ͱ5�UO� 3R `F���H�Yq�Yx�ɱvpP�Sdp���x�X�ٶ%�UJ��S��v��NE�WJOG�GN �DIS��&�KĠL��3T |��AV���`_�CTR!S^�FgLAGf2&�LG�d�U �n�:��3LG_SIZ��Ű���=���FD��I ����Z �ǳ��0�Ʋ� @s��-ֈ�-�=�-����-��0-�ISCH_H��Dq��N?���V��EE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�B�OO)�WL ?`�� ITV���0\�wREC�SCRf �0�a�D^�����MARG��`!P�)�T�/tHy�?I�S�H�WW�I���T�JGM��M�NCH��I�FNK�EY��K��PRG���UF��P��FW�D��HL�STP���V��@�����RESS�H�` �Q�C�T@1�ZbT�R ���U������|R��t�i���G��8PPO��6�F�1�M��FOCU��RwGEXP�TUI��	IЈ�c��n�� n����ePf���!p6��eP7�N���CANAxI�jB��VAIL���CLt!;eDCS_CHI�4�.��O�D|!�S Sxn瘱I�BUFF1�XY��PT�$ �� �v��f�L6q
1YY��P ������pOS1�2�3���_�0Z �  ��aiE�*���IDX�dP�RhrO��+��A&ST��R���Yz�<! Y$EK&CK+���Z&pm&KF�1[ L�� o�0��]PL�6pwq�t�^����w��7�_ \ �`��瀰�7�t�#�0C��] ���CLDP��;eTRQLI�jd.�094FLGz�0r1R3�1DM�R7��LDR5<4R5ORG.���e2(`@���V�8.��T<�3�d^ �q�<4��-4
R5S�`T00m��0D}FRCLMC!D`�?�?3I@��MIC���d_ d���RQzm�q�DSTB	��  �Fg�HAX�;b �H�LEXC#ESZr��rBMup�a%`� �B;doE`�j�`a��F_A�J���$[�O�H0K�db� \��ӂS�$MB既LIБ}SREQUIR�R>q�\Á�XODEBU��oAL� MP�c�ba��P؃ӂ!B�MND���`�`ad�҆�c�cDC1��IN�����`@�(h�?Nz�@q��o�L��TPST8� en�rLOC�RI�p�EX�fA�p��A�oAODAQP�f �X��ON��[rMF �����f)�"I��%�e؃�T��!FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y��RFЭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?
�uD�)�b�	@Ð�i �@CU��V��T0�eRR2�j� Dɐ�Qނ�Bd$OCALI�@F�G�:s�2�RIN��v��<��NTE���k�E���,��b����_Nl��ڂ��kDׄR�m�DIViFDH��@ـn�$V؀�'c!$��$AZ�����~�[���oH �$B�ELTb��!ACC�EL+��ҡ��ICRC�t����T/!���$PS�@#2L  �Ė83������<� ��PATH����D����3̒Vp�A_� Q�.�4�B�Cᐈ��_MGh�$DDxQ���G�$FWh���p��m�����b�DE���PPABNԗR?OTSPEED����00J�Я8��@��~̐$USE_�2�P��s�SY��c�ZA kqYNu@Ag���OFF�q�MO�UN�NGg�K�OL�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I̒��4�\B�ݠVEO�w�Ͳ23�_UPE�߳LOWL���00����D���BwP��� �1RyCʀƶMOSIV��JRMO���@GPE�RCH  �OV ��^��i�<!�ZD <!�c��d@�P��!V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�̒�<�1Ӣ`0 ��RTI$Qx�0 MO���МB@ R�0J��D��s�H�x���b�DUM2(��S_BCKLSH_C̒��>�=�q�#��U��ԑ���2�t�]ACLALvŲ�1n�PN�CHK00'%SD�RTY4�k��y�1r�q_6#2�_UM$Prj�Cw�_�SCL���ƠLMT_J1_�LO��@���q��E������๕�幘S�PC��7������P	Co���H� �PU�m�C/@�"XT_�c�C�N_��N��e���S	Fu���V�&#�����9�̒��=�C�u�SH6#��c����1�Ѩ��o�0�͑
��_�PALt�h�_Ps�W�_10���4�R�01D�VG�Jb� L�@J�OGW����TORQU��ON*�Mٙ�sRHљ�&�_W��-�_=��PC��I��I�I�%II�F�`�JLA.,�1[�VC��0�D�B�O1U�@i�B\J�RKU��	@DBOL_SMd�BM%`�_DLC�BGRV���C��I��H_p� �*COS+\�(LN�7+X>$ C�9)I�9)u*c,)b�Z2 HƺMY@!̳( "TH&-�)TH�ET0�NK23�I��"=�A CB6CB=�C�A�B(261C�616SBC�T25'GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t���B�6���AQ|r�f$NE�DpIB U�\B$5��$!��!A�%Ep(G%(!LPH$U�2׵�2SXpCc%pC�r%�2�&�C�J�&!�V�AHV6H3�YLVhJV�uKV�KV�KV�KV
�KV�IHAHZF`RXM���wXuKH�KH�KH��KH�KH�IO2LORAHO�YWNOhJOuKUO�KO�KO�KO�KO�&F�2#1ic%�d�4GSPBALANgCE_�!�cLEk0H_�%SP��T&�b�c&�br&PFULC��hr�grr%Ċ1k�y�UTO_?�jTg1T2Cy��2N&� v�ϰctw�g�p�0Ӓ~���T��O���� �INSEGv�!�R�EV�v!���DIF���1l�w�1m�
�OB�q
����M�Iϰ1��LCHW3AR����AB&u�?$MECH,1� X:�@�U�AX:�P��pY�G$�8pn 
Z���|���ROBR�C�R̒��N��'��MSK_�`f�p WP Np_��R����΄ݡ�1��ҰТ`΀ϳ��΀"�IN�q��MTCOM_�C@j�q  �L��p��$NOR�E³5���$�r� 8� GR�E�S�D�0ABF�$XYZ_DA5A���DEBU�qI��Q��s �`$�COD��� ��k�F��f�$BUFIN�DXР  ��M{OR��t $-�U��)��r�B��Ӱ�����Gؒu � $SIMULT ৐~�� ���OBJ�E�` �ADJUS<>�1�AY_Ik���D_����C�_FIF�=�T� ��Ұ ��{��p� �����p�@:��D�FRI��ӥMT��RO� ��E�z��͐OPWO��ŀv0��SYS�BU�@ʐ$SOP�����#�U"��pPgRUN�I�PA��DH�D����_OUb�=��qn�$}�/IMAG��ˀ�0�P�qIM����IN��q���RGOVR!Dȡ:���|�P~���Р�0L_6p���i⦄�RB���0��ML���EDѐF� ��%N`M*����̰�SL�`ŀw x �$OVSL�vS;DI��DEXm�g� e�9w�����V� ~�N���w����Ûǖ���M�
͐�q<�>�� x HˁE�^F�ATUS����C�0àǒ��BTMT����If���4����(�ŀy DˀEz�g���PE�r����8�
���EXE��V���E�Y�$Ժ ŀz �@ˁ��UP{�h�$�p��XN���9x�H� �PG"��{ h $SUB��c�@_��01\�_MPWAI��P��&��LO��<�F�p��$RCVFAI�L_C�f�BWD�"�F���DEFSP>up | Lˀ`��D�� U�UNI��S���R`���_L�pP��̐���ā}��� B�~���|�t�`ҲN�`KET��Jy���P� $�~��=�0SIZE���h��{���S<�OR��?FORMAT/p 㰷 F���rEMR���y�UX���@�P�LI7�ā  �$�P_SWI���Ş_PL7�A�L_ �ސR�AR��B�(0C��Df��$Eh����C�_=�U� � �� ���~�J3x�0����TIA4��u5��6��MOM��@���� �B��AD��*��* PU70NRW��W� Q����� A$PI�6���	�� )�4l�}69���Q���c�SPEED�PGq�7�D�>D� ���>tMt[��SAM�`痰8>��MOV���$���p�5��5�D�1�$2�������d{�Hip�IN?, {�F(b+=$�H*�(x_$�+�+GAMM�f|�1{�$GET���ĐH�D����
^pL�IBR�ѝI��$HI��_��Ȑ*B6�E��*8A$>G086LW=e6\<G9�686���R��ٰV��$PDCK�Q�H�_����;"��z�.%�7�4*�9� ��$IM_SRO�D�s"���H�"�LE�O�0\H���6@����U� �ŀ��P�qUR_SC�R�ӚAZ��S_SAVE_D�E��NO��CgA�Ҷ��@ �$����I��	�I�  %Z[� ��RX" �� m���"�q�'"� 8�Hӱt�W�UpS(���Q�M��O㵐 .'}q��Cg���@ʣȳ���S�M�AÂ� ?� $PY��g$WH`'�NGp� ��H`��Fb��Fb��Fb��PLM���	� 0h�H�{�X��O��z�Zp�eT�M���� pS��C��O__0_�B_�a��_%�� | S����@	�v��v  �@���w�v��EM��%G R�fr�B�ː���ftP��PMv��QU� �U�qQ��Af�QTH=��HOL��QHYSf�ES�,�UE�t�B��O#��  -�P0�|�gAQ���ʠu�%��O��ŀ�ɂv�p-�A;ӝROG��a2D�E�Âv�_��ĀZ�INFO&���+����bȜ�OI�킍 ((@SLEQ/�#������$o���S`c0O�0�j01EZ0NUe��_�AUT�Ab�CO�PY��Ѓ�{��@M��N�����1�P�
�M ��RGI�����3X_�Pl�$�����`�W��P��j@��G���EXT_CYCtb���p�����h�_NA�1!$�\�<�RO�`]�?� � m���POR�ㅣ���S�RVt�)����DI �T_l���Ѥ{�ۧP��ۧ �ۧ5٩6٩%7٩8���AS�B�-���$�F6����PL�A�A^�TAR��@E `�Z������<��d� ,(@F1Lq`h��@YNL����M�C���PWR�Ѝ�쐔e�DELiAѰ�Y�pAD#q}X�QSKIP��� ĕ�x�O�`NeT!� ��P_x� ��ǚ@�b�p1�1� 1Ǹ�?� �?��>�@�>�&�>�3�>�9��J2R;쐖 m4��EX� TQ�� ��ށ�Q���[�KF�ܴ��@RDCIf� )�U`�X}�R�#%�M!*�0�)��$RGE7AR_0IO�TJB�FLG�igpER�a��TC݃������2�TH2N��� S1�b��Gq T�0' ����M���`qIb���qREF��1�� l�h��E�NAB��lcTPE ?@���!(ᭀ��� �Q�#�~�+2 H�W�
��2�Қ���"�4�PF�X��P��3�қ{�@��������j�4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:L��7�ҟo@�����j�8�����"4Fj�SMSK������a��E�AX�REoMOTE�������@ "1��Q�IOD�5"%I��P�QRd�9Wi@쐣  �������h�쐤��Y"$�DSB_SIGN�4A�Qi�̰C��>%S�232%�Sb�iDEVICEUS#|�R�RPARIT򱾈!OPBIT�Q���OWCONTR`��Qⱓ�RCU� �M�SUXTASK��3NB��0�$TAT-U�P��S@@쐩�F�6�_�PC}��$FREEFRO�MS]p�ai�GET\N@S�UPDl�ARB��SP%0����� !m$USAࢰ�az9�L�ERI��0f��pRY�5~"_ľ@f�P�1�!�6WR	K��D9�F9Х?FRIEND�Q4b�UF��&�A@TOO�LHFMY5�$L�ENGTH_VT��FIR�pqC�@�yE� IUFIN�R:���RGI�1�OAITI:�xGX�l�I�FG2�7G1a�0���3�B�GPRR�DA���O_� o0e�I1R�ER�đ�3&���TCp���AQJVE�G|�.2���F��1�!d� 9Z�8+5K�+5��E�y�|L0�4�X �0*m�LN�T�3Hz��8P9��%�4�3G��W�0�W�RdD�Z��T�ܳ��K�a3d��$cV 2���1��RI1H�02K2sk3K3Jci�aI�i��a�L��SL��R$V�ؠ�BV�EVk��A (bQ*R��� �,6Lc ���9V2F{/P:B��kPS_�Et�$rr8�C�ѳ$A0��wCPR���v�U�cSk��� {�tЇ4��� 0���VX`�!�tX`A��0P�Ё�
�5�SK!� �-qRH��!0���z�NJ SAX�!h�A�@LlA���A�THIC�1p�������1TFE��|�q>�IF_CH�3�A�I0�����G1@�x������9�Ɇ7_JF҇PR(����RVAT��� �-p��7@����D9O�E��COU(���AXIg��OFF{SE+�TRIG�S K��c���Ѽ�e�[�K��Hk���8�IGMA�o0�A-��ҙ�OR?G_UNEV���� �S�쐮d� �$������GgROU��ݓTO2���!ݓDSP��JO1G'��#	�_P'�2�OR���>P6KE�Pl�IR�0�PML�RQ�AP�Q��E�08q�e���SYSG��"v��PG��BRK*Rd�r�3�-��������ߒ<pAD�ݓJ�B�SOC� N�D?UMMY14�p\@�SV�PDE_OP�3SFSPD_O+VR��ٰCO��&"�OR-��N�0.��Fr�.��OV�S!Fc�2�f��F��!�4�S��RA�"LCH�DL�RECOV(��0�W�@M�յF�RO3��_��0� @�ҹ@VE}RE�$OFS�@3CV� 0BWDG�Ѵ`C��2j�
�TR�!���E_FDO>j�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�<#�8$CA�{�|����8$HBK|1,c��IO��.�:!aPPA"�N�3�^��F���:"�DVC_DB�C��d�w"���D�!��1���ç�3��^��ATIO� �q�0�UC�&CAB�BS�PⳍP��䖁�_0c�SUB'CPUq��S�Pa  aá�}0�Sb��c��r"~ơ$HW_C�����:c��IcA�A-�l_$UNIT��l���ATN�f����CY{CLųNECA���[�FLTR_2_�FI���(��}&��L�P&�����_SCT@SF_��F����G����FS|!�¹�CH�AA/����2��RSD�x"ѡb�r�: ;_T��PRO��OÖ� EM�_��8u�q u�q���DI�0e�RAIL�AC��}RMƐLOԠdC��:anq��wq�����PR��SZQ��pfC�ѷ 	��F�UNCŢ�rRIN�kP+a�0 ��!RA� >R 
Я��ίWAR�BLFQ��A������DA�����L�Dm0�aB9��nqBTIvrbؑ��μPRIAQ1�"AFS�P�!�����`(%b���M�I1UÇDF_j@��y1°L�ME�FA�@HRDiY�4��Pn@RS@Q��0"�MULSE�j@f�b�q �hX��ȑ���$.A[$�1$c1Ó~���� x~��EG�pݓ�q!AR����09>B�%AXE��ROB���W�A4�_�-֣S�Y���!6��&S�'W�R���-1���ST�R��5�9�E��C 	5B��=QB90`�@6������OT�0�o 	$�ARY�8�w20���	%�F�I��;�$LINQK�H��1�a_63��5�q�2XY�Z"��;�q�3@��1��2�8{0B�{`D��� CFI���6G��
�{�_J���6��3aOP_dO4Y;5�QTBmAd"�BC
�z�DU"�z66CTURN3��vr�E�1�9�ҍGFL�`���~ �@�5<:y7�� 1�?0%K�Mc�68Cb�8vrb�4�ORQ��X �>8�#op������wq�Uf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W�� �Tυ� ;����QH� !`�ҽ��U�Q�WkeK#�kecXER��	BGE	0��S�dAWa Ǣ:D���7!�!AX�rB!{q��1 uy-!y�pz�@ z�@z6Pz\Pz�  z1v�y�y� +y�;y�Ky�[y��ky�{y��y�q�yD7EBU��$�����L�!º2WG`  A!B!�,��SV���� 
w���m���w� ���1���1���A���A ��6Q��\Q���!�m@���2CLAB3B��U�����S � ÐER���� �� $�@� Aؑ!p�PO��Z�q0zw�_�_MRAȑ_� d  T��-�ERR��T)Yz�B�I�V3@�cNΑTOQ�d:`L� H�d2�]�X�C[!_ � p�`T}0i��_V1�r�a'�4�2-�2<�����@P�����F�$W���g��V_!�l�$�P����c��q"��	V FZN_CFG_!� 4��?º��|�ų����@�ȲW ��'����\$� �n���Ѵ��9c�Q���(�FA�He�,�XEDM�(�����!s��Q�g�P{RV HE�LLĥ� 5�6�B_BAS!�R�SR��ԣo �#S���[��1r�%��2�ݺ3ݺ4ݺ5ݺ6�ݺ7ݺ8ݷ��ROaOI䰝0�0NLK!ưCAB� ��AC-K��IN��T:�1��@�@ z�m�_PUf!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KA1Rӑ�@��RE~��qP��(��QUE������P
��CSTOPI_AL�����0�&���㰑�0SEM�l�b�|�M��d�TYf|�SOK�}�DI������(���_TM>\�MANRQ�ֿ0�E+�|�$KEY?SWITCH&	����HE
�BEAiT����E� LEҒ���U��FO�����O_HOM�On�REF�PPRzP��!&0��C+�OA��ECO��B�r�IOCM�D8׵��]���8�` � DH�1����U��&�MHx�»P�CFORC��f� ���OM�  � @V��|�U,3P� 1-�`� �3-�4��NPXw_ASǢ� 0Ȱ�ADD����$S�IZ��$VAR\ݷ TIP]�\�
2�A򻡐���]�H_� �"S꣩!Cΐ���FRIF⢞�S0�"�c���NF��V ܻ�` � x�`SI��TES�R6SSG%L(T�2P&��AxU�� ) STMTQ2ZPm 6BW�P*�SHOWb��S�V�\$�� ���A00P�a�6���@�J�T�5��	6�	7�	8�	9�	A�	� �!�'��C@�F�0u�	 f0u�	�0u�	�@uP[Pu%121?U1L1Y1f1sU2�	2�	2�	2�	U2�	2�	2�	2U22%222?U2L2Y2f2sU3P)3�	3�	3�	U3�	3�	3�	3U33%323?U3L3Y3f3sU4P)4�	4�	4�	U4�	4�	4�	4U44%424?U4L4Y4f4sU5P)5�	5�	5�	U5�	5�	5�	5U55%525?U5L5Y5f5sU6P)6�	6�	6�	U6�	6�	6�	6U66%626?U6L6Y6f6sU7P)7�	7�	7�	U7�	7�	7�	7U77%727?U7,i7Y7Fi7sv�VP�UPD��  ��|�԰މ�YSLOǢ� � z��и���o��E��`>�^t��АAL1Uץ����CU���w=FOqID_L�ӿu�HI�zI�$FI�LE_���t��$�`�JvSA��� h����E_BLCK��#�C,�D_CPU<�{�<�o����txJr��R ��g
PW O� ��LA��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ���TBCu�C� ��X -$�LE�Ni��v������I���G�LOW_AXMI�F1��t2X�AM����D�
 ��I��s ��}�TOR�D���Dh��� L=���⇒�s���#�_M�A`�ޕ��ޑTCV����T���&���ݡ����J�����J$����Mo���J�Ǜ R�������2��`� v�����F�JK��CVKi�Ρv�Ρ3���J0�ңJJڣJJ�AALң�ڣ���4�5z�&�NA1-�9���␅�L~��_Vj�������� ` �GROU�pD��B�NFL�IC��REQUwIREa�EBUA�0�p����2¯����c�� \^��APPR��C����
�EN�CL9Oe��S_M v��,ɣ�
���� ��MC�&���g�'_MG�q�C� �p{�9���|�BRKz�GNOL��|ĉ R�Ї_LI|��Ǫ�k�J����P
���ڣ��� ��&���/���6��6���8���p���G� ��8�%�W�<2�e�PATHa�z�@p�z�=�vӥ�ϰ�x�CN=�CA�����6p�IN�UC��bqZ��CO�UM��YZ������qE%���2�������PAYLOA��J2L3pR_A	N��<�L��F�B�6��R�{�R_F2LS3HR��|�LOG�������ӎ���ACRL�_u�������.���H��p�$H{���FWLEX
��J�� :�/��� �6�2�����;�M�_�F16����n���������ȟ��Eҟ��� ��,�>�P�b��� d�{������������$5�T��X��v� ��EťmFѯ� ������&�/�A��S�e�+p�x�� �� ������j�4pA�T����n�EL  ��%øJ���ʰJ�E��CTR�Ѭ�T�N��F&��HAN/D_VB[
�pnK�� $F2{�X6� �rSWi��("�U��� $$Mt�h�R��08��@<b 35��^6A�p3�k��qD{9t�A�̈p��A��AA�ˆ0��U���D�˕D��P��G��IS�T��$A��$AN��DYˀ�{�g4�5D��� v�6�v��5缧�^�@��P�����#��,�5�>�(#�� �&0�_�ER!V9�SQA'SYM��] ������x��ݑ���_SH l�������sT�(����(�:�JA���S�c�ir��_VI�#�Oh9�``V_UNI��td�~�J���b�E �b��d��d�f��n�@��������uN���(!�H�������"CqEN� a�D)I��>�Obtr�DpNx�� ��2IxQA�q��q��-��s �p� s����� ��/OMME��r4r�QTVpPT�P ���qe�i����P�x� ��yT�Pj� $DUMMY9��$PS_��RF�q�  ��:� ps���!~q� X�����K�STs�ʰS�BR��M21_V�t�8$SV_ER�t�O��z���CLR�x�A  O�r?p? O�ր � D �$GLOB���#LO��Յ$�o��P�!SYSADR��!?p�pTCHM0 �� ,����W7_NA��/�e���r�SR��l (:]8:m�K6 �^2m�i7m�w9m��9 ���ǳ��ǳ���ŕߝ �9ŕ���i�L�񝀤�m��_�_�_�Tr�XOSCRE�ƀ�� ���STF���}H�pТ6�sq] _v �AŁ� T����TYP�r�K��u�!�u���O�@ISb�!��tsqUE{tG� ����H�S����!RSM_�XuU?NEXCEPWv��CpS_��{ᦵ�ӕ�p��÷���COU ���� 1�O�U�ET�փr���PR�OGM� FLn!7$CU��PO*q���c�I_�pH;� �� 8��N�_HE�
p��Q��pRY ?���,�J�*���;�OUS�� �� @d���$B�UTT��R@���C�OLUM�íu�S�ERVc#=�PAN�Ev Ł� � N�PGEU�!�F��~9�)$HELP��^WRETER��)� ����Q�������@� P�P �IN��s�PNߠw v��1����� ����LN�� �䟀�_��k�$H��M TEX�#�����FLAn +REL�V��D4p�������M��?,��ӛ$�����P=�USR�VIEWŁ� <�d��pU�p0NFyIn i�FOCU��ni�PRILPm+��q��TRIP)��m�UNjp{t� �QP��XuWARN|Wud�SRTOLS��ݕ�����O|SO;RN��RAUư��9T��%��VI|�zu�� $�P�ATHg��CAC�HLOG6�O�LIMybM���'��"��HOST6�!��r1�R�OBOT,5���IMl� D�C� g!��E�L���i��VCPU_AVA�ILB�O�EX7�!BQNL�(���A�� Q���Q ��ƀ��  QpC���@_$TOOL6�$��_JMP� �<I�u$SS�!$>sqVSHIF��|s�P�p�6�s���yR���OSUR=W�pRADIz��2�_�q�h�g! �q�)�LUza$O�UTPUT_BM��IML�oR6(`�)�@TIL<SC	O�@Ce�;��9 ��F��T��a��o��>�3�����w�2�u�P{t��%�D�JU��|#�WA�IT������%�ONE��YBO�ư �� �$@p%�C�SBn)T;PE��NEC��x"p�$t$���*B_T��R��%�qR� ���s	B�%�tM�+��t�.`�F�R!݀��OPm�wMAS�_DOG�OaT	�D����C3�S�	�O2DELAY���e2JO��n8E� �Ss4'#J�aP6%�����Y_��O2$��2����5��`? �sqZABCS�� � $�2��J�
�sp�$$CLAS>�����AB�xsp'@@VIRT��O.@ABS�$�1� <E� < *A tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R��d�v�����M@[�AX�LրK�*B�dC  ����IN��ā��P#RE������LARMRECO�V <I䂥�N�G�� \K	 �A   J�\�M@PoPLIC�?<E��E�Ha�ndlingTo�ol �� 
V�7.50P/28~[�  �P���
�_SW�� �UP*A� ��F�0ڑ����A����� 20��*A��:����[�FB 7DA�5�� '@�P@��No�ne������ ���Twk*A4_	Oxl�_���V����g�UT�OB�ค����HGAPON8@��LA�ѽU��D 1<EfA����������� Q 1שI Ԁ��Ԑ�:��i�n����#B�)B ���\��HE�Z�r�HTTHKY��$BI�[�m� ����	�c�-�?�Q� o�uχϙϫϽ����� ���_�)�;�M�k�q� �ߕߧ߹�������� [�%�7�I�g�m��� �����������W�!� 3�E�c�i�{������� ��������S/A _ew����� ��O+=[a s������� K//'/9/W/]/o/�/ �/�/�/�/�/�/G?? #?5?S?Y?k?}?�?�? �?�?�?�?COOO1O OOUOgOyO�O�O�O�O �O�O?_	__-_K_Q_���(�TO4�s���DO_CLEAN��|e��SNM  9� �9oKo]ooo��o�DSPDRY�R�_%�HI��m@ &o�o�o#5GY k}����"����p�Ն �ǣ�qX�Մ��ߢ��g�PLU�GGҠ�Wߣ��PRUC�`B`9��o��=�OB��oe�SEGF��K������o %o����#�5�m���LAP�oݎ������ ����џ�����+��=�O�a���TOTA�L�.���USENUʀ׫ �X���R�(�RG_STRI�NG 1��
��M��Sc��
��_ITEM1 �  nc��.�@� R�d�v���������п �����*�<�N�`��r�I/O S�IGNAL���Tryout M�ode�Inp���Simulat{ed�Out��OVERR�`� = 100�In cycl����Prog A�bor�����S�tatus�	H�eartbeat���MH FauylB�K�AlerU� ��s߅ߗߩ߻�����8���� �S�� �Q��f�x���� ����������,�>��P�b�t�������,�WOR������V��
 .@Rdv�� �����*8<N`PO��6� ���o����� //'/9/K/]/o/�/ �/�/�/�/�/�/�/�DEV�*0�?Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO��O�O�OPALT B��A���O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:o�OGRI�p��ra�OLo �o�o�o�o�o�o *<N`r��� ���`o��RB�� �o�>�P�b�t����� ����Ώ�����(��:�L�^�p����PREG�N��.������ ��*�<�N�`�r��� ������̯ޯ����&����$ARG_���D ?	����i�� � 	$��	+[}�]}���Ǟ��\�SBN_CON?FIG i��������CII_SAVE  ���۱Ҳ\�TCEL�LSETUP �i�%HOME�_IO�͈�%M�OV_�2�8�RE�P���V�UTOB�ACK
�ƽFRA:\��� �Ϩ���'`� ��������� ����$�6�c�Z�8lߙ��Ĉ������ �������!凞��M� _�q����2����� ����%�7���[�m� �������@�������`!3E$���J�o�������I�NI�@��ε~��MESSAG�����q��ODE_!D$���O,0.ޜ�PAUS�!�~i� ((Ol� ������� / �//$/Z/H/~/l/�/�'akTSK � q�����UP3DT%�d0;�WSM_CF°�i�еU�'1GRgP 2h�93 |��B��A�/S�XSC�RD+11
1; 	����/�?�?�?  OO$O��߳?lO~O �O�O�O�O1O�OUO_  _2_D_V_h_�O	_X�>��GROUN0O��SUP_NAL��h�	�ĠV_ED�� 11;
 �%�-BCKEDT�-�_`�!oEo$����a��o����,�ߨ���e2no_��o�o�b���ee�o"�o�oED3�o��o ~[�5GED4�n#�� ~�j���ED5Z��Ǐ�6� ~���}���ED6����k�ڏ ~G���!�3�ED7��Z���~� ~�V�şןEDa8F�&o��Ů}p����i�{�ED9���W�Ư
}3�����CRo�����3��տ@ϯ����P�PNO�_DEL�_�RGE?_UNUSE�_�T�LAL_OUT �q�c�QWD_ABOR� �΢Q��ITR_RTN�=���NONSe����CAM_PARAM 1�U�3
 8
SO�NY XC-56� 2345678�90�H � �@���?���(O АV�|[r�u�~�X�HR5k�p|U�Q�߿�R57�����Aff��K�OWA SC31�0M|[r�̀�d @6�|V�� _�Xϸ���V��� ����$�6��Z�l��CE�_RIA_I8j57�F�1��tR|]��_LIO4YW=� ��P<~��F<�GP 1�,���_GYk�*C*  ��CU1� 9� @� G� Z�CLC]� d� l� s�R� ��U[�m� v� � }�� �� C�� ő"�|W��7�HEӰONFI� ��<�G_PRI 1�+P�m®/���������'CHK�PAUS�  1E� ,�>/P/:/ t/^/�/�/�/�/�/�/ �/?(??L?6?\?�?"O�����H�1�_MOR�� y�0�5 	 �9  O�?$OOHO6K�2	"���=9"�Q?55I��C�PK�D3P�������a�- 4�O__|Z
�OG_��7�PO�� ��6_��,,xV�ADB���='��)
mc:cpm�idbg�_`��S:_�  ��P�����Up�_)o�S  ?�  A���Ra�P�_mo8j�"�a�Koo�o9i�(�EՓog�o�o�m��o�f�oGq:I�ZDE�F f8��)��R6pbuf.txAtm�]n�@�����# 	`(Ж�A=L����zMC�21B�=��9���4�=��n׾�Cz  B�HBCCo�C|���CqD���C���C��{iSZE@D���F.��F���E⚵F,�E�ٙ�E@F�N��IU��I?O��I<#I6��I�SY����vqG���Em��(�.��(�(���<�q�G�x2���2� �� a�D�j����ES\E@EX��EQ�EJP �F�E�F� �G�ǎ^F �E�� FB� �H,- Ge���H3Y���  �>�33 ����xV  n2xQ@F��5Y��8B� A�A�ST<#�
� ��_'�%��wRSMO�FS���~2�yT}1�0DE �Of@b 
�(�;�"�G  <�6�z�R���?�j�C4��SZm� W��{�m��C��B-G�Cu�@�$�q��T{�FP?ROG %i����c�I��� �Ɯ�f��KEY_TBL � �vM�u� �	
��� !"�#$%&'()*+,-./01c��:;<=>?@A�BC�pGHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������p����͓���������������������������������耇���������������������!j�LCK��.�j����STAT���_AUTO_DO����W/�INDT_'ENB߿2R��9��+�T2w�XSTO�P\߿2TRLl�L�ETE����_S�CREEN ~ikcsc���U��MMENU �1 i  <g\��L�SU+�U�� p3g���������� ��2�	��A�z�Q�c� ��������������. d;M�q� �����N %7]�m�� �/��/J/!/3/ �/W/i/�/�/�/�/�/ �/�/4???j?A?S? y?�?�?�?�?�?�?O �?O-OfO=OOO�OsO �O�O�O�O�O_�O_�P_Sy�_MANU�AL��n�DBCO�U�RIG���DB'NUM�p��<����
�QPXWORK 1!R�ү�_o�O.o@oRk�Q_AW�AY�S��GCP� ��=��df_AL�P�db�RY��������X_�p 1"�� , 
�^���o( xvf`MT�I^�rl�@�:sONTIM6������Zv�i�
õ�cMOTNE�ND���dRECO_RD 1(R�a��ua�O��q�� sb�.�@�R��xZ��� ����ɏۏ폄��� #���G���k�}����� <�ş4��X���1� C���g�֟�������� ӯ�T�	�x�-���Q� c�u����������>� ���)Ϙ�Mϼ�F� ࿕ϧϹ���:����� ��%�s`Pn&�]�o��� ��~ߌ���8�J���� ��5� ��k����ߡ� ��J�����X��|�� C�U�����������0�����	��dbTO�LERENCqdB�Ⱥb`L�͐PC�S_CFG )��k)wdMC:�\O L%04d.'CSV
�Pc�)s[A �CH� z�P�)~���hMR�C_OUT *��[�`+P SGN� +�e�r��#��10-MAY-�20 09:07~*V17-FEBj�1o9�k PQ�8��)~�`�pa�m��P�JPѬVE�RSION �SV2.0.�8.|EFLOGI�C 1,�[ 	DX�P7)�PF."�PROG_ENB��o�rj ULSew ��T�"_WRST�JNEp�V�r`dEM�O_OPT_SL� ?	�es
 ?	R575)s7)��/??*?<?'�$TO  �-��?&[V_@pEX�Wd�u��3PATH ASA\�?�?O�/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C��SqqF�PMAU�� t/XrMSWR.D�i6.|S/�Z!D_N�O0__T_C_�x_g_�_�tSBL_/FAUL"0�[3w/TDIAU 16M6�p�A12�34567890gFP?BoTofo xo�o�o�o�o�o�o�o ,>Pb�S�p-P�_ ���_s �� 0`����� )�;�M�_�q����������ˏݏ��|)UM�P�!� �^�T�R�B�#+�=�PME�fEI�Y_TEMP9 È�3@�3A �v�UNI�.(YN_BRK 2Y�)EMGDI_S�TA�%W!bՐNC�2_SCR 3��1o"�4�F�X�fv ���������#��ޑ14����)�;������ݤ5��� ��x�f	u�ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/߭P�b�t�� �� xߞ߰���������
� �.�@�R�d�v��� �����������*� <�N���r��������� ������&8J \n������ ��"`�FXj |������� //0/B/T/f/x/�/ �/�/�/�/�/�/4? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�O�O ?�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�O�O�o�o�o
 .@Rdv�� �������*� <�N�`�r����o���� ̏ޏ����&�8�J� \�n���������ȟڟ�����H�ETMO�DE 16���� ��ƨ
�R�d�v�נRROR�_PROG %fA�%�:߽�  ���TABLE  �A������#�L�R�RSEV_NUM�  ��Q���K�S���_AUT�O_ENB  ���I�Ϥ_NOh� �7A�{�R� W *���������	���^�+��Ŀֿ���HISO�͡I�}�_ALM 18A�� �;�����+�e�wωϛϭϿ�r�_H���  A����|��4�TCP_VER !A��!����$EXTL�OG_REQ�9�{�V�SIZ_�QԿTOL  ͡D�z��A Q�_BWD����r���n�w_DI�� 9���}�z�͡m���S�TEP����4��O/P_DO���Ѡ�FACTORY_�TUN�dG�EATURE :�����l�Ha�ndlingTo�ol ��  - �CEngli�sh Dicti�onary��OR�DEAA V�is�� Mast�er���96 H���nalog I�/O���H551���uto Sof�tware Up�date  ��J���matic B�ackup��Pa�rt&�gro�und Edit���  8\apCamera��F��t\j6R�e�ll���LOADnR�omm��shq�ޝ�TI" ��co<��
! o����pane�� 
�!��tyle �select��H�59��nD���onoitor��48�����tr��Reli�ab���adin�Diagno�s"����2�2 ua�l Check �Safety UIF lg\a���hanced Rob Serv �q ct\��lU?ser FrU���DIF��Ext.� DIO ��fi�A d��end.r Err L@��KIF�r��  �����90��FCTN_ MenuZ v'���74� TP I�n��fac  SU (G=�}p��k Excn �g�3��High�-Sper Ski.+�  sO�H9 � �mmunic!�oknsg�teur� 4����V�����conn��2��E�N��Incrs�tru���5.f�dKAREL Cmd. L?�uaA� O�Ru�n-Ti� Env�����K� ��+%�sn#�S/W��74��LicenseT��  (Au* o�gBook(Sy���m)��"
�MACROs,~V/Offse��ap��MH� �����pfa5�Mech�Stop Pro�t��� d�b i��Shif���j545�!xr ��#�ޜ�,^b od�e Switch.��m\e�!o4=.�& pro�4���g��Mult�i-T7G��net.Pos �Regi��z�P>��t Fun����3 Rz1��Numx �����9m�1� � Adjuj��1' J7�7�* ����6tatuq1EI�KRDMto}t��scove�� ��@By- }u'est1�$Go� � �U5\SNPX� b"���YA�"Libr����#��1 �$~@h�pd]0��Jts in V�CCM�����0� 8 �u!��2 R�0��/I�08��TM�ILIB�M J9u2�@P�Acc>��F�97�TPTXl�+�BRSQelZ0�M8 Rm��q%���692��Unex�ceptr mot}nT  CVV�P���KC����+-|��~K  II)�VSP CSXC�&�.c�� e�"�� t��@Wew�A3D Q�8bvr ngmen�@�iP� �a0y�0�pfGr�idAplay �!� nh�@*�3R�1M�-10iA(B2�01 �`2V"  �F���scii�l�oad��83 M��l����Guar��d J85�0�mP�'�L`���stuaPsat�&]$Cyc���|0ori_ x%D7ata'Pqu����ch�1��g`� j6� RLJam�5��|��IMI De-By(\A�cP" #^0�C  etkc>^0asswo%q�)650�ApU�Xsnt��Pven�C�TqH�5�0Y�ELLOW BO�?Y��� Arc�0v�is��Ch�We{ldQcial4Izt�Op� ��gs֛` 2@�a��pofG yRjT1 �NE�#HT� xy�Wb��! �p�`g�d`���p\� =P��JPN ARCP*�PR�A�� O�L�pSup̂fi�l�p��J�� ��cro�670�1C~E�d���SS�pe�teex�$ �P� So7 �t� ssagN5 D<Q�BP:� �9 "0F�QrtQC��P�l0dpn�笔�rpf��q�e�ppma�scbin4ps{yn�' ptx]0�8�HELNCL� VIS PKGsS �Z@MB �&��B J8@IP�E GET_VA�R FI?S (U�ni� LU�OOL�: ADD�@29�.FD�TCm���E�@DVp���`A�Т�NO WTWTE'ST �� &�!���c�FOR ��EC�T �a!� ALS�E ALA`�CP?MO-130��� �b D: HANG FROMg��2���R709 DR�AM AVAIL�CHECKS 5�49��m�VPCS� SU֐LIMC�HK��P�0x�FF� POS� F�� �q8-12 oCHARS�ER6��OGRA ��Z@A�VEH�AME��.#SV��Вאn$���9�m "y�TRC�v� SHADP�U_PDAT k�0���STATI��� �MUCH ���T�IMQ MOTN�-003��@O�BOGUIDE DAUGH���b��@$tou� �@C�y �0��PATH�_�MOVET�� �R64��VMXP�ACK MAY ?ASSERTjS��oCYCL`�TA���BE COR 7�1�1-�AN��RC� OPTIONS�  �`��APSH;-1�`fix��2�SO��B��XO򝡞�C_T��	�i��0j���du�byz p w1a��y�٠HI�����U�pb XSPD� TB/�F� \h�chΤB0���EN�D�CE�06\Q�p�{ smay n�@�pk��L ��tOraff#�	� ���~1from s�ysvar sc�r�0R� ��d�DJ�U���H�!A��/���SET ERR��D�P7����ND�ANT SCRE�EN UNREAO VM �PD�D���PA���R�IO� JNN�0�FI���B��GROUNנD Y�Т٠��h�SVIP 53� QS��DIGIT VERS��ká��NEW�� P06z�@C�1IMAG�hͱ���8� DI`<���pSSUE�5���EPLAN JO�N� DEL���15�7QאD��CAL�LI���Q��m���I�PND}�IMG oN9 PZ�19���MNT/��ES ܏��`LocR Ho�l߀=��2�Pn� P�G:��=�M��ca�n����С: 3�D mE2view� d X��eat1 �0b�pof Ǡ�"HCɰ�ANN�OT ACCESS M cpie�$Et.Qs a� l�oMdFlex)a:z��w$qmo G�s�A9�-'p~0��h0p�a��eJ AUTcO-�0��!ipu@�Т<ᡠIABLE�+� 7�a FPLNs: L�pl m6� MD<�VI�и�WIT HOC�;Jo~1Qui��":��N��USB�@�P�t & remo�v���D�vAxisO FT_7�PGɰ�CP:�OS-1�44 � h s s268QՐOST�p�  CRASH �DU��$P��WO�RD.$�LOG3IN�P��P:	�0��046 issu�eE�H�: Sl�ow st�cB�`6����໰IF��IMPR��SPO�T:Wh4���N1S�TY��0VMGR��b�N�CAT��4�oRRE�� � �58�1��:%�RT�U!Pe -M a�SE�:�@pp���AGpL���m@allء�*0a�OCB W�A���"3 CNTw0 T9DWroO0alarm�ˀm0d t�M�"0�2|�s o�Z@OME<�x� ��E%  #1-�gSRE��M�st}0g     5�KANJI5no� MNS@�IN�ISITALIZf'� E�f�we���6@� dr�@ fp� "��SCII �L�afails �w��SYSTE0[�i��  � Mq��1QGro8�m n�@vA����&���n�0q��RWRI� OF Lk��� �\ref"�
�up�� de-rela��Qd 03.�0S�Schőbetw�e4�IND exm ɰTPa�DO� �l� �ɰGig�E�soperab�il`p l,��H0cB��@]�le�Q0cflxz�Ð���OS {����v4pf;igi GLA�$��c2�7H� lapn�0ASB� If��=g�2 l\c�0���/�E�� EXCE 㰁�P���i�� o0��Gd`]Ц�yfq�l lxt��EFal��#0�i�xO�Y�n�CLOS��SRNq1NT^�F��U��FqKP�ANIOO V7/ॠ1�{8����DB �0���ᴥ�ED��DET�|�'� �bF�NLwINEb�BUG�Tt���C"RLIB���A��ABC JA�RKY@��� rk�ey�`IL���PRr��N��ITGAR� D$�R �Er *�T��a�U�0��h��[�ZE V� T�ASK p.vr��P2" .�XfJ�s�rn�S谥dIBP�	c���B/��BU]S��UNN� j0�-�{��cR'���L�OE�DIVS�CU�Ls$cb����BW !��R~�W`P�����IT(঱tʠ�O=F��UNEXڠ+�Ҧ�p�FtE��SV�EMG3`NML �505� D*�CC_SAFE�P*� �8ꐺ� PET��'P��`�F  !���IQR����c i S>�� K��K�H G_UNCHG��S�/MECH��M���T*�%p6u��tPORY LEAK�9J���SPEgD���2V 74\GR�I��Q�g��CTLN��TRe @�_�p l���EN'�IN�������$���r��T3\)�i�STO�A�s�L��͐X	���qb��Y� ��TO2�J m��0F<�K����SDU�S��O��3 9�J F�&��~�SSVGN-1#�I���RSRwQDAU��Cޱ� �T6�g��� �3�]���BRKCTqR/"� �q\j5�p�_�Q�S�qINVJ0D ZO�Pݲ���s ��г�Ui ɰ̒�a��DUAL� J5�0e�x�RVO117 AW�TH!Hr�%�N�247%�528��|�&aol ���RP���at�Sd�cU���P,�LER��iԗQ<0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�c�豓�{�U��ROP� 2�b�pB��IT�P4M��b !A�Ut c0< � pleste�N@� z1�^qR635 (AccuCal2kA=���I) "�ǰ�1a\�Ps��ǐ� �bЧ0P򶲊���i�g\cbacul "A3p_ �1��ն|���etaca��AT���PC�`����v�_p�.pc!�x���:�circB���5�tl��Bɵ�:�Cfm+�Ί�V�b�����r�upfrm.0����ⴊ�xed��Μ��~�pedA�D �|}b�ptlibB�� �_�rt��	��_\׊ۊ�6�fm �݊�oޢ�e��̆Ϙ�"��c�Ӳ�5�j>���F��tcȐ��	�r�����mm 1��T�sl^0��T�mѡ�#�rm3��ub Y�q�gstd}��pl;��&�ckv�=�r�vf0�䊰��9�vi�����ul�`�0fp�q ��.f��� da�q; i Data Acquisi���n�
��T`��1�89��22 �DMCM RRS�2Z�75��9 3� R710�o5�9p5\?��T ="��1 (D�T� nk@��������E �Ƒȵ��Ӹ�etdmm ��ER�����gE��1�q\mo ?۳�=(G���`[(

�2�` ! �|@JMACRO���Skip/OffCse:�a��V�4oy9� &qR662�H��s�H�
 6Bq�8����9Z�43� J77� 6�J783�o ��n��"v�R5IKC~Bq2 PTLC�vZg R�3 (�s, ��������03�	зJԷ\s�fmnmc "M�NMC����ҹ�%m;nf�FMC"Ѻ|0ª etmcr� ��8���� �,^D&^�   874\Oprdq>,jF0����axisHP�rocess A�xes e�rol�^PRA
�Dp� 5�6 J81j�59� 56o6� ���06w�690 98� [!GIDV�1��2(x2��2ont�0�
� ���m2���?C���etis "IS�D��9�� FpraxRAM�P� D�чdefB�,�G�i�sbasicHB��@޲{6�� 708*�6��(�Acw:� �����D
�/,��AMOX�� ��DvE��?;Td��>Pi� RAFM';�]�!PAM�V�W�E�e�U�Q'
bU�75��.�ceNe� nterface^4�1' 5&!54�K��b(Devam±�/@�#���/<�Tane`�"DNEWE���bt�pdnui �AI��_s2�d_rso!no���bAsfjN�>�bdv_arFvf�`xhpz�}w��hkH�9xstc��gApocnlGzv{�ff� �r���z�3{q�'Td>pcham�pr;e�p� ^59�77��	܀�4}0��m�Ɂ�/�����lf�!�p�cchmp]aMP�&B�� �mpevp�����pcs���YeS�� Macr%o�OD��16Q!)* �:$�2U"_,��Y�(PC ��$_;������o��J�gege=mQ@GEMSW�~Z>G�gesndy��OD�ndda��S��csyT�Kɓ�su^҈����n�m���L�� ' ���9:p'ѳ�޲��spotplusp���`-�W�l��J�s��t[�׷p�key�ɰ�$��s�-����m���\featu 0FEAWD�woolo�srn'!2 p���a�As3���tT.� (N. A.)��!e!�J# (j�,��oBLIB�oD -�.�n��k9�"K��u[-��_���p� "PS�EqW����wop "sEЅ�&�:�J� �����y�|��O8�� 5��Rɺ���ɰ[��X �������%�(
���q HL�0k�
�z�a!�B�Q�"( g�Q�����]�'�.� ����&���<�!ҝ_�#��tpJ�H�~Z��j� ����y������2�� e������Z����V�� !%���=�]�͂��^2n�@iRV� on�IQYq͋JF0� 8ހȖ`�	(^�dQueue���X\1�ʖ`��+F1tpvtsn���N&��ftpJ0v �RDV�	f��J1� Q���v�en���kvstk��m�p��btkclrqq���get�����r��`ka�ck�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�mc�N+v3�_� �����.v�/\=jF��� �`Q��΋ܒ�N50 (F�RA��+��͢fraparm��Ҁ�z} 6�J643p:~V�ELSE
#��VAR $SGSYSCFG.$�`�_UNITS 2��DG~°@�4Jgfr8��4A�@FRL-��0 ͅ�3ې���L�0NE �:�=�?@�8�v�9�~Qx304��;�BP�RSM~QA�5TX�.$VNUM_O�L��5��DJ507���l� Funct�ʂ"qwAP��琉�3# H�ƞ�kP9jQ�QA5ձ� ��@jLJzB J[�6N�kAP���|�S��"TPPR����QA�prnaS�V�ZS��AS8Dj5150U�-�`cr�`8 ���ʇ�DJR`jYȑH�  �Q ��PJ6�a21��4�8AAVM �5�Q�b0 lB�`T�UP xbJ5�45 `b�`616����0VCAM� 9�CLIOn b1�5 ����`MSC8�
rP �R`\sSTY�L MNIN�`J�628Q  �`N�REd�;@�`SCH� ��9pDCSU �Mete�`ORSsR Ԃ�a04 kREIOC �a]5�`542�b9vp�P<�nP�a�`�R�`7��`�MASKg Ho�.r7 �2��`OCO :��r3@��p�b�p���r0X�|�a�`13\mn�a39 HRM"�q��q��LCHK>�uOPLG B��a�03 �q.�pHC�R Ob�pCpPo�si�`fP6 is�[rJ554�òpDSW�bM�D�pqR�ag37 }Rjr0 �1��s4 �R6�7��5�2�r5 �2�r7 �1� P6���Reg�i�@T�uFRKDM�uSaq%�4�`�930�uSNBA��uSHLB̀\suf"pM�NPI��SPVC�J52�0��TC�`"MN�рTMIL�IF�V�PAC W�pT�PTXp6.%�T�ELN N Me��09m3UEsCK�b�`UFR�`ކ�VCOR��VI�PLpq89qSXC��S�`VVF�J�T�P �q��R626.l�u S�`Gސ�2?IGUI�C���PGSt�\ŀH8�63�S�q�����q3u4sŁ684��0�a�@b>�3 :B��s1 T��96 .��+E�51 y�q5�3�3�b1 ���b1� n�jr9 ���`V�AT ߲�q75 �s�F��`�sAWSM<��`TOP u�ŀ�R52p���a80 �
�ށXY q���0� ,b�`885�QXрOLp}�"pE࠱;tp�`LCMD���ETSS���6 |�V�CPE oZ1��VRCd3
�NL:H�h��001m2Epƌ�3 f��p��4 _/165C��6l�ꌰ7PR��008� tB��9 -20-0�`U0�pF�1޲1 ��޲2L"���p���޲4��5 \�hmp޲6 RBC�F�`ళ�fs�8 ��Ҋ��~�J�7 r'bcfA�L�8\PC����"�32m0u�n��K�Rٰn�5 5E7W
n�9 z��g40 kB��3 ���6ݲ�`00iB/���6�u��7�u��8` µ������sU0�`��t �1 05\rb��2 E���K�Ȇ�j���5˰��60 ��a�HУ`:�63�jA0F�_���F�7 ڱ݀�H�8�eHЋ��cU0$��7�p��1u��y8u��9 73��L����D7� ��5t󮊱97 ��8U�1(��2��1�1:���Eh��1np�"��8(�{U1��\pyl���,࿱v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6 B���цp��1�����1�`͵155�ض157 �2��6A2�S����1b�H�2����1Π"�2��&�B6`�1<c�34 7B�5 DR���8_�B/��187y uJ�8 06��90 rBn�1 (���202 0EWE,ѱ2^��2��90�cU2�p�2��2 b��4��2�a"RB4����9\�U2�`w�<l���4 60Mp��7������b�s
5� ��3����pB"9� 3 ����`ڰR,:7 �2��V�2��5���2^��a^	9���qr����n�A5����5᥁"�8a�$Ɂ}�5B���5���B�`UA���� ��86 V�6 S�0��5�px�2�#�529 �2P^�b1P�5~�A2`���&P5��E8��5��u�!�5���ٵ544��5��R��ąP nB^z�c �(�4�����U)5J�V�5��1�1^���%�����5 b�21��gA��58�W82� rb��5N�E�5890r� 1�95 �"���� ��c8"a��|�L ���!J"5|6��^!�6��B�"8�`#��j+�8%�6B�AME�޶"1 iC��62�2�Bu�6V��d� 4���84�`ANRS�P�e/S� C@�5� �6� ��� \� ��6� �V� 3t��� T20CA�R���8� Hf� 1DH�� �AOE� �� ;,|�� �0\�,� �!64K��ԓrA|� �1 (M-7�!/50T�[PM��P�Th:1�C�#Pe�� �3�0� 5`M7�5T"� �D8p� ��0Gc� u�4��i1-O710i�1� Skd�7j�?6�:-HS,� �RN�@�UB�xf�X�=m75sA*A6an���!/CB�B2.6A �0;A�CIB@�A�2�QF1�UB2�21� /70�S� �4�����Aj1�3p�p��r#0 B2\m*A@C��;bi"i1K�u"�A~AAU� imm7c7��ZA@I�@�D�f�A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A �5*A�EA�5B�4>\77
B7=Q�D�2�Q�$B�E7�C�D/qAHEE�W7�_|`jz@�  2�0�Ejc7�`�E"l7�@7�A
1�EH�V~`�W2%Q�R9�.�@0L_�#����"�A���b��H3s=rA/2�R5nR4�74r�NUQ1ZU�A�s\m9
1M92L2�!F!^Y:�ps� 2ci��-?�qhimQ�t  w043 �C�p2�mQ�r�H_ �H20�Evr�QHsXBSt#62�q`s����� x��Pxq350_*AF3I)�2�d�u0�@�� '4TX�0�pa3i1A3sQ25�c&��st�r�VR1%e�q0
��j1��O2� ���A�UEiy�.�‐ ț0Ch20$CXB79�#A�ᓄM Q1]�~�� 9�Q��?PQ��qA !Pvs� 5	15aU����?PŅ���ဝQ9#A6�zS*�7�qb5��1����Q��00P(��V7]u�aitE1�� �ïp?7� !?�z��{rbUQRB1PM=��Qa9��H��QQ�25L�������Q��@�L��8ܰ��y00�\ry�"R2BL��tN  ���; �1D&^�2�qeR�5���_b�3��X]1m1lcqP1�a�E�Q� 5F����!y5���@M-16Q� � f���r��Q�e� p��� PN�LT_�10��i1��9453��@8�e�|�b1l>F1@u*AY2�
��R8�Q0����RJ�J3�D}T� 85
Qg�/0��*A�!P�*A�Ð𫿽�2,ǿپ6t�6=Q��`�Pȓ��� AQ� g�*ASt]1^u�ajr I�B����~�|I�b�L�yI�\m�Qb�I�u�z�A�c3Apa9q� B6S��S��m���}��85`N�N�  �(M���f1��@�6����161��5�s`�SC��U��A�����5\set06�c����10�y�h8��a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��@���5�B��B��h`� F���X0���A:���C�M��AZ��@��4�6@i����� e�O�-	 ���f1��F �ᱦ��1F�Y	���T6HL3��U66~`���U�9dU�9D20Lf0�� Qv� ��fjq��N�� ����0v
� ��i	�\	��72lqQ2������� \chn?gmove.V���d���@2l_arf	�f~��6� �����9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�AX]��V�1\�Qn�BJ�2W�EM!`5���)�#:�64��F�e50S�\��0 �=�PV���e���逕��E�����mw7shqQSH"U��)��9�!A��(����� ,^9�ॲTR1!��&,�60e=�4F���2��2��	 R-��� ��������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2�"�2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D��� 5V��@2cVE����dT��pt갖�1L~E��#�F�Q��9E�#De1/��RT��59���	��A�EiR������9o\m20�20��+�-u�19r4�`�E1 �=`O9`�1"ae���O�2��_$W}am�41�4�3�/d1c_std��1)Ķ!�`_T��r�_ 4\jdg�a�q�PJ %!~`-�r�+bgB���#c300�Y�5j�QpQb1�bq��vB��v25�U������qm43� �Q<W�" PsA��e��� �t�i�P�W.��c��FX.�e�kE14��44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2-a��2A;_2��QW�2�bF�(�V11�2�3�`��X5�Ra21B�J*9�a:88rJ9X�l5�m1a�0���*���(85�&� ������P6���RB,52&A����,fA�9IfI50\u�z�O@V
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq� &ŦP1��vB)e�m�x����1p� �1�D&^�27�F�K�AREL Use{ S��FCTN��� J97�FA+�� (�Q޵�p%�)?��Vj9F?(�j�Rtk208 "Km�6Q�y�j��iæPr��9�s#��v�krcfp�RCFt3���Q~��kcctme�!�ME�g����6�ma�in�dV�� ��r!u��kDº�c���o�����J�dt�F �»�.vrT�f������E%�!��5�FRjK73B�K���UER��HJ�O  J�� (ڳF���F�q�Y��&T��p�F�z��19�tAkvBr���V�h�9p�E�y�<�k������8;�v���"CT��f ����)�
І��)�V 	�6���!��qFF�� �1q���=�����O�?� $"���$��je���TCP Aut�r~�<520 H5��J53E193��9V��96�!8��9���	 �B574��52��Je�(�� Se %!Y�����u��ma�Pqtool�ԕ�������conre�l�Ftrol Reliable�RrmvCU!��H51������ a551xe"�CNRE�I�c�&��it�l�\sfutst �"UTա��"X�\�u��g@�i�6Q]V0H�B,Eѝ6A� �Q �)C���X��Yf�Iȴ1|6s@6i��T�6IU��vR�d�
$e0%1��2�C58�E6���8�Pv�iV4OFH5�8SOeJ� mvBM6E~O58�I�0�E�# +@�&�F�0���F�P 6a���)/++�</N)0\tr1�����P� ,^ɶ�rma;ski�msk�aA����ky'd�h	A	�P��sDisplay�Im�`v����J8�87 ("A��+He<ůצprds��I�T:���h�0pl�2�R�2��:�Gt�@��PRD�TɈ�r�C�@Fpm��D�Q�Asca��� V<Q&��bVvbrl�eې@��^S��8&5Uf�j8710��yl	��Uq���7 �&�p�p��P^@�P�firmQ����Pp� 2�=bk�6�r�3��6���tppl��PL ���O�p<b�ac�q	� �g1J�U�d�J��gait_9e��Y�&���Q���	�Shap���erationx�0��R67451tj9(`sGen� ms�42-f��r�p�50����2�rsgl�E���p�G���qF�205�p�5S���Ձ�ret�sap�BP�O�\s>� "GCR�ö?� �qngda�G ��V��st2axU�b�Aa]��bad�_|�btputl/��&�e���tplibB_��=�2.����5�Ό�cird�v�sl8p��x�hex��v��re?�Ɵx�key��v�pm��x�u9s$�6�gcr��F�������[�q27j92|�v�ollismq�Sk�9O�ݝ� (Gpl.���t��p!o���29$Fo8��cg7�no@�tptcls` CLS�o�b�\�#km�ai_
�s>�v�o	�t�b���ӿ�E��H��6�1en�u501�[m��u�tia|$calm�aUR��CalMa;teT;R51%�i=1]@-��/V� ��Z��� �fq1�9 "KA9E�L����2m��CLMTq�S#��et �LM3!} �:F�c�nspQ�cӞ��c_moq��� ���c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ����N�ve��C�clm��&Ao# �|$fin�de�0ST�D ter Fi?LANG���R��
��n3��z0gCen���r,�� ����J����� ��� K��Ú�=���_Ӛ����r� "FND�R�� 3��f��tguid�䙃N�."��J�tq�� ��������������J����_@������c��	m��Z��\fndr. ��n#>
B2p��Z�CP Ma�����C38A��� c��6� (���N�B����� �� 2�$�81��!m_���"ex�z 5�.Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$ �r*$��*$r*$%/s#�C�d/.,P�/0*ʲDPN��$���$�*�Gr�$k Ex�c�'IF�$MAS}K�%93 H5�%�H558�$548 H�$4-1�$��#21(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�4�9�0�4a�3�9j0"�M�49�4  �x�4�4tpsh��x�4�P�4- DQ� @�3�Q�4�R�4�pR%0 �2�r�4.b
E\���5�A�4��3adq\>�5K979":E�a~jO l "DQ^E^�3i�Dq ��4�R�O ?R�? ��q�5 ��T��3rAq�O�L#st�5~��7p�5��0REJ#�2�@av^Eͱ��F���4��.�5y �N� �2il(in8�4��31 JH1�2�Q4�251ݠ�4rmal� �3)�REo� Z_�æOx����4��^F�?onorTf��7_�ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4�REM���4yݱ"u@�RER5932fO��4�7Z��5lity,��U��e"Dil\��5��o ��798�7�?�25 �3hk9 10�3��FE�0=0|P_�Hl\mhm�5 ��qe�=$�^�
E���u�IAymptm`�U��BU��vste� y\�3��me�b�DvI� [�Qu�:F�Ub�*_��
E,�su��_ Er��ox���4�huse�E-�?�s�n�������FE��,�b#ox�����c݌," �������z��M�x�g��pdspw)� 	��9���b���(��1���c��Y� R�� �>�P���W��� �����'�0ɵ��[��͂���  ߤ ,@� ��A�bum�pšf��B*�Bo!x%��7Aǰ60�BB�w���MC� (6�,�f�t I�s� ST��*��}B���z��w��"BBF
��>�`���)��\bbk968 "�X4�ω�bb�9vas69����etbŠb��X�����ed	��F��u�f� �seDa"������'�\��@,���b�ѽ�o6�$H�
�x�$�f���!�y���Q[�! tp�err�fd� T�Pl0o� Reco�v,��3D��R642 � 0��C@}s�� N@��(U�rr�o���yu2r���  �
  |����$$CLe�? �������������$z�_D�IGIT��������.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo�$j��+c:PRO�DUCTM�0\P_GSTKD��V&o�hozf99��D����$FEAT?_INDEX��xd���  �
�`ILECO_MP ;���#���`�cSETU�P2 <�e~�b�  N �a��c_AP2BCK� 1=�i  #�)wh0?{%&c����Q�xe%� I�m���8�� \�n����!���ȏW� �{��"���F�Տj� ��w���/�ğS���� �����B�T��x�� ����=�үa������ ,���P�߯t������ 9�ο�o�ϓ�(�:� ɿ^���Ϗϸ�G� ��k� �ߡ�6���Z� l��ϐ�ߴ���U��� y����D���h��� ���-���Q������ ���@�R���v���� )�����_�����* ��N��r��7 ��m�&�3�\�i
pP 2>#p*.VRc�*��� /���PC/1/OFR6:/].��/+T�`�/�/F%�/��,�`r/?�*.F�8?	H#&?e<��/�?;STM @�2�?�.K �?�=�iPendant Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OoO�O_:JPG  _J_�56_�O_�_��	PANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W �o�o�o)�Z4�o[��WI��
T�PEINS.XM)L��0\����qCustom Toolbar	���PASSWO�RDyFRS�:\L�� %P�assword ?Config��� ֏e�Ϗ�B0���T� f����������O�� s������>�͟b�� [���'���K��򯁯 ���:�L�ۯp����� #�5�ʿY��}��$� ��H�׿l�~�Ϣ�1� ����g��ϋ� ߯��� V���z�	�s߰�?��� c���
��.��R�d� �߈���;�M���q� �����<���`���� ��%���I������ ��8����n���! ��W�{"� F�j|�/� Se��/�/T/ �x//�/�/=/�/a/ �/?�/,?�/P?�/�/ �??�?9?�?�?o?O �?(O:O�?^O�?�O�O #O�OGO�OkO}O_�O 6_�O/_l_�O�__�_ �_U_�_y_o o�_Do �_ho�_	o�o-o�oQo �o�o�o�o@R�o v��;�_� ��*��N��G��� ���7�̏ޏm���� &�8�Ǐ\�돀��!� ��E�ڟi�ӟ���4� ßX�j��������į S��w������B�#���$FILE_D�GBCK 1=���/���� ( �)
�SUMMARY.�DGL���MD:����Dia�g Summar�y��Ϊ
CONSLOG�������D��ӱConsol�e logE�ͫ���MEMCHEC�K:�!ϯ���X�M�emory Da�ta��ѧ�{)}��HADOW���ϵ�J���Sha�dow Chan�gesM�'�-�?�)	FTP7Ϥ��3ߨ���Z�mme?nt TBD��ѧ�0=4)ETHERNET��������T�ӱEthe�rnet \�fi�guration�U�ؠ��DCSVR�F�߽߫�����%��� verif�y all��'�1�PY���DIFF������[���%��diff]�����1R�9�K��� ����X��CHGD������c��!r����2ZAS� ���GD���k��8z��FY3bI[� �/"�GD���s/�����/*&UPDA�TES.� �/���FRS:\�/�-�ԱUpdates� List�/��P�SRBWLD.C	M(?���"<?�/Y��PS_ROBOWEL��̯�?�?��? &�O-O�?QO�?uOO nO�O:O�O^O�O_�O )_�OM___�O�__�_ �_H_�_l_o�_�_7o �_[o�_lo�o o�oDo �o�ozo�o3E�o i�o���R� v���A��e�w� ���*���я`����� ����O�ޏs���� ��8�͟\�����'� ��K�]�쟁����4� ��ۯj������5�į Y��}������B�׿ �x�Ϝ�1���*�g� ����Ϝ���P���t� 	�ߪ�?���c�u�� ��(߽�L߶��߂�� ��(�M���q� ��� 6���Z������%��� I���B�����2������h����$FI�LE_� PR� ���������MDON�LY 1=.�� 
 ���q�� ��������~ %�I�m� 2��h��!/� ./W/�{/
/�/�/@/ �/d/�/?�//?�/S? e?�/�??�?<?�?�? r?O�?+O=O�?aO�? �O�O&O�OJO�O�O�O�_�O9_�OF_o_
VISBCKL6[*.VDv_�_.P�FR:\�_�^�.PVision� VD file �_�O4oFo\_joT_�o o�o�oSo�owo �oB�of�o�+ �������+� P��t������9�Ώ ]�򏁏��(���L�^� ������5���ܟk�  ���$�6�şZ��~������
MR_G�RP 1>.�L��C4  B���	 W������*u����RHB ��2� ��� ��� ���B�����Z� l���C���D��������Ŀ��K�PJ���_I���T����F�5UPǎ?����ֿ �E�M.G��E$��;n߇�:G��@O����@��;@�A��f�@�F�B@�#�*λ� F@ ��������J��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<?,6\b��+�@&�(�a�L߅�p�A��A��߲�v���r��� ���
�C�.�@�y�d� �������������`�?�Z�lϖ�BH�� �Ζ��������
0�PS@�P��I$��ܿ� �B�x��/ ��@�33:���.�gN�UUU�U��q	>u.�?!rX���	�-=[z��=�̽=V6�<�=�=��=$q�����@�8�i7G���8�D�8@9!�7�:�����D�@ D�Ϡ Cϥ��C�
�����'/0-��P/ ����/N��/r��/�� �/�??;?&?_?J? \?�?�?�?�?�?�?O �?O7O"O[OFOOjO �O�O�O�O�гߵ��O $_�OH_3_l_W_�_{_ �_�_�_�_�_o�_2o oVohoSo�owo�o�i ��o�o�o��); �o_J�j��� ����%��5�[� F��j�����Ǐ��� ֏�!��E�0�i�{� B/��f/�/�/�/���/ ��/A�\�e�P���t� �������ί��+� �O�:�s�^�p����� Ϳ���ܿ� ��OH� �o�
ϓ�~ϷϢ��� �������5� �Y�D� }�hߍ߳ߞ������� �o�1�C�U�y��� ������������� -��Q�<�u�`����� ����������; &_J\����� �����ڟ�F� j4������� ��!//1/W/B/{/ f/�/�/�/�/�/�/�/ ??A?,?e?,φ?P� q?�?�?�?�?O�?+O OOO:OLO�OpO�O�O �O�O�O�O_'__K_ �o_�_�_�_l��_0_ �_�_�_#o
oGo.oko Voho�o�o�o�o�o�o �oC.gR� v�����	�� �<�`�*<��` �����ޏ��)�� M�8�q�\�������˟ ���ڟ���7�"�[� F�X���|���|?֯�? �����3��W�B�{� f�����ÿ������� ��A�,�e�P�uϛ� b_�����Ϫ_��߀� =�(�a�s�Zߗ�~߻� ��������� �9�$� ]�H��l������ ������#��G�Y� � B�������z������� 
ԏ:�C.gRd ������	� ?*cN�r� ����/̯&/� M/�q/\/�/�/�/�/ �/�/�/?�/7?"?4? m?X?�?|?�?�?�?�? ��O!O3O��WOiO�? �OxO�O�O�O�O�O_ �O/__S_>_P_�_t_ �_�_�_�_�_�_o+o oOo:oso^o�o�op� �o�� ��$�� o�o�~��� ����5� �Y�D� }�h�������׏�� ��
�C�.�/v�<� ��8������П��� �?�*�c�N���r��� �����̯��)��? 9�_�q���JO����� ݿȿ��%�7��[� F��jϣώ��ϲ��� ����!��E�0�i�T� yߟߊ��߮��߮o�o ��o>�t�>�� b�����������+� �O�:�L���p����� ��������'K 6oZ�Z�|�~�� ���5 YD i�z����� �/
//U/@/y/@� �/�/�/�/���/^/? ??Q?8?u?\?�?�? �?�?�?�?�?OO;O &O8OqO\O�O�O�O�O��O�O�O_�O7_���$FNO ����VQ_�
F0fQ kP� FLAG8�(�LRRM_CHKT_YP  WP��^P�WP�{QO=M�P_MIN�P�����P�  �XNPSSB_CF�G ?VU ��_���S� ooIUTP_DEF_OW  ���R&hIRCOM��P8o�$GENO�VRD_DO�V��6�flTHR�V �d�edkd_ENB�Wo k`RAVC_GRP 1@�WCa X"_�o_ 1U<y�r� ����	��-�� =�c�J���n������� �ȏ����;�"�_�pF�X���ibROU�`�FVX�P��&�<b&�8�?���埘�������  D?�јs���@@g�B�7�p�)�ԙ���`SMT�cG��mM���� �LQHoOSTC�R1H����P��at�S5M��f�\���	127.0��=1��  e��ٿ �����ǿ@�R�d��vϙ�0�*�	ano?nymous����0�������/�[��
 � �����r��� �ߨߺ�����-��� &�8�[�I�π��� ����1�C��W� y���`�r������ߺ� ������%�c�u�J \n�������� �M�"4FX�� i������7 //0/B/T/��� m/��/�/�/?? ,?�/P?b?t?�?�/�? ��?�?�?OOe/w/ �/�/�?�O�/�O�O�O �O�O=?_$_6_H_kO Y_�?�_�_�_�_�_'O 9OKO]O__Do�Ohozo �o�o�o�O�o�o�o
 ?o}_Rdv�� �_�_oo!�Uo*� <�N�`�r��o������ ̏ޏ�?Q&�8�J��\���>�ENT 1=I�� P!􏪟  ����՟ğ �������A��M�(� v���^�����㯦�� ʯ+�� �a�$���H� ��l�Ϳ�����ƿ'� �K��o�2�hϥϔ� �ό��ϰ������� F�k�.ߏ�R߳�v��� ���߾���1���U���y�<�QUICCA0��b�t����1������%���2&����u�!ROUTE�Rv�R�d���!P�CJOG����!�192.168�.0.10��w�N�AME !��!?ROBOTp��S_CFG 1H��� ��Auto-sta�rted�tFTP������ � 2D��hz ����U��
/ /./�v���/� ��/�/�/�/�/�!? 3?E?W?i?�/?�?�? �?�?�?�?���AO �?eO�/�O�O�O�O�? �O�O__+_NO�OJ_ s_�_�_�_�_
OO.O oB_'ovOKo]ooo�o P_>o�o�o�o�oo �o5GYk}�_�_ �_��8o��1� C�U�$y�������� ӏf���	��-�?�� ���Ə���ϟ� ����;�M�_�q� ��.�(���˯ݯ�� P�b�t�����m����� ����ǿٿ�����!� 3�E�h��{ύϟϱ� ���$�6�H�J�/�~� S�e�w߉ߛ�jϿ��� �����*߬�=�O�a��s��YT_ERR� J5
���PDUSIZ  ��^J����>��W�RD ?t���  guest}��%�7�I��[�m�$SCDMN�GRP 2Kt;�������V$�K�� 	P01.14 8���   y�����B    �;����� ��������
 �������������~����C�.gR|��� � i  � � 
��������� +��������
���l .Vr���"�l��� m
d�������_GROU��L.�� �	�����07EQUPD � 	պ�J�T�Ya ����TT�P_AUTH 1�M�� <!i?Pendany���6�Y!KAREL:*��
-�KC///A/ �VISION SCETT�/v/�" �/�/�/#�/�/
??�Q?(?:?�?^?p>�C?TRL N�����5�
�FF�F9E3�?�F�RS:DEFAU�LT�<FAN�UC Web S_erver�:
� ����<kO}O�O�O�O��O��WR_CON�FIG O�� ��?��IDL_�CPU_PC@��B��7P�BH�UMIN(\��<TGNR_IO��������PNPT_SI�M_DOmVw[T�PMODNTOL�mV �]_PRTY��X7RTOLNK 1P����_o!o�3oEoWoio�RMAS�TElP��R�O_gCFG�o�iUO�|�o�bCYCLE�o��d@_ASG 19Q����
 ko, >Pbt����������sk�bN�UM����K@�`I�PCH�o��`RTRY_CN@oR���bSCRN����Q���� �b�`�bR���Տ��$J2�3_DSP_EN�	����OBP�ROC�U�iJO�GP1SY@��8�?�!�T�!�}?*�POSRE�~zVKANJI_�` ��o_�� ��T�L�6�͕����CL_L�GP<�_���EYLO�GGIN�`����LANGUA�GE YF7R�D w���LG��U��?⧈�x� ������=P��'0���$ NMC�:\RSCH\0�0\��LN_DISP V��
�ј������OC�R.RD�zVTA{�OGBOOK W
{��i0��ii��X���@��ǿٿ�����"��6	h������e�?�G_BUFF� 1X�]��2 	աϸ��������� ��!�N�E�W߄�{� �ߺ߱�����������J���DCS �Zr� =��� �^�+�ZE��������a�IO 1[
{# ُ!� �!�1� C�U�i�y��������� ������	-AQ cu�������EfPTM  �d �2/ASew� ������// +/=/O/a/s/�/�/��NSEV����TYP�/??y͒�RS@"���>��FL 1\
������?�?�?�?�?��?�?/?TP6���">�NGNAMp�ե�U`�UPS���GI}�𑪅mA_�LOAD�G �%�%DF_M�OTN���O�@MA?XUALRM<��@J��@sA�Q����WS ��@C �]m�-_����MP2�7�^
{ �ر�	�!P�+bʠ�;_/��Rr�W�_�WU�W�_��R 	o�_o?o"ocoNoso �o�o�o�o�o�o�o �o;&Kq\�x �������#� I�4�m�P���|���Ǐ ���֏��!��E�(� i�T�f�����ß��ӟ ���� �A�,�>�w� Z�������ѯ����د ���O�2�s�^��� ����Ϳ���ܿ�'���BD_LDXDI�SAX@	��MEM�O_APR@E ?=�+
 � *� ~ϐϢϴ���������~�@ISC 1_�+ ��IߨT��Q� c�Ϝ߇��ߧ����� w����>�)�b�t�[� ����{�������� ��:���I�[�/���� ��������o�����6 !ZlS��s ����2�A S'�w���� g��.//R/d/��_MSTR `��-w%SCD 1am͠L/�/H/�/�/? �/2??/?h?S?�?w? �?�?�?�?�?
O�?.O ORO=OvOaO�O�O�O �O�O�O�O__<_'_ L_r_]_�_�_�_�_�_ �_o�_�_8o#o\oGo �oko�o�o�o�o�o�o �o"F1jUg �������� �B�-�f�Q���u������ҏh/MKCFG� b�-㏕"L_TARM_��cL�w� σ�Q�N�<�METPU�I�ǂ���)NDSP_CMNTh�p��|�  d�.���ς�ҟܔ|�P�OSCF����PSTOL 1e'�{4@�<#�
5� ́5�E�S�1�S�U�g� ������߯��ӯ��� 	�K�-�?���c�u������|�SING_C�HK  ��;�ODAQ,�f��Ç�~�DEV 	L��	MC:!�HS�IZEh��-��T�ASK %6�%�$1234567�89 �Ϡ��TR�IG 1g�+ l6�%���ǃ�����8�p�YP[� ���EM_INF 1�h3� �`)AT&FVg0E0"ߙ�)���E0V1&A3&�B1&D2&S0�&C1S0=��)�ATZ������H@�����A���AI�@q�,��|���� � ��ߵ�����J���n� �����W��������� ��"����X��/� ���e������ 0�T;x�=� as��/�,/c =/b/�/A/�/�/�/ �/��?���^? p?#/�?�/�?s?}/�? �?O�?6OHO�/lO? 1?C?U?�Oy?�O�O3O  _�?D_�OU_z_a_�_~�ONITOR���G ?5�   	EXEC1Ƀ��R2�X3�X4�X5��X���V7�X8�X9Ƀ�RhBLd�RLd�R Ld�RLd
bLdbLd"b�Ld.bLd:bLdFbLc2�Sh2_h2kh2wh2��h2�h2�h2�h2��h2�h3Sh3_h3��R�R_GRP_�SV 1in���(�����C?BP�P�A4�>%���gY�>r���x�_D=R^���PL_NAME �!6��p�!�Default �Personal�ity (fro�m FD) �R�R2eq 1j)T?UX)TX��q��X dϏ8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|������2'�П������*�<�N�`�r��< ��������ү����@�,�>�P�b� �Rdrg 1o�y �\�O, �3����� @D�  ��?������?䰺��A�'�6����;��	lʲ	 �xJ������ �<� �"�� ��(pK�K ���K=*�J����J���JV����Z������rτ́p@j�@wT;f���f���ұ]�l��I��7�������������b��3��´7  ��`�>�����bϸ�z���=�����Jm��
� B�H�˱]����q�	� p� W P�pQ�p��p|  Ъ�g����c�	'� � ���I� � � ����:����
�È=����"�nÿ�	�ВI  �n @B� cΤ�\��ۤ��q��y�o�N���  '������@2�@�����/��C��C�C�@ �C������
��A��* # W @<�P�R�%
h�B�b�A��j������������Dz ۩��߹�����j���( �� -��C���'�7L������Y������ �?�ff ���gy ����o�:a��
�>+�  PƱj�( ����7	���^|�?����xZ��p<
6b<���;܍�<����<� <�&Jσ�AI�ɳ+�|���?fff?I��?&�k�@�.���J<?�` �q�.�˴fɺ�/ ��5/����j/U/�/ y/�/�/�/�/�/?�/0?q��F�?l? ?�?/�?+)�?�?ؿE�� E�I�G+� F��?)O �?9O_OJO�OnO�Of�BL޳B�?_h�.� �O�O��%_�OL_�?m_ �?�__�_�_�_�_�
��h�Îg>���_Co�_goRodo��o�GA�ds�q�C��o�o�o|���ؠ$]Hq���D���pC���pCHmZZ7t���6q�q���ܶN'�3A�A��AR1AO��^?�$�?��K/�±
=ç�>����3�W�
=�#�W��eۣצ�@�����{����<�����(�B�u���=B0������	L���H�F�G����G��H�U�`E���C�+����I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3�l� W���{��������՟ ���2��V�A�z��� w�����ԯ������ ��R�=�v�a����� �������߿��<� '�`�Kτ�oρϺϥ� �������&��J�\� G߀�kߤߏ��߳��� ����"��F�1�j�U� ��y���������� ��0��T�?�Q�����(���3/E�y���u����<��M3�8�����M4Mgs&�IB+2D�a���{�^^	�@�����uP2	P7Q4_A��M00bt��R��`����/   �/�b/P/�/t/�/  *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?��?�?O 2 F;�$�vGb�/�Aa��@�a�`�qC��C�@�o�Ot���KF�� DzH@�� F�P D���O�O�ys<O!_3_E_�W_i_s?���@U@pZ�422�!2~
  p_�_�_�_	oo-o?o Qocouo�o�o�o�o��Q ��+��1���$MSKCF�MAP  �5?� �6�Q��Q"~�cONREL7  
q3��bEXCFENB�?w
s1uXqFNC�_QtJOGOVLKIM?wdIpMrd�bWKEY?w�u�bWRUN�|�u�bSFSPDTY�xavJu3sSIGN?>QtT1MOT�Nq��b_CE_GRoP 1p�5s\r���j�����T�� ⏙������<��`� �U���M���̟��� ���&�ݟJ��C��� 7�������گ��������4�V�`TCOM_CFG 1q}��Vp�����
P�_/ARC_\r
jyUAP_CPL���ntNOCHECK� ?{  	r��1�C�U�g� yϋϝϯ����������	��({NO_WA�IT_L�	uM�NMTX�r{�[m�o_ERRY�2sy3� &��������r�c� ��T_�MO��t��, �j#$�k�3�PAR�AM��u{��	�[���u?�� =�9@345678901��&���E�W� 3�c�����{������������=��UM_RSPAC�E �Vv��$ODRDSP���jx�OFFSET_C�ARTܿ�DIS���PEN_FI�LE� �q��c֮�O�PTION_IO���PWORK kv_�ms �(P(�R�@�6$j.j	 ��Hj(�6$�p=�_DSBL'  �5Js�\���RIENTTO>p9!C��PqfA�� UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?p]a]�D�WcUa쪋l;�	�lmb�`�x7J�`�p����a�< ���`�m�a��H(���H3k7HSM�5G�22G���Gp
��
��c�'|��CR�	>�>q�GsuaT��3���  �4 spBpyr  ]o�*S�B_����j�]��t�q� ��rna �,����6  ��P�Q�|N��M�,k���	'� �� ��I� �  ��%�=��ͭ���ba�	���I  �n @��~���Dp�������N	 W�  '!o�:q�pC	 C�@@sBq�t|��� m�
�!*�h@ߐ�n����*�B	 �A���p�G �-�qbz��P��t�_�������( �� -��恊�n�ڥ[A"]Ѻ�b4�'!5�(p? �?�ff� ��
����OZ�R*��85�z���>΁  	Pia��(5���@����ک�a�c�dF#?��5�x��*�<
6�b<߈;܍��<�ê<� <�&�o&�)��A�lcΐI�*�?f7ff?�?&c����@�.uJ<?�`��Yђ^� nd��]e��[g��Gǡd <����1��U�@�y� dߝ߯ߚ����߼�	� ��-������&��"�E�� E��G+� Fþ����� �������&��J�5��bB��AT�8�ђ ��0�6���>���J� n�7��[m�0���h��1��>��M�I
��@��A�[��C�-�)��?�A��� /�YĒ�a�Jp��vav`CH/�������}!@I��Y�'�3A��A�AR1AO��^?�$�?�����±
=���>����3�?W
=�#����+�e��ܒ������{����<�����.(�B�u���=B0������	��*H�F�G����G��H�U�`E���C�+��-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�?O �?3OOWOBOTO�OxO �O�O�O�O�O�O_/_ _S_>_w_b_�_�_�_ �_�_�_�_oo=o(o aoLo�o�o�o�o�o�o �o�o'$]H �l������ �#��G�2�k�V��� z���ŏ���ԏ��� 1��U�g�R���v��� ��ӟ�������-���(�������y�a����Q�<c�,!3�8�}���,!4Mgs����ɢ�IB+կ篴a���{���A�@/�e�S���w��P!�	P�������7��0ӯ�ϑ�R9�K�`��oχϓϥ�  ���χ����)��M� �����z���{߉ߛ���ߒߤ�������  )�G�q�_����2 F;�$�&Gb���n�a�[ZjM!C�s��@j/�A�S�=�F�� Dz��� F�P D��W����)������������x?���@U@
9�=�=���=��
  v������ �*<N`�*�P ���˨�1���$PARAM�_MENU ?�-�� � DEFP�ULSEl	W�AITTMOUT��RCV� �SHELL_W�RK.$CUR_oSTYL�,�OPT�/PTB�./("C�R_DECSN���,y/�/ �/�/�/�/�/?	??�-?V?Q?c?u?�?�U�SE_PROG �%�%�?�?�3C�CR�����7_HOST !�#!�44O�:T̰�?�PCO)ARC�O�;_�TIME�XB� � �GDEBU�GV@��3GINP?_FLMSK�O�IqT`��O�EPGAPe �L��#[CH�O^�HTYPE����?�?�_�_�_�_�_ oo'o9obo]ooo�o �o�o�o�o�o�o�o :5GY�}�� �������1��Z��EWORD ?}	7]	RS`�_	PNS�$斂JOE!>�TE�s@WVTRACEC�TL 1x-�� �� ������ɆD/T Qy-��䀿D � ��7�4�P  :�L :�GP:�D :�@ :�8�,�>�P�b��� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� V�(�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_d��_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�_���*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p�������� //$)�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �#|"DEF�SPD |�,l!!J �8 IN �TRL }�-�" 8�%�!PE_C�ONFI� ~g%O�g!�$�%��$LID�#�-~74GRP 1�7�Q!�#!A ����&ff"!A+�33D�� D]�� CÀ A@+6�!�" d�$�9�9�*1*0� 	 �+9�(�&�"�? ´	C�?�;B@3AO�?�OIO3OmO"!>�T?�
5�O�O�N��O =��=#�
�O_�O_J_5_ n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_Roxoco�o �o�o�o�o�o�o�>)bM��;
�V7.10bet�a1�$  �A�E�rӻ��A " �p?!G�^�q>���r��0��q�ͻqBQ��qA\�p�q�4�q*�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏� ��4��1�j�U���y� ����֟������0� �T�?�x�c������� ү����!o�,�ۯP� ;�M���q�����ο�� �ݿ�(��L�7�p�x+9��sF@ �� �ͷϥ�g%������ +�!6I�[߆������� �ߠ���������!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ���=(aL ^������ �'9$]�Ϛ��� ��������/<� 5/`�r߄ߖߏ/>�/ �/�/�/�/?�/1?? U?@?R?�?v?�?�?�? �?�?�?O-OOQO<O uO`O�O�O�O�O���O _�O)__M_8_q_\_ n_�_�_�_�_�_�_o �_7oIot���o�o ���o�o�o(/!L/ ^/p/�/{*o��� ������A�,� e�P�b���������� Ώ��+�=�(�a�L� ��p������Oߟ񟠟 � �9�$�]�H���l� ~�����ۯƯ���#� No`oro�on��o�o�o �oԿ���8J\ ng����vϯϚ��� ����	���-��Q�<� u�`�r߫ߖ��ߺ��� ����;�M�8�q�\� ��������z������ %��I�4�m�X���|� ����������:�L� ^���Z�������� ���$�6�H�S wb����� ��//=/(/a/L/ �/p/�/�/�/�/�/? �/'??K?]?H?�?�� �?�?f?�?�?�?O�? 5O OYODO}OhO�O�O �O�O�O�O&8J4_ F_����_�_��_ �_"4-o�O*oco No�oro�o�o�o�o�o �o)M8q\ �������� �7�"�[�m��?���� R�Ǐ���֏�!�� E�0�i�T���x����� ���_$_V_ �2�l_�~_�_�����R�$P�LID_KNOW�_M  �T������SV� ��U͠�U��
��.� ǟR�=�O�����mӣ�M_GRP 1�T�!`0u��T@ٰ)o�ҵ�
���P зj��`���!�J� _�W�i�{ύϟϱ���`������߱�MR��Ņ��T��s�w�  s��ߠ޴߯߅��ߩ� ������A���'�� ����������� ��=���#����������}������S��ST^��1 1��U# ����0�_ A  .��,>Pb�� ������3 (iL^p���(��2*��'�<-/3/)/;/M/4f/x/�/�/�5�/�/�/�/6 ??(?:?7S?e?w?�?8�?�?�?�?~MAD  d�#`PARN_UM  w�\%OSCH?J ME�
�G`A�Iͣ�EUP�D`OrE
a�OT_CMP_��B@�P@�'˥TER_C;HK'U��˪?R�$_6[RSl�¯��_#MOA@�_�U_�_RE�_RES_G � �>�oo8o+o\o Oo�oso�o�o�o�o�o@�o�o�W �\�_ %�Ue Baf�S�  ����S0��� �SR0��#��S�0>� ]�b��S�0}������R�V 1�����rB@�c]��t�(@�c\����D@�c[�$���RTHR_INRl�DA��z˥d,�MASS9�� ZM�MN8�k�M�ON_QUEUE� ���˦��x� URDNPUbQN{�P[��END���_ڙ�EXE�ڕ�@BE��ʟ��OPTIO�Ǘ�[��PROGR�AM %��%�ۏ�O��TASK�_IAD0�OCFG� ���tO��ŠD�ATA���Ϋ@��27�>�P�b�t� ��,�����ɿۿ������#�5�G���INFOUӌ�������� �Ͽ���������+� =�O�a�s߅ߗߩ߻�@�������^�jč�� yġ?PDIT� �ίc���WE�RFL
��
RG�ADJ �n�A	����?����@���?IORITY{�QV}���MPDSPH������Uz����O�TOEy�1�R�� (!AF4�E��P]���!tc�ph���!ud|��!icm���ݏ6�XY_ȡ��R��ۡ)� *0+/ ۠�W :F�j���� ��%7[B��*��PORTT#�BC۠�����_CARTREP�
�R� SKSTA�z��ZSSAV����n�	2500H863���r�$!�U�R����q��n�}/�/�'� URGeE�B��rYWF� #DO{�rUVWV��$��A�WRUP_DELAY �R�>�$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?3A_QSKIP!�n�;l#x 	1/+O + OROdOvO9Hn��O �G�O�O�O�O�O_�O _D_V_h_._�_z_�_ �_�_�_�_
o�_.o@o Roovodo�o�o�o�o �o�o�o*<L�r`���n��$�RCVTM���]��pDCR!�L�ЈqB��C�*J�C$�>��$ >5?-;���04M¹�O���ǃ�������~��9On�Y��<
6b<߈�;܍�>u.��?!<�& {�b�ˏݏ��8���� �,�>�P�b�t����� ����Ο���ݟ�� :�%�7�p�S������ ʯܯ� ��$�6�H� Z�l�~�������ƿ�� �տ���2�D�'�h� zϽ��ϰ��������� 
��.�@�R�d�Oψ� �߅߾ߩ������� ��<�N��r���� ����������&�8� #�\�G�����}����� ������S�4FX j|������ ���0T?x �u����'/ /,/>/P/b/t/�/�/ �/�/�/�/�?�/(? ?L?7?p?�?e?�?�? ��?�? OO$O6OHO ZOlO~O�O�O�?�?�O �O�O�O __D_V_9_ z_�_�?�_�_�_�_�_ 
oo.o@oRodovo�X��qGN_ATC �1�� AT&FV0E/�� ATDP/6/9/2/9�h�ATA�n,�AT%G1%B�960/�++U+�o,�aH,�q�IO_TYPE � �u�sn_�oR�EFPOS1 1}�P{ x�o�Xh_�d_��� ��K�6�o�
���.�ාR����{{2 1�P{���؏V�ԏxz����q3 1���$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����<�>��S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB��-�f��S8 1� ����Y�������y��SMASK 1��P  
9�G��XNOM���a~߈�~�qMOTE  h��~t��_CFG ᢥ����рrPL_�RANG�ћQ��POWER ��e���SM_DRYPRG %i��%��J��TART� �
�X�UME_PRO'�9��~t�_EXEC_EN�B  �e��GS�PD������c��T3DB���RM���MT_!�T����`OBOT_NA_ME i�����iOB_ORD_�NUM ?
��\qH863�  �T���������bPC_TIMoEOUT�� x�`oS232��1��k� LTEA�CH PENDA1N �ǅ�}����`Mainte�nance Co#ns�R}�m
"{�d?KCL/Cg��Z� ��n� ?No Use}�8	��*NPO��Ѯ����(C7H_L��������	�mMAVA#IL��{��ՙ��SPACE1 2��| d��(>��&���p��M,?8�?�ep/ eT/�/�/�/�/�W/ /,/>/�/b/�/v?�? Z?�/�?�9�e�a�=? ?,?>?�?b?�?vO�O�ZO�?�O�O�Os�2�/O*O<O�O`O �O�_�_u_�_�_�_�_[3_#_5_G_Y_o }_�_�o�o�o�o�o[4.o@oRodovo $�o�o����"�	�7�[5K]o� �A����	�̏�?�&�T�[6h�z��� ����^�ԏ���&�� ;�\�C�q�[7���� ����͟{���"�C�@�X�y�`���[8�� ��Ưدꯘ��0�?π`�#�uϖ�}ϫ�[Gw �i� ��:�
G� ���� $�6�H�Z�l�~ߐ��8  ǳ�����߈��d(���M�_�q�� ����������?� ��2�%�7�e�w����� ��������������� !�RE�W����� �����?�Q `�� @ 0��ߖrz	�V_�����
/ L/^/|/2/d/�/�/�/ �/�/�/?�/�/�/*? l?~?�?R?�?�?�?�?@�?�?�?2O�?
���O[_MODE � �˝IS �"��vO,*ϲ��O-_��	M_v_#dCWORK_AD�M���%aR  ���ϰ�P{_�P_?INTVAL�@�����JR_OPTI[ON�V �EBp�VAT_GRP �2����#(y_Ho �e_vo �o�oYo�o�o�o�o�o *<�bOoNDp w������	� ��?�Q�c�u����� /���ϏᏣ����)� ;���_�q��������� O�ɟ���՟7�I� [�m�/�������ǯٯ 믁��!�3���C�i� {���O���ÿտ��� ϡ�/�A�S�e�'ω� �ϭ�oρ������� +�=���a�s߅�Gߕ� �����ߡ���'�9� K�]��߁����y� ���������5�G�Y���E�$SCAN_GTIM�AYuew��R �(�#(�(�<0.a+aPaP
TqA>��Q��oX�����OO�2/��:	d/JaR��WY��^��p�^R^	r  P���� � � 8�P�	�D��GYk} ��������Qp/@/R/x/)P;�o\T���Qpg-�t�_DiKT��[  � lv%��� ���/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OWW �#�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o lO~Od+No`oro�o�o �o�o�o�o�o& 8J\n����8��u�  0�"0g �/�-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q�����$o ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E��� ��Do��������ҿ� ����,�>�P�b�t� �ϘϪϼ���������w
�  58�J�\� n߀ߒߜկ������� ��	��-�?�Q�c�u�p����� �� -����� �2�D�V�@h�z�������������������& ���%	123�45678�" +	��/� ` r������� �(:L^p ������� / /$/6/H/Z/l/~/� �/�/�/�/�/�/? ? 2?D?V?h?�/�?�?�? �?�?�?�?
OO.O@O o?dOvO�O�O�O�O�O �O�O__*_YON_`_ r_�_�_�_�_�_�_�_ ooC_8oJo\ono�o �o�o�o�o�o�oo "4FXj|���������	���s3�E�W�{�C�z  Bp��  � ��2���z��$SCR_GRP� 1�(�U8(�\x^ �@  �	!�	 ׃�� �"�$� ��-��+���R�w����D!~�����#����O����M-10i�A 890990�5 Ŗ5 M61CA >4��Jׁ
� ���0�����#�1�	"�z���О���¯Ҭ � ��c���O�8�J� ������!�����\ֿ��B�y����������A��$�  !@��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ �϶�������%��I� 4�m��<�l߃ߕ��߹�B���\���� 1��U�@�R��v�� ����������;���*<=�
F���?�<d�<�>7�����s@�:��� B����ЗЙ���EL�_DEFAULT�  �����B�MIP�OWERFL  ��$1 WFD�O $��ER�VENT 1������"�pL!�DUM_EIP���8��j!AF�_INE �=�!'FT���9!��4 ��[�!RPC_MAIN\>�J�n'VISw=���o!TP�PU��	d�?/!
PM�ON_PROXY@/�e./�/"Y/��fz/�/!RDMO_SRV�/�	g�/�#?!R C?�h,?o?!
pM�/��i^?�?!RLSgYNC�?8�8�?>O!ROS�.L�4�?SO"wO�#DO VO�O�O�O�O�O_�O 1_�OU__._@_�_d_ v_�_�_�_�_o�_?o�ocoiICE_K�L ?%y (�%SVCPRG�1ho8��e���o�m3��o�o�`4 �`5�(-�`6PU�`7@x}�`���l9��{�d:?��a�o� �a�oE��a�om��a ���aB���aj叟a ���a�5��a�]� �a����a3����a[� ՟�a�����a��%��a ӏM��a��u��a#��� �aK�ů�as���a�� mob�`�o�`8�}�w� ������ɿ���ؿ� ��5�G�2�k�VϏ�z� �Ϟ����������1� �U�@�y�dߝ߯ߚ� �߾�������?�*� Q�u�`������� �����;�&�_�J� ��n������������sj_DEV ~y	�MC:���_OUT�",REC� 1�Z� d �   	�    ��@�� ����A�����
 �PS?D#6 r��UO� �� �� `��� �Z�{� �r� *�  +X�- � I- �- !
- � �X�YZ��PSJ;4 ��?  (� E � ��R ���� E- �� �/e/�l!4�/��� X� (,/>/P/�/�/*�""4� =�!� � ؀  ?"S1h��'!�/���("- ��\?�?$=�= �?�?�?"OOFO4OjO |O^O�O�O�O�O�O�O �O_ __T_B_x_f_ �_�_�_�_�_�_�_o ooPo>oto�oho�o �o�o�o�o�o(
 L:\�p���w,����4� "�X�F�|���p����� ֏ď����0��@� f�T���x�����ҟ� Ɵ���,��<�b�P� ��h�z������ί� �(�:��^�L�n�p� ������ܿ�п� � 6�$�Z�H�jϐ�rϴ� �����������2�D� &�h�Vߌ�z߰ߞ��� ��������
�@�.�d��R��ZjV 1��w P����j� 
�� ��<��
TYPEV�FZN_CFG ;��5d��4�GRP 1��A�c ,B� A�� D;� B����  B4�RB21HE�LL:�(
��?x���<%RS'! ��H3lW� {������`2Vh������%w�����#!�1�����7�2�0d�����HK 1��� �k/f/x/�/�/�/ �/�/�/�/??C?>?�P?b?�?�?�?�?��OMM ����?���FTOV_ENB� ���+�HOW_R�EG_UIO��I_MWAITB�.JKOUT;F��LIwTIM;E���O�VAL[OMC_UN�ITC�F+�MON�_ALIAS ?�e�9 ( he ��_&_8_J_\_B_ �_�_�_�_j_�_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]n��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� ���������ӟ~��� 	��-�?��c�u��� ����V�ϯ����� �;�M�_�q������ ��˿ݿ����%�7� I���m�ϑϣϵ�`� ������ߺ�3�E�W� i�{�&ߟ߱������� ����/�A�S���w� ����X������� ���=�O�a�s���0� ������������' 9K]���� b���#�G Yk}�:��� ���/1/C/U/ / f/�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_O
O�O�O�O �O�OvO�O__%_7_��C�$SMON_�DEFPRO ����`Q� *SY�STEM*  d�=OURECAL�L ?}`Y (� �}*copy� mdb:*.*� virt:\t�mpback\=�>inspiron:5076 �V��_�_�_	o  }.=x�Rfr:\�_*`@�]�_`oro�oe/ ea(o:o�PPo�o�o�d
xyzrate 61 �o�o�o�`r�e w�X4060 :L����h3!ds:or�derfil.dat�_�zS�e�w��� `�_:��uK�܏� � o%o8�sϏ`�r��� �o(�:��pP���� �*���Ώ_�q����������L�ݯ���6� �2�emp�P192.168.4E�?46:795�f�px���� �*.d4��F�O����1 �����Ͽ`�rτ���y;�6 @�R��������tpdisc 0�ϼ¿���b��t߆��tpconn 0 )�;�M� ������'߹���\� n���ҩ�9�K������ ��ϥ�N�6244����b�t����+��=�O������)�792����as��9 �2�*<����0���3
�btĆ�4 ���=4 pU��
/ }5�� ���g/y/�/0/�B/T/�/�/	?��580 �/�/c?u?�? ��567�?�?�? "�?58�?bOtO�O���?5�O 1652  WO�O�O�O���O�I�O `_r_�_�/)�;_M_�_ �_o?'?�T�_�_co uo�o�?�?5O�G�o�o �oO"O�o�H�obt ���/�/KtV�� �/��>`�h�z� ��o�o:����
� ��Aӏd�v�������$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1����?���%֟ ��&�	��\�?�f� ��u��������ϯ�� "��F�)�;�|�_��� ����ֿ��˿��� B�%�f�I�[Ϝ�Ϧ� �ϵ�������,��6� b�E߆�i�{߼ߟ��� ��������L�/�V� ��e��������� ���6��+�l�O�v� �������������� 2V9K�o� ������& R5vYk��� ��/��<//F/ r/U/�/y/�/�/�/�/ ?�/&?	??\???f? �?u?�?�?�?�?�?�? "OOFO)O;O|O_O�O �O�O�O�O�O_�O_ B_%_f_I_[_�__�_ �_�_�_�_�_,oo6o boEo�oio{o�o�o�o �o�o�oL/V �e������ ��6��+�l�O�v��������PARAM� ����� ��	��P�����OFT_K�B_CFG  �⃱���PIN_S_IM  ����C�U�g�����RVQSTP_DSB,��򂣟����SR ��/�� & gCAR������TOP_ON_E�Rސ���P_TN /�@��A	�RIN�G_PRM� ���VDT_GRP� 1�ˉ�  	������������Я �����*�Q�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߣߠ� ������������0� B�i�f�x������ �������/�,�>�P� b�t������������� ��(:L^p �������  $6HZ�~� ������/ / G/D/V/h/z/�/�/�/ �/�/�/?
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O�__&_8___\_��V�PRG_COUN�T��@���RENBU��UM�S��__UPD 1�/�8  
s_�o o*oSoNo`oro�o�o �o�o�o�o�o+& 8Jsn���� �����"�K�F� X�j���������ۏ֏ ���#��0�B�k�f� x���������ҟ���� ��C�>�P�b����� ����ӯί������UYSDEBUG��P�P�)�d�YH�S�P_PASS�U�B?Z�LOG ���U�S)��#�0�  ��Q)�
MC:\��6���_MPC���U�ϒ�Qñ8� �Q�S_AV �����lǲ%�ηSV;��TEM_TIMEw 1��[ (�P��Ty�ؿT1S�VGUNS�P�U'��U���ASK_?OPTION�P�U��Q�Q��BCCF�G ��[u� n�X�G�`a�gZo� �߃ߕ��߹������ �:�%�^�p�[��� ������� �����6� !�Z�E�~�i���������%�������&8 ��nY�}�?� �ԫ ��( L:p^���� ���/ /6/$/F/ l/Z/�/~/�/�/�/�/ �/�/�/2?8 F?X? v?�?�??�?�?�?�? �?O*O<O
O`ONO�O rO�O�O�O�O�O_�O &__J_8_n_\_~_�_ �_�_�_�_�_o�_ o "o4ojoXo�oD?�o�o �o�o�oxo.T Bx��j��� �����,�b�P� ��t�����Ώ��ޏ� �(��L�:�p�^��� ����ʟ��o�� 6�H�Z�؟~�l����� ��د���ʯ ��D� 2�h�V�x�z���¿�� �Կ
���.��>�d� Rψ�vϬϚ��Ͼ��� ����*��N��f�x� �ߨߺ�8�������� �8�J�\�*��n�� �����������"�� F�4�j�X���|����� ��������0@ BT�x�d��� ��>,Nt b������/ �(//8/:/L/�/p/ �/�/�/�/�/�/�/$? ?H?6?l?Z?�?~?�? �?�?�?�?O�&O8O VOhOzO�?�O�O�O�O �O�O
__�O@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<o^o�o ro�o�o�o�o�o�o  J8n$O�� ���X���4��"�X�B�v��$TB�CSG_GRP �2�B���  �v� 
 ?�  ������ ׏�������1��U��g�z���ƈ�d�, ���?v�	 �HC��d�>�����e�CL  Bጙ�Пܘ������\)��Y  3A�ܟ$�B�g�B�#Bl�i�X�ɼ���>X��  D	J���r�����C����үܬ���D�@v�=�W� j�}�H�Z���ſ���������v�	�V3.00��	�m61c�	�*X�P�u�g�p�>�d��v�(:�� ���p͟�  O�����p�����z�JCFoG �B���Y ���������=��=�c�q� K�qߗ߂߻ߦ����� ���'��$�]�H�� l������������ #��G�2�k�V���z� ������������ �p*<N���l� ������#5 GY}h��� �v�b��>�// / V/D/z/h/�/�/�/�/ �/�/�/?
?@?.?d? R?t?v?�?�?�?�?�? O�?*OO:O`ONO�O rO�O�O��O�O�O_ &__J_8_n_\_�_�_ �_�_�_�_�_�_�_o Fo4ojo|o�o�oZo�o �o�o�o�o�oB0 fT�x���� ���,��P�>�`� b�t�����Ώ����� ��&�L��Od�v��� 2�����ȟʟܟ� � 6�$�Z�l�~���N��� ��دƯ�� �2�� B�h�V���z�����Կ ¿����.��R�@� v�dϚψϪ��Ͼ��� ����<�*�L�N�`� �߄ߺߨ����ߚ�� �����\�J��n�� ���������"��� 2�X�F�|�j������� ��������.T Bxf����� ��>,bP �t�����/ �(//8/:/L/�/�� �/�/�/h/�/�/�/$? ?H?6?l?Z?�?�?�? �?�?�?�?O�?ODO VOhO"O4O�O�O�O�O �O�O
_�O_@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<oro`o �o�o�o�o�o�o�o &�/>P�/�� �������4� F�X��(���|����� ֏����Ə0��@� B�T���x�����ҟ�� ����,��P�>�t� b������������� ��:�(�^�L�n��� ����2d�����̿ �$�Z�H�~�lϢϐ� �������Ϻ� ��0� 2�D�zߌߞ߰�j��� �������
�,�.�@� v�d��������� ����<�*�`�N��� r������������� &J\�t�� B������ F4j|��^����/�  2 6# 6&J/6"��$TBJOP_�GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� ƞ6$ @2 �"	� �C�� �&b�  Cق'�!�!>ǌ��
559>��0+1�33=��CL� fff?>+0?�ffB� J1��%Y?d7�.��/>;��2\)?0��5���;��h{CY� �  @� ~�!B�  A�P?��?�3EC�  D��!�,�0*BO���?�3JB��
:�/��Bl�0��0�$��1�?O6!Aə�3AДC�1D�G6Ǌ=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__<�O�O>B�\JU�O�HH�1ts�A@g33@?1� C�� ��@�_�_&_8_>��D�UV_0�LP�Q30O<{�zR� @�0 �V�P!o3o�_<oRifo Po^o�o�o�oRo�o�o �o�oM(�ol��p~��p4�6&��q5	V3.0}0�#m61c�$�*(��$1!6�A�� Eo�E���E��E���F��F�!�F8��FT��Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G,�IR�CH`�C��dTDU�?D���D��DE�(!/E\�E���E�h�E��ME��sF�`F+'\F�D��F`=F�}'�F��F��[
F���F���M;S@;Q�U�|8�`rz@/&�8�6&<��1��w�^$ESTPAR�S  *({ _#H�R��ABLE 1%�p+Z�6#|�Q�Q � 1�|�|�|��5'=!|�	|�
|��|�˕6!|�|�:|���RDI��z!ʟܟ� ��$���O������¯ԯ�����S��x# V���˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���U-����ĜP�9� K�]�o��-�?�Q�c��u���6�NUM  ��z!� �>  Ȑ����_CF�G �����!@�b IMEBF_T�T����x#��a�VE�R��b�w�a�R {1�p+
 (3�6"1 ��  6!�� �������� �9�$�:� H�Z�l�~���������@������^$��_���@x�
b MI_�CHANm� x� >kDBGLV;0o��x�a!n ETHE�RAD ?�
� �y�$"�\&�n ROUT��!�p*!*�SN�MASK�x#�255.h�fx�^$OOLOFS_�DI��[ՠ	OR�QCTRL � p+;/���/+/=/ O/a/s/�/�/�/�/�/���/�/�/!?��PE?_DETAI���PON_SVOF�F�33P_MON� �H�v�2-9S�TRTCHK ����42VTCOMPATa8�24�:0FPROG =%�%CA)&O~�3ISPLAY���L:_INST_M�P GL7YDUS8���?�2LCK�LPKQUICKMEt ��O�2SCRE�@}�
tps�@�2�A�@�I��@_Y����9�	SR_GR�P 1�� ���\�l_zZg_@�_�_�_�_�_�^�^� oj�Q'ODo/ohoSe ��oo�o�o�o�o�o �o!WE{i�������	1234567�h�!���X�E1�V[�
 �}ipn�l/a�gen.htmno��������ȏ�~�Panel� setup̌}��?��0�B�T�f� ��񏞟��ԟ� ��o����@�R�d�v� �����#�Я���� �*���ϯůr����� ����̿C��g��&� 8�J�\�n�����϶� ��������uϣϙ�F� X�j�|ߎߠ����;� ������0�B��*N�UALRMb@G ?�� [��� ���������� ��%� C�I�z�m�������v�SEV  �����t�ECFG CՁ=]/BaA$�   B�/D
 ��/C�Wi{� ������4 PRց; �To�\o�I�6?K0(%����0���� �//;/&/L/q/\/`�/�/�/l�D ��Q�/I_�@HIS�T 1ׁ9  �(  ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,153,1�?v?�?�?�?�� >?P=962c?�?
O`O.O�?�?�136�? |O�O�O�OAOSOeO�O __0_�HM___q_�_ �_�_�_H_�_�_oo %o7o�_[omoo�o�o �oDo�o�o�o!3E ��a81�ou� �����o��� )�;�M��q������� ��ˏZ�l���%�7� I�[���������ǟ ٟh����!�3�E�W� ���������ïկ� v���/�A�S�e�P b������ѿ����� �+�=�O�a�s�ϗ� �ϻ�������ߒ�'� 9�K�]�o߁�ߥ߷� �������ߎ�#�5�G� Y�k�}�������� �������1�C�U�g� y���v����������� 	�?Qcu� �(���� )�M_q��� 6���//%/� I/[/m//�/�/�/D/ �/�/�/?!?3?�/W? i?{?�?�?�?�����? �?OO/OAOD?eOwO �O�O�O�ONO`O�O_ _+_=_O_�Os_�_�_ �_�_�_\_�_oo'o 9oKo�_�_�o�o�o�o �o�ojo�o#5G Y�o}�������?��$UI_P�ANEDATA �1������  	�}�0�B�T�f�x��� )����mt�ۏ� ���#�5���Y�@�}� ��v�����ן����� ��1��U�g�N������ �1��Ïȯ گ����"�u�F��� X�|�������Ŀֿ=� �����0�T�;�x� _ϜϮϕ��Ϲ������,ߟ�M��j�o� �ߓߥ߷������`� �#�5�G�Y�k��ߏ� ������������� �C�*�g�y�`����� ����F�X�	-? Qc����߫�� ��~;"_ F��|���� �/�7/I/0/m/�� ���/�/�/�/�/�/P/ !?3?�W?i?{?�?�? �??�?�?�?O�?/O OSOeOLO�OpO�O�O �O�O�O_z/�/J?O_ a_s_�_�_�_�O�_@? �_oo'o9oKo�_oo �oho�o�o�o�o�o�o �o#
GY@}d ��&_8_���� 1�C��g��_������ ��ӏ���^���?� &�c�u�\�������ϟ ���ڟ�)��M�� ���������˯ݯ0� ����7�I�[�m�� ��������ٿ�ҿ� ��3�E�,�i�Pύϟ�����Ϫ���Z�l�}����1�C�U�g�yߋ�) ߰�#������� �� $�6��Z�A�~�e�w� �����������2� �V�h�O�����v�p���$UI_PAN�ELINK 1��v�  ��  ��}�1234567890����	-? G ���o���� �a��#5GD�	����p&���  R����� Z��$/6/H/Z/l/ ~//�/�/�/�/�/�/ �/
?2?D?V?h?z?? $?�?�?�?�?�?
O�? .O@OROdOvO�O O�O �O�O�O�O_�O�O<_�N_`_r_�_�_�0, ���_�X�_�_�_ o2o oVohoKo�ooo�o�o �o�o�o�o��, >r}������� �����/�A�S� e�w��������я� ��tv�z����=� O�a�s�������0S�� ӟ���	��-���Q� c�u�������:�ϯ� ���)���M�_�q� ��������H�ݿ�� �%�7�ƿ[�m�ϑ� �ϵ�D��������!� 3�Eߴ_i�{�
�߂� ���߸������/�� S�e�H���~��R~ '�'�a��:�L�^� p���������������  ��6HZl~ ���#�5���  2D��hz�� ���c�
//./ @/R/�v/�/�/�/�/ �/_/�/??*?<?N? `?�/�?�?�?�?�?�? m?OO&O8OJO\O�? �O�O�O�O�O�O�O[� _��4_F_)_j_|___ �_�_�_�_�_�_o�_ 0ooTofo��o��o ��o�o�o,> 1bt����K ����(�:��� �{O������ʏ܏� uO�$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v�������� п���ϕ�*�<�N� `�rτ��O�Ϻ�Io�� �������8�J�-�n� ��cߤ߇����߽��� �o1�oX��o|�� ������������ 0�B�T�f�������� ������S�e�w�,> Pbt��'�� ���:L^ p��#����  //$/�H/Z/l/~/ �/�/1/�/�/�/�/?  ?�/D?V?h?z?�?�? �???�?�?�?
OO.O ��ROdO�߈OkO�O�O �O�O�O�O_�O<_N_ 1_r_�_g_�_7O�M�m�$UI_Q�UICKMEN � ���_AobRESTO�RE 1��  � |��Rto�o�im�o�o �o�o�o:L^ p�%����� �o����Z�l�~� ����E�Ə؏����  �ÏD�V�h�z���7� ������/���
��.� @��d�v�������O� Я�����ßͯ7� I���m�������̿޿ ����&�8�J��n� �ϒϤ϶�a������� Y�"�4�F�X�j�ߎ� �߲������ߋ����0�B�T�gSCRE�`?#muw1sco`u2��U3��4��5��6���7��8��bUSE�Rq�v��Tp���k�s����4��5��6���7��8��`ND�O_CFG ܶ#k  n` `P�DATE ���Noneb�SEUFRAME�  �TA�n�R�TOL_ABRT8y�l��ENB����?GRP 1�ci/aCz  A��� ��Q�� $6H!Rd��`U����~��MSK  ��4���Nv�%�U��%���bVISCAND_MAX��I��FAI�L_IMG� �P��P#��IMRE/GNUM�
,[gSIZ�n`�A��,VONTMOiU��@����2��a��a�����FR:�\ � �MC:\�\LO�G�B@F� !��'/!+/O/�Uz? MCV�8#oUD1r&EX{+�S�PPO64�_��0'fn66PO��LIb�*��#V���,f@��'�/� =	�(S�ZV�.����'W�AI�/STAT' ����P@/�?��?�:$�?�?��2�DWP  ���P G@+b=���� H�O_JMPERR 1�#k�
  �2345?678901dF�� �O{O�O�O�O�O�O_ �O*__N_A_S_�_
� MLOWc>
 ��_TI�=�'�MPHASE � ��F��PSoHIFT�1 9�]@<�\�Do�U #oIo�oYoko�o�o�o �o�o�o�o6l CU�y���� � ��	�V�-�e2�����	VSFT]1�2	VM��� �5�1G� ���~%A�  B8̀̀�@ pكӁ˂1�у��z�ME@��?�{��!c>&%�JaM1��k�0�{ ��$`0TDINE#ND��\�O� �z����S��w��P����ϜRELE��Q��Y���\�_ACTIV��:�R�A ��e���e��:�RD� ���YBOX �9�د�6���02���190.0.��83��25�4��QF�	 ��X�j��1��robot��� ?  p�૿�5pc��̿������7�����-�f�ZWABC�����,]@ U��2ʿ�eϢωϛ� �Ͽ����� ���V�@=�z�a�s߰�E�Z��1�Ѧ