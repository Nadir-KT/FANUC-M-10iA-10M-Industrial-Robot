��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  "� �ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1�� H PCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $� � N�O�PS_SPI�_INDE��$��X�SCREE�N_NAME {�SIGN���� PK_F�IL	$THK�YMPANE� � 	$DUMM�Y � u3|4�|�RG_STR�1 � $T�ITP$I��1�{������5�6�7�8
�9�0��z�P����1�1��1 '1
'2"�S�BN_CFG1 � 8 $CN?V_JNT_* |�$DATA_C�MNT�!$FL�AGS�*CHE�CK�!�AT_C�ELLSETUP�  P $HOME_IO,�G�%�#MACR=O�"REPR�(-�DRUN� D|�3SM5H UTO�BACKU0 �� $ENAB���!EVIC�T]I � D� �DX!2ST� ?0B��#$INTERV�AL!2DISP_�UNIT!20_D�On6ERR�9FR�_F!2IN,G�RES�!0Q_<;3!4C_WA�471��8�W+0�$Y �$DB� 6COMW!2MO� H.o	 \rVE�1�$F�RA{$�O�UDcB]CTMP�1_FtE2}G1_��3�B�2�XD��#
 d $�CARD_EXI�ST4$FSS�B_TYP!AH�KBD_SNB�1A�GN Gn $�SLOT_NUM��APREV4D�EBU� g1G ;1_�EDIT1 �� 1G=� S<�0%$EP�O$OP�U0LETE_OK�B{US�P_CR�A�$;4AV� 0LACIw1�R�@k ܢ1$@MEN�@$D�V�Q`PvVAl{� BL� OU&R ,A�0�!� =B� LM_O�
e=R�"CAM_;1� xr$A�TTR4�@� AN�NN@5IMG_H�EIGH�AXcWI7DTH4VT� �U�U0F_ASPE�C�A$M�0EX�P�.@AX�f�C�F�D X $�GR� � S�!.@B�PNFLI�`�d� �UIRE 3T!GI�TCH+C�`N� S&�d_LZ`AC�"�`SEDp�dL� J�4S�0� <za�!p;�G0 � 
$WARNM�0f�!p�@� -s�pNST� �CORN�"a1FL{TR{uTRAT� �T}p  $ACCa1�p��|{�r�ORI�P�C�kRTf0_S~B\qHG,]I1 [ T�`4�"3I�pTYD�@*2 3`#@� �!,�B*HDDcJ* C�d�2_�3_�4_�5�_�6_�7_�8_�9�4? �CO�$ <� �o�o�hK3 1#`�O_Mc@AC t� � E#6NGPvABA� �c1�Q 8��`,��@nr1�� d�P�0e�]p� cvnpUP&Pb26h���p�"J�p_R�r�PBC��J�rĘߜJV�@U� B��s}�g1��"YtP_*0OFS�&R @� RO_�K8T��aIT�3T�N'OM_�0�1p�38W >��D �� Ќd@��hPV��mEX�p�� �0g0ۤ�p�r
�$TF�2C$MDM3i�TO�3�0U� ^F� ��Hw2JtC1(�Ez�g0#E�{"F�"F�40CPh@�a2 �@$�P�PU�3N)�ύRևAX�!DU���AI�3BUFp�F=�@1 |pp����pPIT� PP�M�M�y��}F�SIMQSI�"ܢVAڤT�\�?�w T�`(zM��P�B�qFACTb�@EW�P1��BTv?�MC�5 �$*1JB`p脎*1DEC��F��� �=�� �H0CHNS_EMP1�G$G��8��@_4��3�p|@P��3�TC c�(r/�0-sx��ܐ�� MBi��!����JR|� i�SEGFR���Iv �aR�TpN�C��PVF4>�bx &��f{u Jc!�Ja��� !28�ץ8�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb��Ӏq�۽�н����Lp�3�B���CRC�e�3CCp����c� �mcҞb�1J�cѿ�.�T���D$ICb�Cq��5r�ե��@v�'���E�V���zF��_��FR,pN��ܫ�?�84�0A�! �r�� �h�Ϩ��p�2�͕a�� �د"P	�Cx Ϗ��oH"27�!ARV�O`C�'$LG�pV�B�1�P��@�t�aA�0'�|�b+0Ro�� MEp`0"1 CRA 3 CAZV�g6p�O �#FCCb�`�`F�`K�8������ADI��a �A�bA'�.p��p�`�c�`S4PƑ�a�A�MP��-`Y�3P�M��]pUR��QUA1 � $@TITO1�/S@S�!����"0�D�BPXWO��B0!5�$SK���2�P�x q�!"�"�PR�� 
� =����!g# @q1$2�S$z���L�)$�/H���� %�/�$C�!9&?�$ENE�q.c'*?�Ú RE�p�2(H ��O��0#$L|3$$@�#�B[�;���FOs_D��ROSr��#������3RIG7GER�6PApS��>��ETURN�2�c�MR_8�TUw�\�0EWM��M�cGN�P���BLAH��<E���P��&$�P� �'P@�Q3�CkD{��DQ���4�1�1��FGO_AWA�Y�BMO�ѱQ#!��DCS_�)7  �PIS� I  gb {s�C��A��[ �B$�S��AbP�@r�EW-�TNTVճ�BV�Q[C�(c`�UW�r�P�J��P�$0��S�AFE���V_SV>�bEXCLU�砝nONL2��SY��*a&�OT�a'�HI_V�4��B����_ *P0� 9�_�z��p �TSG�� +nrr�@�6Acc*b��G�#@E�V�.iHb?fANNUNX$0.$fdID�U�2�SC@�`�i�a��jP�f��z��@I$2,O��$FibW$}�OT�9@�1 $DUMMYT��da��dn��� � �E- ` ͑HE4(sg�*b��SAB��SUFFI�W��@CA=��c5�g6r�!MS�W�E. 8Q�KE3YI5���TM�10s�qA�vIN���ї!���/ D��HOST_P!�rT��t�a��tn��tsp�pEMpӰV��� SBLc �ULI�0  p8	=ȳ�r�DTk0~�!1 � $S�>�ESAMPL��j� ۰f璱f���I�0��>[ $SUB�k��#0�C��T�r#a�SAVʅ��c���C�,�P�fP$n0E�w �YN_B#2 0&Q�DI{dlpO(��v9#$�R_I��� �ENC2_9S� 3  5�C߰�f�- �SpU�����!4�"g�޲�1T���5X�j`ȷg��0�0K�4�AaŔAVER�qĕ9g�gDSP�v��PC���r"��(���ƓVA�LUߗHE�ԕM�+�IPճ��OPP ��TH��֤��"P�S� �۰F��df�J� ���aC1+�6 H�bLL_DUs�~a3@{��3:���OTX"���s��r�0NOAUTO�!7�p$)�$�*�R�c4�(�C� 8��C, �""�L�� �8H *8�L H <6����c"�`,  `Ĭ�kª�q��q��Psq��~q��7��8���9��0����1��1�̺1ٺ1�1�1� �1�1�2(�2T����2̺2ٺ2�U2�2 �2�2ʕ3(�3��3��̺3�ٺ3�3�3 �3��3�4(�B'q���?��!9 <�9�&�z��I��1��׌M��QFE@'@� :� ,6��Q? ��@P?`$�5�9�E�@A�a�A� �;p$TP�$VARI:�Z���7UP2�P< ���TDe���K`Q�縡�!��BAC�"=# T�p��e$)_,�b8n�kp+ IFIG�kp�H  ��P���@|`�!>t ;E�4�sC�ST�D� D���c�<� 	 C��{��_���l����R  ���FORC�EUP?b��FLUS�`H�N>�F ��^�RD_CM�@E������� ��@vMP��REMr F�Q��1k@P���7Q
K4	NJ��5EFFۓ:�@I�N2Q��OVO�O{VA�	TROV���DTՀ�DTMX� ��@�
ے_P`H"p��CL��A_TpE�@�pK	_(�FY_T��v(��@%A;QD� �����`�!0tܑ0RQ��"�_�a����M�7�sCL�dρRIV'��{��EARۑIOFHPC�@����B�Bƅ�CM9@���R ��GCLF�e!DaYk(M�ap#5Tu�DG��� �%��FsSSD �s? P�a(�!�1���P_�!�(J�!1��E�3�!3�+=5�&�GRA��7��@��;�PW��OyNn��EBUG_S�D2H�P{�_E �A L�뀏���TERM`5B�i5?��ORI�#e0Ci5L��SM�_�P��e0Di5}���TA�9Ei5$Z ��UP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1젎4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ��E�p %B`�'EC����AR$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"�r�A��?���ERV��XQ�Y�� mG>@�BN��U\���R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`�0SMT6�G�3�GR��13�aPA�L@���`�q�uH �� ���TOC�A�`P	P�`$O�P����p�ѡ�`�0O��RE�`R�4C�AO�p낎Be��`R�Eu�h�A��eo$PWR�IMu��RR_�c��q=B �I&2H���p_A�DDR��H_LE�NG�B�q�q�q$�Rj��S�JڢSS��SKN��u\��u̳�uFٳSE�A�jrS��[MN�!K���0��b����OLX���p����`ACRO 3pJ�@��X�+��Q���6�OUP3�b_"�IX��a�a1��}� ������(��H��D���ٰ��氋�IO�2S�D�����<
�7�L $l��`�Y!_OFFr�P�RM_���aT�TP_+�H:�M (|pOBJ]"�p��[$��LE~Cd�>��N � ��֑�AB_�TqᶔSؙ`H�LVh�KR�"uHITCOU���BG�LO�q ���h�����`��`sSS� ���HW��#A:�Oڠ<`IN�CPU2VISIOW�͑��n��to��t�o�ٲ �IOLN.��P 8��R��p�$SLob P7UT_n�$p���P& ¢��Y F_AuS�"Q��$L������Q  U�0	P4Aa��^���ZPHY��0-��a��UOI �#R `�K����$�u�"pPpk�`��$�����Y�UJ5��S-���NE6WJO9GKG̲DIS���1Kp���#T (�uAqVF�+`�CTR�C�
�FLAG2�LG�dU ���؜�~13LG_SIZ�����b�4�a��a�FDl�I`�w� m�_�{0 a�^��cg���4������Ǝ���{0��� SC#H_���a7�N�d�VW���E�"����D4��UM�Aљ`LJ�n@�DAUf�EAU��p��d|�r�GH�bܢ0��BOO��WgL ?�6 IT㸰�y0�REC��S#CR ܓ�D
�\���MARGm�!��@զ ��d%�����S�����W���U� �JG=M[�MNCHJ���_FNKEY\�K��7PRG��UF��7Pn��FWD��HL��STP��V��=@��,�А�RS��HO`����C9T��b ��7�[�UL���6�(RD� �d���Gt��@PO���������MD�FOC�U��RGEX��TKUI��I��4� @�L�����P� ���`��P��NE��C�ANA��Bj�VA�ILI�CL !�UDCS_HII4��s"�O�(!�S��³S��a���BU�FF�!X�?PTH$m���v`��P�@��a�!Y�?Pp��j�3��`OS1Z�2Z3Z8�� Z � ��[aEȤ\��ȤIDX�dPSR�rO���zA�ST�L�R}�Y&�� /Y$E�C����K�&&z�� [ LQ��+00�	P�� �`#qdt
�U�dw<���?_ \ �`4Р��\��Ѩ#\0C4�]{ ��CLDPL�>�UTRQLI��d8ڰ�)�$FLG&�� �1�#�D���'B�LqD�%�$�%ORGڰ 5�2�PVŇVY8�s�T8�r�$}d^ ���$(6��$�%S�`T� ��B0�4�6RCLM�C�4]?o?�9세�M9I�p}d_ d=њ�RQ��DSTB�p� ;F�HH�AX�R JHdLE�XCESr1!BM!p�a`��/B�T8�B��`a�p=F_�A7Ji��KbOtH� K��db \Q���v$�MBC�LI|�)SREQUIR�R�a.\<o�AXDEBUZ�ALt M��c�b�{Ph����2ANDRф�`�`d;�2�ȺSDC��N�INl�K�x`��X� N&��aZ����UPST� �ezrLOC�RI,rp�EX<fA�p�n9A���`AQ��7f XY�OND�rMF,Łf�s"��`}%�e/� ���FX3@�IGG�� g ��t"��ܓs#N�s$R�a%��iL��h�L�v�@�DATA#?pE�%�tR��Y��Nh t $+MD`qI}�)nv� ytq�ytHP`�Pxu��<(�zsANSW)�yt(@��yuD+�)Yr��ܵ0o�i �@CU�w�V�p 09AARR2��j Du�{Q��~7Bd$CALIA@���G��2��RI�N��"�<E�NTE��Ck�r^�آ�]���_N�qlk���9��*����Bm��DIVFFDH�@���qnI�$V,��S�$��$Z�X�o��*����oH ?�$BELT�u!_ACCEL�.�~�=�IRC�� ����D�T�8�$PS�@�"L�@�r��#�^�S�Eы T�PAT!H3���I���3x�p�A_W��ڐ���2n�C��4�_MG��$DD��T���$FW�Rp9��I�4���DE7�PPAB�N��ROTSPE!E�[g�� J��[��C@4��@$US�E_+�VPi��S�YY���1 qYNr!@A�ǦOFF�qnǡMOU��NG����OL����INC �tMa6��HB��0HBENCS+�8q9Bp�X4�FDm�IN�Ix�0]��B��VE��#�>y�23_UP񕋳/LOWL���p� B���Du�9B#P`��x ���BCv�r�MO3SI��BMOU��@��7PERCH  ȳOV��â
ǝ� ���D�ScF�@MP����� Vݡ�@y�j��LUk��Gj�p�UPp=ó���ĶTRK�>�AYLOA�Qe� �A��x�����N`�F��RTI�A$��MO UІ�HB�BS0�p7D5����ë�Z�DU�M2ԓS_BCKLSH_Cx�k�� ��ϣ���=���ޡ< �	ACLAL"q�p�1м@��CHK� :�S�RTY���^�%E1Qq_�޴_�UM�@�C#��S�CL0�r�LMT_OJ1_L��9@H��qU�EO�p�b�_�e�k�e�SPC��u�L��N�PC�N�Hz �\P��C�0~"XT\��CN_:�N9�L�I�SF!�?�V����U�/���x�T���CB!�SH�:��E� E1T�T����y���T�f�PA ��_P��_� =������!����J6 L�@���OG�G�TORQU��ONֹ��E�R0��H�E�g_W2��ā_郅���I*�I�I��Ff`xaJ�1�~1�VC3�0BD:B�1�@SBJRKF9~�0DBL_SM�:�2M�P_DL2GRV�����fH_��d���CcOS���LNH ��������!*,�aZ���fcMY�_(�TH���)THET0��N�K23���"��C-B�&CB�CAA�B��"��!��!�&SB8� 2�%GTS�Ar�CIMa�����,4#<97#$DU���H�\1� �:Bk62�:AQ�(rSf$NE�D�`I ��B+5��$̀�!�A�%�5�7���LCPH�E�2���2S C%C%�2-&FC0JM&̀V�8V�8߀LUVJV!KV/KV=KUVKKVYKVgIH�8@FRM��#X!KH/KUH=KHKKHYKHgI�O�<O�8O�YNO�JO!KO/KO=KO*KKOYKOM&F�2�!�+i%0d�7SPBA?LANCE_o![c�LE0H_�%SP�c� &�b&�b&PFULC�h�b�g�b%�p�1k%�UTO_<��T1T2�i/�2N��"�{�t#�Ѡ�`�0�*�.�T��O�À<�v INSEG"�ͱREV4vͰl�gDIF�ŕ�1lzw6��1m��OBpq�ь�?�MI{���nL�CHWARY�_�A�B��!�$MEC�H�!o ��q�AX���P����7Ђ�`n� 
�d(�U�RO�B��CRr�H���8'�MSK_f`��p P �`_���R/�k�z�����1 S�~�|�z�{���z��q�INUq�MTC�OM_C� �q � ���pO�$ONOREn����p�Ђr 8p GRle�uSD�0AB��$XYZ_DAx�1a���DEBUUqX������s z`$��wCOD�� L����p�$BU�FINDX|� � <�MORm�t $فUA��֐�Ф�
y��rG��u� � $SIMUL  S�*�Y�̑a��OBJE�`̖AD�JUS�ݐAY_	IS�D�3���_FI�=��T u 7�~�6�'��p} =��C�}p�@b�D��FRiIr��T��RO@ �\�E}��y�OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1�0e��M��ED}�*�p ��N�PMֲ���&c�w�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B��2�G�B�_�M�� �q�E� �x Hw��p��AT+USW���C�0o��s���BTM�ǌ�I
�k�4��x�԰q�y Dw�E&���@E�r��7��жЗ�EXE��ἱ���8��f q�z @w���3UP'��$�pQ�XN����������� �PG΅{ h? $SUB�����0_���!�MPW�AIv�P7ã�LO�R���F\p˕$R�CVFAIL_C���BWD΁�v��DEFSP!p | Lw���Я�\���UNI+�����bH�R�+�}_L\pAP��x�t���p�}H��> �*�j�(�s`~�NN�`KETB�%�J�PE Ѓ~��J0SIZE����X�'����S�OR��FORMAT�`��c ��WrEM�t��%�UqX��G��PLI��~p�  $ˀP_SWI�pq�J�_PL��AL_ S�����A��B���� C��D�$E���.�C_�U��� � � ���*�J3K0�����TIA4��5��6��MOM������h���ˀB��AD����������PU� NR��������m��� A$PI�6q��	���� �K4�)6�U��w`���SPEEDgPG ��������Ի�4 T�� � @��SAMr`��\�]��MOV_�_$�np t5��5���1���2��������'�S�Hp�IN�'�@ �+����4($4+T+GAMMWf�1'�$GET`�p����Da���

pLIB�R>�II2�$HIB=�_g�t��2�&E;�b�(A�.� �&LW�- 6<�)56�&]��v�p���V��$PGDCK���q��_?�����q�&���7��4���9+� �$IM_SR�p�D�s�rF��r�rLE����Om0H]��0�p���pq��PJq?UR_SCRN�FA����S_SAVEc_D��dE@�NOa�CAA�b�d@�$q�Z �Iǡs	�I� �J�K�  ����H�L��>�" hq������ɢ� � bW^US�A�u�
�M4���a��)q `��3�WW�I@v�_�q��.MUAo�� � �$PY+�$W�P�vNG�{��P�:��RA��RH��RO�PL�����q� ��s'�%X;�OI�&�Zxe ���m�� p��ˀ�3s�O�O�O�O�O�a:a�_т� |��q� d@��.v��.v��d@��[wFv��E���%s�tJ;B�w�|�tP���PMA�QUa ���Q8��1�Q�TH�HOLG�Q7HYS��ES��q�UE�pZB��Oτ�  ـPܐ(�A��(��v�!�t�O`�q���u�"���FA��IR#OG�����Q2����o�"��p��INF�Oҁ�׃V����R�vH�OI��� (�0SLEQ������ Y�3����Á��P0QOw0���!E0sNU��AUT�A�COPY�=�/�'��@Mg�N��=�}1h������ ��RG���Á���X_�P��$;ख�`��W��P���@�������EX_T_CYC b�Qȝ�RpÁ�r��_N�Ae!А���R�Ov`	�� � 9���POR_�1�\E2�SRV �)_�6I�DI��T_�k��}�'���dЇ�����5*��6��7��8i�H�iSdB���2�$��)F�p��GPLeAdA
�TAR�Б@����P�2�裔d� �,�0FL`�o@Y�N��K�M��Ck��GPWR+�9ᘐ��ODELA}�dY�p�AD�a��QSwKIP4� �A�Z$�OB`NT�} ��P_$�M�ƷF@\b Ipݷ�ݷ�ݷd�� ��빸��Š�Ҡ��ߠ�9��J2R�� ��� 4V�EX� TQQ����TQ������� ��`�H�RD�C�V� �`��X)�R�p�����r��~m$RGEAR_� sIOBT�2FLG��LfipER�DTC����Ԍ���2TH2N�S}� 1� ���G T\0 I���u�M\Ѫ`I�\d"�REF�1Á� l�h��ENA9B��cTPE�04� ]����Y�]��ъQn#���*��"���ҡ���2�Қ�߼��������
�3�қ'�9�K�]�(o���4�Ҝ������������5�ҝ�!�3�E�W�i�{��6�Ҟ������������
�7�ҟ-?Q(cu�8�Ҡ�������SMSKÁ� �p�0���EkA��EMO[TE6�����@0�݂TQ�IO}5��ISTP�POW@��� �pJ���������E�"$�DSB_SIGN�1UQ�x�C\�TP����RS232����R�iDEVICE�US�XRSRPAR�IT��4!OPBI�T�QI�OWCONTR+�TQ��?SR�CU� MpSUXTASK�3N�p�0p$oTATU�P�IS�0�����p_XP�C)�$FREEFROMS	pna��GET�0��UPD2�A�2��SP� :�ߧ� !$USAN�na&�����ERI�0�RpRY$q5*"_j@�Pm1�!N�6WRK9KD����6��QFRIEND�Q�RUFg�҃�0oTOOL�6MY�t�$LENGTHw_VT\�FIR�p�C�@ˀE> +IUF�IN-RM��RGyI�1ÐAITI�b$GXñ3IvFG2v7�G1���p3�B�GP1R�p�1F�O_n 0��!RE��p�53҅�U�TC��3A�A�F ��G(��":��� e1n!��J�8�%���%�]��%�� 74�XS O0�L��T�3�H&��8���%b453G�E�W�0�WsR�TD ����T��M����Q�T�]�$V 2�����1�а91�8�02*�;2k3�;3�:i fa�9-i�aQ��NS���ZR$V��2BVwEVD�2AQ�B;�����&�S�`��F�"�kX�@�2a�PS�E���$r1C��_$Aܠ6wPR��7vMUb�cS�t '�F"619�� 0G�aV`��p�d`���50�@ԍ�-�
25S��� ��aRW����4B�&�N�AX�!��A:@LAh��rTHIC�1I���X�d1�TFEj��q�uIF'_CH�3�qI܇7�Q�pG1RxV���]�t�:�u�_JF~��PRԀƱ�RVA=T��� ��`����0RҦ�DOfE��CsOUԱ��AXI���OFFSE׆TRIGNS���c����h�����H�Y�䓏IGMA0PA�p�J�E�ORG_UNsEV�J� �S��~���d �$C�z��J�GROU��Ɖ�TOށ�!��DSP��JOGӐ�#��_Pӱ�"O�q�����@�&KEP�IRȼ�ܔ�@M}R��AP��Q^�Eh0��K�ScYS�q"K�PG2�BRK�B��߄�p�Y�=�d����`ADx_�����BSOC����N��DUMMY�14�p@SV�PD�E_OP�#SFS�PD_OVR-�b��C��ˢΓOR٧3N]0ڦF�ڦ��OV��SF��p���F+�r!���CC��1�q"LCHDL��R�ECOVʤc0��Wbq@M������RO�#䜡Ȑ_+��� @�0�e@VER�$7OFSe@CV/ �2WD�}��Z2����TR�!���E�_FDO�MB_�CM���B��BL �bܒ#��adtVQRҐ$0p���G$�7�A�M5��� eŤ��_�M;��"'����8$�CA��'�E�8�8$�HBK(1���IO�<�����QPPA ������
��Ŋ����?DVC_DBhC;�@�#"<Ѝ�r!S�1[���S�3[֪�ATIEOq 1q� ʡU�3���CABŐ�2�C@vP��9P^�B���_� ~�SUBCPU�ƐS�P �M�)0NS��cM�"r�$HW_C��U��S@��S�A�A�pl$UNI5Tm�l_�AT����e�ƐCYCLq�N�ECA���FLT?R_2_FIO�7(��)&B�LPқ/�.�o_SCT�CF_`�aFb�l���|�FS(!E�e�CHA�1��4�8D°"3�RSD��$"�}����_Tb�PcRO����� EMi�_��a�8!�a 1!�a��DIR0�?RAILACI�)RMr�LO��C���Q�q��#q�դ�PRJ=�S�AC/�zc 	��FUNCq�0rRINP�Q�0���2�!RAC �B ��[���[WAR�n���BL�Aq�A0����DAk�\���LD0���Q���qeq�TI�"r��K�hPRIA,�!r"AF��Pz!=��;��?,`�RK���MrǀI�!�DF_@�B�%1n�LM�FA�q@HRDY�4_�P�@RS�A�0� �MULSE@���a� ��ưt���m�$�1$�1�$1o����7� x*�EGE �����!AR���Ӧ�0�9�2,%� 7�AXE.��ROB��WpA��_l-��SY[�W!‚�&S�'WRU�/-1��@�STR�����:�Eb� 	�%��J��AB� ���&9���֐�OTo0 	$��ARY�s#2��Ԛ��	ёFI@��$LINK|�qC1%�a_�#���%kqj2XYZ��t;rqH�3�C1j2^8'0	B��'�4����+ �3FI���7�q����'��_Jˑ���O3N�QOP_�$;5��F�ATBA�QBC��&�DUβ�&6��TURN߁"r�E11:�p��9GFL�`_��Ӑ* �@�5�*7��Ʊ W1�� KŐM���&8���"r��ORQ��a�(@#p =�j�g�#qXU�����NmTOVEtQ:�M���i���U��U��VW �Z�A�Wb��T{�, �� @;�uQ���P\�i��U�uQ�We�e�SE)Rʑe	��E� O���UdAas��4S�0/7����AX��B �'q��E1�e��i� �irp�jJ@�j�@�j�@ �jP�j@ �j�!�f� �i��i��i��i� �i�y�y�'y�x7yTqHyDEBU8�$32���qͲf2G + AB����رrnSVS�7� 
#� d��L�#�L��1W��1 W�JAW��AW��AW�Q�W�@!E@?D2�3LAB�29U4�Aӏ�ޮC  o�ER|f�5� � $�@�_ A��!�PO���à�0#�
�_M�RAt�� d r� T��ٔERR��L��;TY&���I��qV�0�cz�TOQ�d�PL[ �d�"�� ?�|w�! � pp`qT)0���_V1VrP�aӔ����2ٛ2薈E����@�H�E����$W�����V!��$�P��o�cI���aΣ	 HELL�_CFG!�� 5��B_BAS�q�SR3��� Ea#Sb���1�U%��2��3��4��U5��6��7��8����RO����I0�0NL�\CAB+�����ACK4�����,�\@p2@�&�?�_PUﳳCO. U�OUG�P�~ ����m�������T=Pհ_KAR�l�&_�RE*��P���|�QUE���uP�����CSTOPI_AL7�l�k0��h��]�l0SEM�4�(��M4�6�TYN�SO���DIZ�~�A������m_TM�MA'NRQ��k0E�����$KEYSWI�TCH���m���H=E��BEAT��|�E- LE~�����U±�F!Ĳ���B�O_�HOM=OGREFUPPR&��y!� �[�C��O��-EC�OC��Ԯ0_IOC�MWD
�a�'8k��� � Dh1���UX���M�βgP�gCFORC��� �	�m�OM.  �� @�5(�U��#P, 1��, 3���45	�NPXw_ASt�� 0���ADD���$S�IZ��$VAR\���TIP/�.�
�A�ҹM�ǐ��/�H1�+ U"S�U!Cz����FRIF��J�S0���5Ԓ�NF��܍� � xp`SIƗ�TE�C���CSG%L��TQ2�@&���x�� ��STMT��2,�P �&BWuP���SHOW4���S�V�$�� �Q�A00�@Ma}����� �����&���5���6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G�� 0G���0G���@GP��PG��1	1	U1	1+	18	1E	U2��2��2��2��U2��2��2��2��U2��2��2	2	U2	2+	28	2E	U3��3��3��3��U3��3��3��3��U3��3��3	3	U3	3+	38	3E	U4�4��4��4��U4��4��4��4��U4��4��4	4	U4	4+	48	4E	U5�5��5��5��U5��5��5��5��U5��5��5	5	U5	5+	58	5E	U6�6��6��6��U6��6��6��6��U6��6��6	6	U6	6+	68	6E	U7�7��7��7��U7��7��7��7��U7��7��7	7	U7	7+	78	7Ev��VP��UPDs��  �`NЦ��
��YSLOt�� � L��d���A�aTA�0d��|��ALU:ed�~�CU�ѰjgF!aID_L��ÑeHI�jI��$FILE_���d��c$2�
�cSA>�� hO��`E_B�LCK��b$��hD_CPUyM�yA���c�o�d�b����R ;�Đ
PW��!�[ oqLA��S=�8ts�q~tRUN�q st�q~t���qst�q�~t �T��ACC�s��X -$�qLEN;��tH��p�h�_�I��ǀLOWo_AXI�F1�q
�d2*�MZ���ă���W�Im�ւ�aR�TOR��pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v�������TCV��؁��T��ي�����t�V�H���V�Jj�R�MA�"��J��m�u�b����q2j�#�U�{�t�6K�JK��VK;���4H���3��J0�����JJ��JJ��AAAL��ڐ��ڐԖ4Օ5���N1���ʋƀW�LP�_(�g��Ѽ�pr�� `�`GGROUw`��B�ПNFLIC��f�R�EQUIRE3�E�BU��qB���w�2�����p���q5�p��� \��APPRҒ�C}�Y�
ްEN�٨CLO7��S_!M��H���u�
�qu�o� ���MC��8���9�_MG��C��Co��`M�в�N�B;RKL�NOL|�N�:[�R��_LINђ�$|�=�J����Pܔ�� ���������������6ɵ�̲8k�C����� ��
��q�)��7�PATH 3�L�B�L��H�wࡠm�J�CN�CA��ؒ�ڢB�IN�rUChV�4a��C!�UM��!Y,���aE�p�����ʴ���PAYL�OA��J2L`R'_AN�q�Lpp����$�M�R_F2�LSHR��N�LO�ԡ�Rׯ�`ׯ�ACRL_G�ŒЛ� �r�Hj`߂$HM�^��FLEXܣ�q}J�u� :� ������������1�F1�V�j�@�@R�d�v�������E�� ��ȏڏ����"�4� q���6�M���~��U��g�y�ယT��o�X ��H������藕?� ����ǟِݕ�ԕ�����%�7���J�� � V�h�z����`AT�採@�EL��� S��J|��v��JEy�CTR���~�TN��FQ��H�AND_VB-����v`�� $��Fa2M����ebSW���q'��� $$	MF�:�Rg�(x�,4�%��0&A�`�=���aM)F�AW�Z`i�A�w�A��X X�'pi�D*w�D��Pf�G�p�)CSTk��!x��!N��DY�pנM�9$`%� ��H��H�c�׎���0� ��Pѵڵ�쵠�������J��� ���1��R�6���QASYMvř����v��J���cі�_SH>��ǺĤ�ED� ���������J�İ�%��C�IDِ�_VI�!X�2PV_UCNIX�FThP�J�� _R�5_Rc�cTz�pT�V ��@���İ�߷��U I�������Hqpfˢ��aEN��3�DI����O4d8D�`J�� x g"IJAAȱz�aabp�c�oc�`a�pdq�a� ���OMME��м �b�RqT(`PT@�@� S��a7�;�Ƞ��@�h�a�iT�@<�� $DUMMY}9Q�$PS_���RFC�  S�v� �p���Pa� �XƠ���STE�SBRY�M21�_VF�8$SV_�ERF�O��LsdsC+LRJtA��Odb`�O�p � D $GLOBj�_LO���u�q�cAp��r�@aSYS�qA�DR``�`TCH>  � ,��ɩ�b�W_NA����7�A�SR���l ���
* ?�&Q�0"?�;'?�I) ?�Y)��X���h���x� �����)��Ռ�Ӷ�;� �Ív�?��O�O�O�D>D�XSCRE栘p5����ST��s#}y`����/u_HA�q� TơgpTYP�b���PG�aG���Od0�IS_䓀d�UEMd� ����ppyS�qaRSM_�q�*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCO�U��S�Ԕ 1�!�UE&��Ubwr���PROGM�FL�@$CUgpPO��Q��� UI_�`H>� � 8�� �_HE�PS�#��`?RY ?�qp�b���dp5��OU}S�� � @6p~�v$BUTTp��RpR�COLUMxq�e��SERV5��PANEH�q�� � �@GEU���Fy��)$H�ELPõ)BETERv�)ෆ���A� � � ��0��0�L�0ҰIN簪c�@QN��IH�1���_� ֪�LNN�r� �qpձ_ò�=�$H��TEqXl����FLA@^��RELV��D`���������M��?�,�ű�m����"��USRVIEWN�q� <6p�`U�`��NFI@;�F�OCU��;�PRI�� m�`�QY�TR�IP�qm�UN<`Md� #@p�*e�WARN)e6�SRWTOL%��g��Ẵ�ONCORN��R�AU����T���w��VIN�Le� {$גPATH9��גCACH��LO9G�!�LIMKR�����v���HOSTN�!�b�R���OBOT�d�IM>� �� ����Zq�Zq;�VCPU?_AVAIL�!�+EX	�!AN����q��1r��1r��1 ��ѡ�p�  #`C�����@$TOO�L�$��_JMP�� ���e$�SS����SHI9F��Nc�P�`ג��E�ȐR����OS�UR��Wk`RADILѮ��_�a��:�`9a��`a�r��LULQ�$OUTPUTg_BM����IM��AB �@�rTILNSCO��C7� ������&�� 3��A���q����m�I�2G�n�y@Md��}��yDJU��N_�WAIT֖�}Ҵ�{�%! NE�u��YBO�� ��� $`�t�S�B@TPE��NE�Cp�J^FY�nB_T��R�І�a$�H[YĭcB��dM� ��F� �p�$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"g�"��[���P?���U�ZABC~%��  $�"�R��
�p�$$C�LAS�������!pϐ� � VI�RT]��/ 0ABS�����1 5�� < �!F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZi{0�-�AXL�p��"�n63  �{tIN��qztPRE�����v��p�uLARMRECOV 9l�rwtNG�� .;	 A   �|.�0PPLIC���?5�p��Handlin�gTool o� �
V7.50P�/23-�  �P�f��
��_S�Wt� UP�!�� x�F0��t���A�ϐv� 86m4�� �it	���{� r2 �7DA5�� ��� Qfy@��o�Noneis�ͅ˰ ��T����!LAe+x>�_l�V�uT�:�s9�UTO�"����t�y��HGAPO�N
0g�1��Uh�D� 1581�����̟ޟry����Q 1���p� ,�蘦��ր;�@��q�_��"�" �3c�.�H����D�HTTHKY X��"�-�?�Q���ɯ ۯ5����#�A�G�Y� k�}�������ſ׿1� ����=�C�U�g�y� �ϝϯ�����-���	� �9�?�Q�c�u߇ߙ� �߽���)�����5� ;�M�_�q����� ��%�����1�7�I� [�m����������! ����-3EWi {������ )/ASew� ���/��/%/ +/=/O/a/s/�/�/�/ �/?�/�/?!?'?9? K?]?o?�?�?�?�?O��?�?�?O#O]���T�O�E�W�DO_C�LEAN��7��CN�M  � ��__/_A_S_�D?SPDRYR�O��HIc��M@�O�_�_ �_�_oo+o=oOoao�so�o�o���pB��v �u���aX�t����|��9�PLUGG����G��U�PRCvPB��@��_�orOxr_7�SEGF}�K[mwxq�O�O������?rqLAP �_�~q�[�m������ ��Ǐُ����!�3�>x�TOTAL�f y�x�USENU�p©� �H���B��RG�_STRING �1u�
��Mn�S5�
ȑ_�ITEM1Җ  n5�� ��$�6�H� Z�l�~�������Ưد����� �2�D��I/O SIGN�AL̕Try�out Mode�ӕInp��Simulatedב�Out��O�VERR�P = �100֒In �cycl��בP�rog Abor���ב��Stat�usՓ	Hear�tbeatїM?H Faul��Aler'�W�E�W� i�{ύϟϱ������� �CΛ�A���� 8�J�\�n߀ߒߤ߶� ���������"�4�F�pX�j�|���WOR{p Λ��(ߎ����� �� $�6�H�Z�l�~����� ���������� 2PƠ�X ��A {������� /ASew������SDEV [�o�#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y?PALTݠ1�� z?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O��O�O�O_�?GRI �`ΛDQ�?_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|�� �������0�xB�T��oPREG�> �� f���Ə؏��� � �2�D�V�h�z��������ԟ���Z���$ARG_��D �?	���;���  w	$Z�	[O��]O��Z�p�.�SB�N_CONFIG� ;��������CII_SAV/E  Z������.�TCELLSE�TUP ;�%�HOME_IO�Z�Z�%MOV_8��
�REP�lU��(�UTOBACK�ܠ��F�RA:\z� X\�z�Ǡ'`�z����ǡi�INI�0�z���n�MESSAG���ǡC���ODE_D�������%�O�4�n�PAU�SX!�;� ((O>��ϞˈϾ� �����������*� `�N߄�rߨ߶�g�l ?TSK  wͥ�<_�q�UPDT+���d!�A�WSM_kCF��;���|'�-�GRP 2:�V?� N�BŰA�߾%�XSCRD1�1�
7� �ĥĢ ����������*��� ����r����������� 7���[�&8J\�n��*�t�GRO�UN�UϩUP_kNA�:�	t�n�_ED�17��
 �%-BCKEDT-�2�'LK�`���-t��z�q�q�z���2t1������q�k�(/��ED3/��/�.a/8�/;/M/ED4�/t/�)?�/.?p?�/�/ED5`??�?<?.�?8O�?�?ED6O�?�qO�?.MO�O'O9OED7�O`O_�O.�O8\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o�_�	-9o�oo%oCR _ 9]�oF�o��k� � NO_DE�L��GE_UN�USE��LAL_OUT �����WD_ABO�Rﰨ~��pITR�_RTN��|N'ONSk���˥�CAM_PARA�M 1;�!�
 �8
SONY �XC-56 234567890� ਡ@����?��( АP\�
���{����^��HR5q�̹��ŏR�57ڏ�Aff���KOWA S_C310M
�x�}̆�d @<� 
���e�^��П\ ����*�<��`�r��g�CE_RIA_UI�!�=�F��}�z� ��_�LIU�]���ꋐ<��FB�GP ]1��Ǯ��M�_�q�0�C*  �����C1��9��@Ҩ�G���CR�C]���d��l��s��R������[Դm��vꨰ������� +C����(������=�HE�`ONFI�ǰ�B�G_PRI 1�{V���� �ϨϺ����������CHKPAUS��w 1K� ,!u D�V�@�z�dߞ߈ߚ� �߾������.��R��<�b���O��x������_MOR��� �^Biqy-���� 	 �� ���*��N�`����"���?��q?;�;�I���K��9�P����ça�- :���	�

��M����pU�ð��<��,,~��DB���튒�)
mc:cpm�idbg�f�:��������¥�p��/�  �$���pH�� ��s>��p��p�0U�?�8�R��Ug�/������Uf�M/w�O/�
D�EF l��s)��< buf.t�xts/�t/��ާ��)�	`�����=�L���*MC��1�����?43��1���t�īCz � BHH�CPUe�B�_B�y�;��>C����CnY
K�E?�{hD]^Dٿ�?r���1D���^�=G	���F��F���Cm	fF�O�OF�ΫY	���&�w�1���s�J��.�p��ዐ�BDLw�M@x8��1Ҩ�����g@D�p@�0E�Y�1X�E�Q�EJP F��E�F� G��:F^F E��� FB� H�,- Ge��H�3Y��:�  >�33 ���N~  n8�~@��#5Y�E>�ðA��Yo<#�
"Q ����+_�'RSMOF�S�p�.��'T1>��DE ��F� 
Q��;�(P � B_<_��R��X��	op6C4P�Y
�s@ ]AQ�2s@CR�0B3�MaC{@@*c�w��UT�pFPROG %�z�o�o�igI�q���v��ldK�EY_TBL  ��&S�#� �	
��� !"#�$%&'()*+�,-./01i�:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������vq���͓���������������������������������耇���������������������p`LCK�l4�p`�`�STAT ��S_A�UTO_DO����5�INDT_ENB!���R�Q?�1��T2}�^�STOP�b���TRLr`LE�TE��Ċ_SCREEN �Z�kcsc��U���MMENU 1� �Y  < �l�oR�Y1�[���v� m���̟�����ٟ� 8��!�G���W�i��� �����ïկ��4�� �j�A�S���w����� 迿�ѿ����T�+� =�cϜ�sυ��ϩϻ� ������P�'�9߆� ]�o߼ߓߥ������ ��:��#�p�G�Y�� ����������$��� �3�l�C�U���y��� �������� ��	V�Y)�_MANUA�P���$DBCO�[�RIGڇ
�DB'NUM� ��B1 e�
�PXWORK 1!�[�_�U/4FX�_AW�AY�i�GCP�  b=�Pj_AL� #�j�Y��܅ `��_�  1"�[/ , 
�odP�&/~&lMZ�IdP�x@P@#ONTImMه� d�`&�
�e�MOTN�END�o�REC�ORD 1(�[8g2�/{�O��!�/ ky"?4?F?X?�(`? �?�/�??�?�?�?�? �?)O�?MO�?qO�O�O �OBO�O:O�O^O_%_ 7_I_�Om_�O�_ _�_ �_�_�_Z_o~_3o�_ Woio{o�o�_�o o�o Do�o/�oS�o L�o����@� ��+�yV,�c�u� �������Ϗ>�P�� ���;�&���q���� ����P�ȟ�^���� ��I�[����� ����$�6�������jTOLERENCwsB���L�͖ �CS_CFG �)�/'dMC�:\U�L%04dO.CSV�� c���/#A ��CH��z� //.ɿ��(S��RC_OUT �*���SGN� +��"��#��10-FEB-�20 18:23~015-JANp��0:51+ P/Vt�ɞ�/.���f�pa�m���PJPѲ��V�ERSION �Y�V2.0�.84,EFLOG�IC 1,� 	:ޠ=�ޠL���PROG_ENqB��"p�ULSk'� ����_WRS�TJNK ��"fE�MO_OPT_S�L ?	�#
 	R575/# =�����0�B����TO  �ݵϗ��V_F EX�d��%��PATH ;AY�A\����\�5+ICT�Fu�-�j�#�egS�,�STBF_TTS�(�	d����l#!w�� MAqU��z�^"MSWX��.��4,#�Y�/�
!J�6%Z�I~m��$SBL__FAUL(�0�^9'TDIA[�1<��� ���1�234567890
��P��HZ l~������ �/ /2/D/V/h/�Z� P� ѩ� yƽ/��6�/�/�/? ?/?A?S?e?w?�?�?��?�?�?�?�?�,/�U3MP���� �A�TR���1OC@PM�El�OOY_TEM=P?�È�3F���G�|DUNI��.�Y�N_BRK 2�_�/�EMGDI_�STA��]��ENC�2_SCR 3�K7(_:_L_^_l& _�_�_�_�_)��C�A14_�/oo/oAo�Ԣ�B�T5�K� ϋo~ol�{_�o�o�o '9K]o� �������� #�5��/V�h�z��л` ~�����ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T���x��������� ү�����,�>�P� b�t���������ο� ���(�f�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������:� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ���*<N` r������� &8J\n� ���������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?��?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O��O__NoETMO�DE 16�5��Q �d�X
�X_j_|Q�PRROR�_PROG %fGZ%�@��_  �U�TABLE  �G[�?oo)oRjR�RSEV_NUM�  �`WP��QQY`�Q_AUT�O_ENB  ��eOS�T_NOna �7G[�QXb W *��`��`��`	��`d`+�`�o�o�o�dHISUc�QOP�k_ALM 18G[� �A��l�P+�ok}����r�o_Nb�`  G[��a�R
�:PTCP_VER !GZ�!�_�$EXTL�OG_REQv9�i\�SIZe�W��TOL  �QD�zr�A W�_BWD�p��xf́t�w_DI�� 9�5��d�T�QsRֆS�TEP��:P�O/P_DOv�f�P�FACTORY_�TUNwdM�EATURE :�5�̀rQHa�ndlingTo�ol �� \sf�mEngli�sh Dicti�onary��ro�duAA V�is�� Mast�er����
EN�̐nalog I�/O����g.fd�̐uto Sof�tware Up�date  F �OR�matic Backup���H596,�g�round Ed�itޒ  1 H�5Camer�a�F��OPLG�X�ell𜩐II�) X�ommՐs�hw���com��c9o���\tp����pane��  o�pl��tyle �select��a�l C��nJ�Ցo�nitor��RD�E��tr��ReOliab𠧒6U�Diagnos(��푥�5528�u���heck Sa�fety UIF���Enhance�d Rob Se�rv%�q ) "�S�r�User F�r[�����a��xt�. DIO �f�iG� sŢ��en]dx�Err�LF�� pȐĳr됮� ܻ���  !��FCTN Menu`��v-�ݡ���TP �Inېfac� � ER JG�C�pבk Exczt�g��H558��igh-Spex��Ski1�  2�
P��?���mmuwnic'�ons���&�l�ur�ې��S�T Ǡ��con�n��2��TXPL��ncr�str�u����"FAT�KAREL C�md. LE�ua�G�545\��Ru�n-Ti��Env��d
!���ؠu++�s)�S/W���[�Licen3seZ��� 4T�0��ogBook(S�yڐm)��H54�O�MACROs,~\�/Offse��7Loa�MH�������r, k�Mec�hStop Pr�ot���� lic�/�MiвShif8����ɒMixx���)���xStS�Mo�de Switc�h�� R5W�Mo��:�.�� 74 H���g��K�2h�?ulti-T=�M����LN (P{os�Regiڑ�������d�ݐt Fun�ǩ�.������Num~����� l�ne��ᝰ Ad�jup�����  �- W��tatu�w᧒T�RD�Mz�ot��sco+ve U�9����3Ѓ�uest 492�*�o������62;�SNPX yb ���8 J7`���Libr��J�48���ӗ� �Ԅ�
��6O�� Part�s in VCCMt�32���	�{�ޤ�J990��/I�� 2 P��TM/ILIB��H���P�AccD�L�7
TE$TX�ۨ�7ap1S�Te����pkey��wգ��d��Unex�ceptx�mot�nZ���������є�� O���� �90J�єSP CSXC<�f��Ҟ�� Py�We}���P3RI�>vr�t��men�� ��iPɰa�����v�Grid�pla�y��v��0�)�H1��M-10iA(_B201 �2\�� 0\k/�Ascii�l�Т�ɐ/��Col��ԑGuaMr� 
�� /P-��ޠ"K��st{P�at ��!S�Cyqc�҂�orie�v�IF8�ata- quҐ�� ƶ��moH574��RL���am���Pb�HM/I De3�(b����PCϺ�Pas�swo+!��"PE�? Sp$�[���tp\��� ven��Tw��N�p�YELLO�W BOE	k$Ar�c��vis��3�*�n0WeldW�cGial�7�V#tѓOp����1y� �2F�a�portN�(�p�T1�T� ��� ��xy]�&T5X��tw�igj�1�� b� ct\�J�PN ARCPS�U PR��oݲO�L� Sup�2fi�l� &PAɰאcr=o�� "PM(�����O$SS� eвtex�� r���=�=t�ssagT��	P��P@�Ȱ�锱�rtW��H'>r��dpn��n1
�t�!� z ��as�cbin4psy�n��+Aj�M H�EL�NCL V�IS PKGS �PLOA`�MB ��,�4VW�RI�PE GET_V�AR FIE 3�\t��FL[�OO�L: ADD R�729.FD \Kj8'�CsQ�QE���DVvQ�sQNO �WTWTE��}PD�  �^��biRFwOR ��ECTn��`��ALSE A�LAfPCPMO-�130  M" �#h�D: HAN?G FROMmP��AQfr��R709� DRAM AV�AILCHECK�SO!��sQVPCS� SU�@LIMC�HK Q +P~dFF� POS��F�Q �R5938-12 CHARY��0�PROGRA �W�SAVEN`A�ME�P.SV��7��$En*��p?FU��{�TRC|� SH�ADV0UPDAT� KCJўRSTA�TI�`�P MUC�H y�1��IMQ� MOTN-00�3��}�ROBOG�UIDE DAU�GH�a���*�toQu����I� Šhd��ATH�PepMOV�ET�ǔVMXP�ACK MAY ?ASSERT�D���YCLfqTA�rB�E COR vr�*Q3rAN�pRC OPTIONSJ1�vr̐PSH-1k71Z@x�tcǠSU1�1Hp^9R!�Q�`C_T�P��'�j��d{tby app wa 5I�~d�P�HI���p�aTEL��MXSPD TIB5bLu 1��UB6@��qENJ`CE2�6�1��p��s	�ma�y n�0� R6�{�R� �Rtraf�f)�� 40*�p���fr��sysv�ar scr Jq7��cj`DJU���bH V��Q/�PS?ET ERR`J`� 68��PNDA�NT SCREEN UNREA��4'�J`D�pPA���p=R`IO 1���P�FI�pB�pGROUN�PD��G��R�P|�QnRSVIP !p��a�PDIGIT �VERS�r}BLo��UEWϕ P06s  �!��MAGp0�abZV�DI�`� SSUE�ܰ��EPLAN JO�T` DEL�pݡ#�Z�@D͐CALLOb�Q ph��R�Q�IPND��IMGޏR719��MN�T/�PES �pV:L�c��Hol�0Cq����tPG:�`C�M��canΠ��pg�.v�S: 3D �mK�view d2�` �p��ea7У�b� of �Py����ANNOT AC?CESS M��Ɓ�*�t4s a��lyok��Flex/�:�Rw!mo?�P�A?�-�����`n�p�a SNBPJ AUTO-�06f����TB��PIABL�E1q 636��P�LN: RG$�pl�;pNWFMDB�V�I���tWIT 9tx�0@o��Qui#0|�ҺPN RRS?p�USB�� t &� remov�@ �)�_��&AxEPFT�_=� 7<`�pP:��OS-144 ���h s�g��@O�ST� � CRASH DU 9���$P�pW� .}$��LOGIN���8&�J��6b046� issue 6� Jg��: Sl�ow �st��c (Hos`�c��z�`IL`IMPRWtSPOT:Wh:0\�T�STYW ./ЏVMGR�h�T0C�AT��hos��EP�q��� �O�S�:+pRTU' k�-�S� ����E:��ppv@�2�� t\hߐr��m ��all���0�  $�H� WA�͐��3 CNT0s T�� WroU�alarm���0s�d � �0SE1���r: R{�OMEBp����K� 55��RE�àSEst��g  �   �KAN�JI�no���I�NISITALI1Z-p�dn1weρ<�6�dr�� lx`��SCII L�f�ails w�� <��`�YSTEa���8o��Pv� IIH����1W�Gro>Pm 7ol\wpSh@�P���Ϡn cflx�L@АWRI �OF� Lq��p?�F�u�p��de-rel}a�d "APo �SY�ch�Abet�we:0IND t0$gbDO���r�y `�GigE�#�operabilf  PAbHi�H`���c�lead�\e�tf�Ps�r�OS� 030�&: fig��GLA )P ���i��7Np tps�wx�B��If�g�������5aE�a EXCE#dU�_�tP�CLOS��"ro�b�NTdpFaU�c�!���PNIO_ V750�Q1�8�Qa��DB ��P� M�+P�QED�D�ET��-� \rk~��ONLINEhSBUGIQ ߔĠi`�Z�IB�S apA�BC JARKY�Fq� ���0MILT�`� R�pNД �p�0GAR��D*pR8��P�"! jK�0c�T�P�Hl#n�a�Z�E V�� TASK�$VP2(�4`
��!�$�P�`WIBP�K05�!FȐB/���BUSY RUNN�� "�򁐈�2�R-p�LO�N�wDIVY�CUL���fsfoaBW �p���30	V���ˠIT`�a505�.�@OF�UNE�X�P1b�af�@�E���SVEMG� N�MLq� D0pCC_SAFEX 0c�0u8"qD �PET�`9N@�#J87����RsP�A'�M�K��`K�H GUN�CHG۔MECH��pMc� T�  y�, g@�$ ORY LEAKA�;��ޢSPEm�Ja��V�tGRIܱ�@�oCTLN�TRk��FpepR�j50�E�N-`IN�����p `�`�Ǒk!��T3/d\qo�STO�0A�#
�L�p �0�@�Q��АY�&�;pb1TO8pP�s���FB�@YpL`�`DU��aO�sHupk�t4 � P�F� �Bnf�Q�PSVG�N-1��V�SRS	R)J�UP�a2�Qx�#D�q l O��~�QBRKCTR5� ��|"-�r�<pc�j!�INVP�D ZO�� ��T`h#�Q�cHs�et,|D��"DU�AL� w�2*BRV�O117 A]�T�Nѫt�+bTa247`3��q.?��sAUz��i�B�comple�te��604.�� -�`hancZ�U� F��e8�'�  ��npJtPd!�q��`��� 5h596p�!5d�� "p �P�P�Q�0�P2�p�A�� xP��R(}\xPeJ� aʰI���E���1��p� j  �� xSt��^t �A�ApxP�q 5 sig��a��"AC;a��p
�bCexPb_p���.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o�dxPX�b]o2�� �cb�c��ixP�jupfrmp�dxP�o�`exe�ax�oFdxPtped}o���u`�cptlibxzxP�lcr�xrxP�\�blsazEdxP_fm�}gcxP�x���o�|sp�o�mc(��ob_jzop�u6�wQf��t��wms�1q���sld�)��jmc�o\�n��nuhЕ��|cst�e��>�pl�q�p�iwck���uv�f0uߒ��lvisyn�CgaculwQ�
E F  ! �Fc.fd�Qv�� �qw���Data Acquisi���nF�|1�RR631�`��TR�QDMCM� �2�P75H�1��P583xP1��7�1��59`�5�P5�7<PxP�Q����(0���Q��o pxP!/daq\�oA���@�� ge/�etd�ms�"DMER"؟,�pgdD���.��m���-��qaq.<᡾xPmo��h����f{�u�`13��MA�CROs, Sk�saff�@z����03��SR�Q(��Q6��1"�Q9ӡ�R�ZSh��P^xPJ643�@7ؠ�6�P�@�PRS�@����e �Q�UС PI�K�Q52 PTLqC�W��xP3 (��p/O��!�Pn ��xP5��03\s�fmnmc "M�NMCq�<��Q��\$AcX�FM���ci ,Ҥ�X����cdpq+�6
�sk�SK�xP�SH560,P���,�y�refp "GREFp�d�A�jxP6	�of�OFc�<g6y�to�TO_���<�ٺ���+je|�u��caxis2��xPE�\�e�q"IS�DTc��]�prax ��MN��u�b�isde܃h�\��w�xP! isba�sic��B� P�]��QAxes�R�6������.�(Ba�Q�ess��xP����2�D�@�z�atis���(�{����h��~��m��FMc��u�{�
ѩ�MNIS ��ݝ����x����xٺ��x� j75���Devic�� Interfac�R<ȔQJ754��� xP�Ne`��xP��ϐ2�б����d=n� "DNE���~
tpdnui5cUI��ݝ	bd�b�P�q_rsof�Ob
dv_ar�o��u�����stchkc��z	 8�(}onl��G!ffL+H�J(��"l"/�n�b���z�hamp��T�C2�!i�a"�59��S�q��0 (�+P�o��u�!2��xpc_2p�cchm��CHMqP_�|8бpevwsp��2쳌pcsF���#C SenxPa�cro�U·�-�R6�Pd�xPk�����p���gT�L��1d M �2`��8�1c4ԡ�3v qem��GEM,�\i(��Dgesnd��5���H{�}Ha�@s1y���c�Isu�xD��Fmd��I��7�4����u���AccuC�al�P�4� ��ɢ7TޠB0��6+6f�6��99\aFF q�SA(�U��2�
X�p�!�Bd��cb_�SaU=L��  �� ?��ܖto��otplus\tsrnغ(�qb�Wp��t���1���Tool (N. A.)�[K�7�Z�(P�m����bdfcls� k94��"K4p��qtpa=p� "PS9H�>stpswo��p�L7��t\�q���� D�yt5�4�q��w�qк�� �M�uk��rkey����s��}tҾsfeatu6�E!A��� cf)t\Xq��0���d�h5����LRC0�md�!�587���aR�(����d2V��8c?u3l\�pa3}H�&r-�Xu�b��t,�� �q "�q �Ot��~,���{�/��1c�}����y�p�r� �5���S�XAg�-�y����Wj874�-? iRVis���Queu�� Ƒ� -�6�1���(����u���tӑ����
��tpvtsn "VTSN�3C�+�� v\pRDV����*�/prdq\�Q�&�vstk=P����Ƥ�nm&_�դ�cl�rqν���get@�TX��Bd���aoQ8Ͽ�0qstr�D[�� ��t�p'Z����nqpv��@�enlIP�0��D!x�'�|���s1c ߸��tvo/�� 2�q���vb��� �q���!���h]���(� Contr{ol�PRAX�P�5��556�A@5m9�P56.@56@�5A�J69$@9�82 J552 IDVR7�hqA����16�H���La��� ��Xe�frl�parm.f�FRL�am��C9�@(F�����w6{����A��QJ643�� 50�0LSE�
_pVAR $�SGSYSC��R�S_UNITS ��P�2�4tA�TX.�$VNUM_OLD 5�1�xP{��50+�"�` Funct���5tA� }�(�`#@�`3�a0�cڂb��9���@H5נ� �P���(�A���� �۶}����ֻ}���bPRb�߶~ppr4�TPSPI�3�}�r�10�#;A� t��
`���1���96 �����%C�� Aف��=J�bIncr�	�� ��\���1o5q{ni4�MNINp	�xP�`���!��Ho�ur  r� 2�21 �?AAVM����0 ��TUP� ��J545� ��6162��VCAM  (��CLIO ��R6�N2��MSC "P ~�STYL�Cv�28~ 13\��NRE "FHR�M SCH^��DCSU%ORSsR {b�04 ��EIOC�1 �j 542 � o�s| � egis�t�����7�1~�MASK��934"7 ��O�CO ��"3�8Ļ�2���� 0 �HB��� 4�"39�N� Re�� �L�CHK
%OPLG�%��3"%MHCR&.%MC  ; 4? ���6 dPI�54��s� DSW%MDr� pQ�K!637�0Ƚ0p"�1�Р"4 ��6<27 CTNY K � 5 ���"I7��<25�%/�T�%OFRDM� �Sg!<��930 FB( �NBA�P� ( HL�B  Men�S�M$@jB( PVC ���20v��2HT�C�CTMI�L��\@PAC 116U�hAJ`SAI \@�ELN��<29s�?UECK �b�@�FRM �b�OR\���IPL��Rk0�CSXC ���V�VFnaTg@HTTsP �!26 ���G�@obIG{UI"%IPGS�r>� H863 qb�!8�07r�!34 �r�84 \so`! QLx`CC3 Fb�21��!96 rb!51� ���!53R% 1�!s3!��~�.p"9�js VATFUJ7�75"��pLR6^RP�WSMjUCTO��@xT58 F!80����1XY ta3!7�70 ��885&�UOL  GTSo
�<{` LCM �r| gTSS�EfP6 W�>\@CPE `��0cVR� l�QNL"���@001 imrb�c3 =�b�0����0�`6 w�b-P-� R-�b8n@5EW�b9 �Ґa� ����b�`ׁ�b2 20�00��`3��`4*5�`5!�c�#$�`�7.%�`8 h60�5? U0�@B6E�"aRp7� !Pr8� t�a@�tr2 'iB/�1vp3�vp�5 Ȃtr9Σ�a4r@-p�r3 F�Ⴐr5&�re`u��r7� ��r8�U�p9 �\h738�a�R/2D7"�1f���2&�7� �3 7)iC��4>w5Ip�NOr60 C�L�1bE6N�4 I�pyL�uP0��@N�-PJ8�N�8NeN�9 H�r`��E�b7]�|���88�Вࠂ9 2��a�`0�qЂ5�%U0O97 0��@1�0����1 (�q�3 5R���0���@mpU��0�0�7*��H@(q�\P"RB6�q124�b;��@����@06� x�3 pB/x�u ��x��6 H606�a1x� ��7 6 ����p�b155 �����7jUU162� �3 g��4�*�65 2e "_��P�4U1`���B�1���`0'�174� �q��P�E186g R ��P�7 ��P�8&�3 (�9o0 B/�s191�����@202��6� 3���A�RU2x� d��2 b2h`��4�᪂2�4����19v Q�2��u2Jd�Tpt2� ��H�a�2hP�$�5���!U2�p�p
�2�p��@!5�0-@��8 @��9��TX@�� �e5N�`rb26Af�2^R��a�2Kp��1y�b5(Hp�`
�5�0@�gqGA���a52ѐ�Ḳ-6�60ہ5� ׁ�2��8�E��9�EU)5@ٰ\�q5hQ`S*�2ޖ5�p\w�۲��pJ �-P��5�p1i\t�H�4��PCH�7j��phiw�@��P��x��559 ldu� P�D���Q�@������� �`.��P>�:��8�581�"�q�58�!AM۲T�Aw iC�a589��0@�x����5 �a��12׀0.�1���,��2����,�!P\h8���Lp ��,�7��6��0840\� ANRS 0C}A��p���{��ran��FRA��Д�е�� �A%���ѹ�Ҍ��� ��(����Ќ���� ����������ь�����$�G��1��ը���������� sxS�`q�  ������`64��M��iC/50T-H��`����*��)p46���� C��N����m7;5s֐� Sp���b46��v����Г/M-71?�7�З����42������C�2��-�а�70�r�E��/h����`O$��rD���c7c7C�q��Ѕ����L��/��2\imm7c7�g������`���(��e� ����"�������a0 r��c�T,�Ѿ�"��,�� ��x�Ex�m77t����k����5�����)�iC��-HS-�  B
_�>���+�Т�7U�]���Mh7
�s��7�������-9?�/260L�_������Q��������]�9pA/ @���q�S�х����h621��c��92����8��.�)92c0�g $�@�����)$��5$���pylH"O"
��21���t?�350����p��$�0�
�� �350!����0��9�U/0\{m9��M9A3�P��4%� s��3M$���X%u���"him�98J3����� i d �"m4~�103p�� <����h794̂�&R���H�0����\� ��g�5AU��՜��0�� �*2��00��#0�6�АՃ�է!07{r ���������kЙ@����EP �#������?��#!��;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/��?�ҽCD25L����u0�"l�2BL
#��B��\20�2_�r �re���X��1��N����A@��z��`C��pU��`��04H��DyA�\�`fQ���sU���\�5  ��� p�g�^t��<$85��p�+P=�ab1l��G1LT��lA8�!puDnE(�20T��qJ�1 e�bH85��h�b�Ռ�5[�16B@s��������d2�8�x��m6t!`Q ����bˀ���b#�(�6iB;S�p�!��3 � ��b�s��-`Є_�W8�_����6�I	$�X5�1�U85��R�p6S����/ �/+q�!�q��`�6o���5m[o)�m6s�W��Q�?��setC06p ��3%H�5��10p$����g/��JrH��  9��A�856���d�F�� ���p/2��@h�܅�✐)�5���̑v��(��m6���Y�H�ѝ̑m�6(�Ҝ��a6�DM����#-S�+��H2��� ��Ҽ�� �r̑���✐��l���p1����F���2�\t6h T6H����� ��'Vl���ᜐ�V@7ᜐ/����;3A7��p~S��������4�`圐�V���!3��2�PM[��%�ܖO�chn��ve�l5����Vq���_a�rp#��̑�.���2l_hemq$�.�'�6415���5����?����F�����5 g�L�ј[���1���𙋹1����M7NU�М��eʾ����Euq$D;��-�4��3&H�f�c�Ĝ�h�� ����u���〜���ZS�!ܑ4���M	-����S�$̑�ք �� 0��<�����.07shJ�H�v�� ��sF��S*󜐳����̑���vl�3�A�T��#��QȚ�Te��q�p�r����T@75j�5 �dd�̑1�(UL�&�(� ,���0�\�?���̑�a��� xSt ���a�e�w�2��(�2	�2�C��A/����\�+p�����21 9(ܱ�CL S���� B̺��7F���?�<�lơ1L����c�� ���u9�0����e!/q��O���9�K��r9 (��,�Rs���ז�5�G�m20Ac��i��w�2��:�0`�$��2�2l�0�@k�X�S� ,�ι2��hO���1!41w����2T@� _std ��G�y� �ң�H� jdgm����w0\�  �1L���	�P�~� W*�b��t 5�������3�,���E {������L��5\L��3�L�|# ~���~!���4�#�� O����h�L6A�������2璥����44�����[6\j4s��·���#��ol�E"w�8Pk��� ��?0xj�H1�1Rr��>��]�2a�2AHw�P ��2��|41�8 ��ˡ��{� �%�A<��� +�?�l��0�&�"��|�`Am1�2������3�HqB�� K�R��ˑb�W���Fs ���)�ѐ�!���ah�1����5��16�16C��C����0\imBQ��d���(�b��\B5�-���DiL���O�_�<��PEtL�E�RH�ZǠP8gω�am1l��u� ��̑�b�<����<�$�T�̑�F����I ̑�Dpb��X"�ᒢް�p� ���^�t��9�0\� j9�71\kckrcfJ�F�s�����c��e "CTME�r������!�a�`mai�n.[��g�`run}�_vc�#0�w��1Oܕ_u����bctme��Ӧ�`ܑ��j735�- K�AREL Use% {�U���J��(1���p� Ȗ�9��B@��L�9��7j�[�atk208 C"K��Kя��\��9��a��̹����c�KRC�a�o ��kc�qJ�&s�����Gr ſ�fsD��:y��s���A1X\j|хrdtdB�, ��`.v�q��� �sǑIf�Wfj�52�TKQuto� Set��J� �H5K536(�9i32���91�58(�i9�BA�1(�74O�,A$�(TCP A@k���/�)Y� ��\tpqtool�.v��v���! �conre;a#�C�ontrol R�e�ble��CNRE(�T�<�4�2���pD�)���S�552��q(g�� (򭂯4X��cOux�\sfu;ts�UTS`�i�栜���t�棂���? 6�T�!�SA OO+D6������ ���,!��6c+� igt�t6i��I0�TW8 ���la��vo58�o�bFå����i�Xh��!Xk�|0Y!8\m6e�!G6EC���v��6��@�������<16�A���A�6s����U�`g�T|ώ���r1�qR��˔Z4�T��� ��,#�eZp)g����<ONO0���uJ��t�CR;��F�a� xS�t�f��prdsuGchk �1��2&&$?���t��*D%$�r (�✑�娟:r��'��s�qO��<scr�c�C�\At�trld J"o�\�V�����Paylo�nf�irm�l�!�87���7��A�3ad �! �?ވI�?plQ��3��3"�q��x pl�`���d7��l�calC�uDu�8��;��mov������initX�:s8�O��a�r4 ��r6�7A4|�e Generatiڲ���q7g2q$��g R�� (Sh��c ,D|�bE��$Ԓ\P�:�"��4��4�4,�. sg��5�F�$d6"e�!p "�SHAP�TQ n7gcr pGC�a(��&"� ��"GDAL¶��r6�"aW<�/�$dataX:s�"tpad��[q�%tput;a__O7;a��o8�1�yl+s�r �?�:�#�?�5x�?�:	c O�:y O�:�IO�s`O%g�qǒ�?��@0\��"o�j92�;!�Ppl.Col�lis�QSkip #��@5��@J��D��@@\ވ�C@X�7���7�|s2��ptcls�LS�DU�yk?�\_ ets�`�< \�Q��@��d�`dcKqQ�FC;�b�J,�n��` (�D�4eN����T�{ ���'j(�c�q���/�IӸaȁ��̠H������зa�e\�mcclmt "�CLM�/��� ma�te\��lmpA�LM�?>p7qmc?����2vm�q��%�3s��_sv90�_x�_msu�2L^v_0� K�o�{in�8(|3r<�c_log8r��rtrcW�E �v_3�~yc롘�d�<�te��d�er$cCe� F	iρ�R��Q�?|�l�enter߄�|��(Sd��1�T�X�+fK�r�a99�sQ9+�5�r\t�q\� "FNDR����STD~n$LANG�Pgui��D⠓�S������sp�!ğ֙uf�ҝ�s����$�����e+�=����������������w�H�r\fn_�ϣ��$`x��tcpma��- �TCP�����R638 R�Ҡ��+38��M7p,���� ��$Ӡ�8p0Р�VS,�6>�tk��99�a�� B3���PզԠ��D�2�����UI��t���hq B���8��������p����re�ȿ��exe@4φ�B���e38�ԡG�rmpWXφ�var@�φ�3N�����vx�!ҡ��qҿRBT $c�OPTN as�k E0��1�R �MAS0�H593>/�96 H50�i�+480�5�H0��Dm�Q�K��7�0�g��Pl�h0ԧ�2�OR�DP��@"��t\mas��0�a��"�ԧ�����k�գR����ӹ`m��b��7Г.f��u�d��r>��splayD�E����1w�UPDT |Ub��887 (��Di{���v�Ӛ�� �⧔��#�B��㟳��o  ����a������60q��B���>��qscan��B���ad@�������q`�䗣�#���8��`2�� vlv�䀃Ù�$�>�b���!y S��Easy/���Util��룙�511 J�����9R7 ��Nor֠��inc),<6Q�� �`c��"4�[���G986FVRx S1o����q�nd6��� �P��4�a\ (��
  �������d��K�b9dZ���men7���o- Me`tyF���Fb�0�TUa�'577?i3R��\�5�u?��!� n���f������l\mh�Ц�űE|hmn�	��<!\O���e�1�� l!��y��Ù�\|p����B�����mh�@��:. aG!���/�t�55�`6�!X�l�.us��|Y/k)ensubL�
��eK�h�� �B \1;5g?y?�?�?D��?�*rm�p�?Ktbox O2K|?�G��C?A%ds���?1ӛ#� �TR��/��P� 4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?Ă�Q23t.�P׀al��Pr+OP517��#IN0a��Q(}g�N�PESTf3ua�P B�l�ig�h�6�aq���P � xS���`  n�0mb�umpP�Q969�g�69�Qq��P0�b�aAp�@Q� BOqX��,>vche�s�>vetu㒣=w/ffse�3����]�;u`aW��:zol�sm<ub�a-��]D�K�ibQ�c����Q<t�waǂ tp�Q҄T�aror Rec�ov�b�O�P�642����a�q��a�⁠QErǃ�Qry�з`�P'�T�`�aarൄ����	{'�pak7971��71��m0���>�pjot��P�Xc��C�1�adb -v�ail��nag��<�b�QR629�a�Q���b�P  �
�  �P��$�$CL[q �����������$�PS_DIGI�T��� "�!�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv��������*璬�1:PRODUC�T�Q0\PGST�K�bV,n�9�9�\���$�FEAT_IND�EX��~��� 搠ILECOMP ;���)��"��SETUP2 <����  N� !�_AP2B�CK 1=� � �)}6/E+%,/i/��W/�/~ +/�/O/�/s/�/?�/ >?�/b?t??�?'?�? �?]?�?�?O(O�?LO �?pO�?}O�O5O�OYO �O _�O$_�OH_Z_�O ~__�_�_C_�_g_�_ �_	o2o�_Vo�_zo�o o�o?o�o�ouo
�o .@�od�o�� �M�q���<� �`�r����%���̏ [�������!�J�ُ n�������3�ȟW�� ����"���F�X��|� ���/���֯e����� �0���T��x���� ��=�ҿ�s�ϗ�,Ϡ��9�b�� P/� 2) *.VRiϳ�!�*�����0�����PC�7�>!�FR6:"�c��χ��T��߽߀Lը��ܮx���G*.F��>� �	N��,�k��ߏ��STM �����Qа����!�iPend�ant Pane	l���H��F���4�p�����GIF��������u����JPG&P��<�����	PANELO1.DT���� �����2�Y@�G��
3w������//�
4 �a/�O///�/��
TPEINS.�XML�/���\��/�/�!Custo�m Toolba�r?�PASS�WORD/�F�RS:\R?? %�Passwor�d Config �?��?k?�?OH�6O �?ZOlO�?�OO�O�O UO�OyO_�O�OD_�O h_�Oa_�_-_�_Q_�_ �_�_o�_@oRo�_vo o�o)o;o�o_o�o�o �o*�oN�or� �7��m��&� ��\�����y��� E�ڏi������4�Ï X�j��������A�S� �w�����B�џf� ������+���O���� �����>�ͯ߯t�� ��'���ο]�򿁿� (Ϸ�L�ۿpς�Ϧ� 5���Y�k� ߏ�$߳� �Z���~�ߢߴ�C� ��g�����2���V� ���ߌ���?���� u�
���.�@���d��� ����)���M���q��� ��<��5r� %��[�& �J�n��3 �W���"/�F/ X/�|//�/�/A/�/ e/�/�/�/0?�/T?�/ M?�??�?=?�?�?s? O�?,O>O�?bO�?�O O'O�OKO�OoO�O_ �O:_�O^_p_�O�_#_ �_�_Y_�_}_o�_�_�Ho)f�$FILE�_DGBCK 1�=��5`��� ( ��)
SUMMAR�Y.DGRo�\M�D:�o�o
`D�iag Summ�ary�o�Z
CONSLOG�o�o�a�
J�aConsole logK��[�`MEMCH�ECK@'�o��^qMemory �Data��W��)�qHADO�W���P��sS�hadow Ch�angesS�-c-���)	FTP�=��9����w`qm�ment TBD�׏�W0<�)ETHERNET̏��^�q�Z��aEthernet bp�figurati�on[��P��DCSVRFˏ��Ïܟ�q�%�� verify allߟ�-c1PY���DI�FFԟ��̟a��p{%��diffc���q��1X�?�Q��� ����X��CHGD��¯ԯ�i��px��� ���2p`�G�Y�� ��� �GD��ʿܿq���p���Ϥ�FY3ph�O�a��� ��(�GD������y���p�ϡ�0�UP?DATES.�Ц�~�[FRS:\������aUpdates List����kPSRBWLD'.CM.��\��B���_pPS_ROBOWEL���_���� o��,o!�3���W��� {�
�t���@���d��� ��/��Se��� ��N�r�  =�a�r�& �J���/�9/ K/�o/��/"/�/�/ X/�/|/�/#?�/G?�/ k?}??�?0?�?�?f? �?�?O�?OUO�?yO O�O�O>O�ObO�O	_ �O-_�OQ_c_�O�__ �_:_�_�_p_o�_o ;o�__o�_�o�o$o�o Ho�o�o~o�o7�o 0m�o� ��V �z�!��E��i� {�
���.�ÏR����� �����.�S��w�� ����<�џ`������ +���O�ޟH�������8���߯n����$�FILE_��PR����������� �MDONLY 1=4�~� 
 ��� w�į��诨�ѿ���� ���+Ϻ�O�޿sυ� ϩ�8�����n�ߒ� '߶�4�]��ρ�ߥ� ��F���j�����5� ��Y�k��ߏ���B� ����x����1�C��� g������,���P��� ������?��Lu~�VISBCKR�|<�a�*.VD||�4 FR:\���4 Visi�on VD file� :Lbp Z�#��Y�} /$/�H/�l/�/ �/1/�/�/�/�/�/ ? �/1?V?�/z?	?�?�? ??�?c?�?�?�?.O�? ROdOO�OO�O;O�O �OqO_�O*_<_�O`_��O�__%_�_�MR_GRP 1>4��L�UC4  ;B�P	 ]�o�l`�*u����RHB ���2 ��� �?�� ���He�Y �Q`orkbIh�oJd�o�Sc�o�oL�D��L҄bJ��cF�5U�aSLみ�o�o E��PoE��E�i.#G9C�e>w�_}�Ay�AnW��lq?�J�AnK��xq0~�� F�@ �r�d�a}J���NJk�H9��Hu��F!���IP�s}?��`�.9�<9��896�C'6<,6�\b�}B���Bǥ�Casd�B�n;B���B��{-�(���A��;B����A���AƯ�A�v���,fp�PA�����|�ݏx����%���p�A6Β@U��{ �v�a�������П�� ��ߟ��<���i{~;BH�P �a`�<Q��QA[K����ï�T
6�P=��PJ�M˯�o�o�B��P5���@�3�3@���4�m�,�@�UUU��U�~w�>u.�?!x��^��ֿ���3��=�[z�=�̽=�V6<�=�=�=$q��~���@8�i7�G��8�D�8@9!�7���@Ϣ���cD�@ D�� CϫoV��C��P��P'� 6��_V� m�o��To�� xo�ߜo������A� ,�e�P�b����� ��������=�(�a� L���p���������^� ������*��N9r ]������� �8#\nY� }�������/ ԭ//A/�e/P/�/p/ �/�/�/�/�/?�/+? ?;?a?L?�?p?�?�? �?�?�?�?�?'OOKO 6OoO�OHߢOl��ߐ� ���O�� _��G_bOk_ V_�_z_�_�_�_�_�_ o�_1ooUo@oyodo vo�o�o�o�o�o�o Nu�� �������;� &�_�J���n������� ݏȏ��%�7�I�[� "/�描�����ٟ�� �����3��W�B�{� f�������կ����� ��A�,�e�P�b��� �����O�O�O��O �OL�_p�:_������ ���������'��7� ]�H߁�lߥߐ��ߴ� ������#��G�2�k� 2��Vw�������� ���1��U�@�R��� v������������� -Q�u��� r��6��) M4q\n��� ���/�#/I/4/ m/X/�/|/�/�/�/�/ �/?ֿ�B?�f?0� BϜ?f��?���/�?�? �?/OOSO>OwObO�O �O�O�O�O�O�O__ =_(_a_L_^_�_�_�_ ���_��o�_o9o$o ]oHo�olo�o�o�o�o �o�o�o#G2k V{�h���� ���C�.�g�y�`� ���������Џ�� �?�*�c�N���r��� �����̟��)�� M�_�&?H?���?���? �?�?����?@�I�4� m�X�j�����ǿ��� ֿ����E�0�i�T� ��xϱϜ�������� �_,��_S���w�b߇� �ߘ��߼������� =�(�:�s�^���� �������'�9� � ]�o����~������� ������5 YD V�z����� �1U@yd ��v�����/Я */��
/�u/��/�/ �/�/�/�/�/??;? &?_?J?�?n?�?�?�? �?�?O�?%OOIO4O "�|OBO�O>O�O�O�O �O�O!__E_0_i_T_ �_x_�_�_�_�_�_o �_/o��?oeowo�oP� �oo�o�o�o�o+ =$aL�p�� �����'��K� 6�o�Z������ɏ�� 폴� ��D�/ / z�D/��h/ş���ԟ ���1��U�@�R��� v�����ӯ������ -��Q�<�u�`���`O �O�O���޿��;� &�_�J�oϕπϹϤ� �������%��"�[� F��Fo�ߵ����ߠo ��d�!���W�>�{� b������������ ��A�,�>�w�b��� �������������=��$FNO ����\��
F0�l q  FLAG�>�(RRM_C�HKTYP  r] ��d �] ���OM� _MI�N� 	���� ��  XT SSB_CFG ?\ �����OTP�_DEF_OW � 	��,IR�COM� >�$G�ENOVRD_D�O��<�lTH�R� d�dq_�ENB] qR�AVC_GRP s1@�I X( / %/7//[/B// �/x/�/�/�/�/�/? �/3??C?i?P?�?t? �?�?�?�?�?OOO�AO(OeOLO^O�OoR�OU�F\� ��,�B,�8�?���O�O�O	_|_���  DE_��Hy_�\@@m_B��=�vR/��I�O�SMT�G�SUoo|&oRHOSTC�s1H�I� ���zMSM�l[�bo�	127�.0�`1�o  e�o�o�o#z�o�FXj|�l60s	�anonymou�s������Q�ao�&�&��o �x��o������ҏ� 3��,�>�a�O�� ��������Ο�U%�7� I��]����f�x��� �����ү����+� i�{�P�b�t������ ������S�(�:� L�^ϭ�oϔϦϸ��� ���=��$�6�H�Z� ����Ϳs�������� ��� �2���V�h�z� ��߰���������
� �k�}ߏߡߣ���� ����������C�* <Nq�_���� ��-�?�Q�c�eJ ��n����� ��/"/E�X/j/ |/�/�/�%'/ ?[0?B?T?f?x?� �?�?�?�?�??E/W/�,O>OPObO�KDaEN�T 1I�K P�!�?�O  �P �O�O�O�O�O#_�OG_ 
_S_._|_�_d_�_�_ �_�_o�_1o�_ogo *o�oNo�oro�o�o�o 	�o-�oQu8 n������� �#��L�q�4���X� ��|�ݏ���ď֏7����[���B�QUICC0��h�z�۟���1ܟ��ʟ+���2�,���{�!ROUTER|�X�j�˯!PCJOG̯���!192.�168.0.10���}GNAME �!�J!ROBO�T�vNS_CFG� 1H�I ��Auto-started�$/FTP�/���/ �?޿#?��&�8�J� �?nπϒϤ�ǿ��[� �����"�4ߵ&���� ������濜������� ���'�9�K�]�o�� �����������/ �/�/G���k��ߏ��� ����������1 T���Py���� �"�4�	H-|�Q cu�VD��� �/�;/M/_/q/ �/����/
/�/> ?%?7?I?[?*/?�? �?�?�/�?l?�?O!O 3OEO�/�/�/�/�?�O  ?�O�O�O__�?A_ S_e_w_�O4_._�_�_ �_�_oVOhOzO�O�_ so�O�o�o�o�o�o�_ '9Kno�o� ����o*o<oNo P5��oY�k�}����� pŏ׏����0����C�U�g�y���_�T_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
 �.�FFF9E3����FRS:D�EFAULT��FANUC W�eb Server�
������q��������������WR�_CONFIG ;O�� ����IDL_CPU_kPC"��B���= �BH#MIN�.�BGNR_I�O��� ���% NP�T_SIM_DO�s}TPMOD�NTOLs �_�PRTY�=!O�LNK 1P�� �'9K]o>�MASTEr ��|���O_CFG�ƟUO����CY�CLE���_A�SG 1Q���
 q2/D/V/h/z/ �/�/�/�/�/�/�/
?�?y"NUM�x��Q�IPCH���£RTRY_C�N"�u���SCRQN������ ���R����?���$J23_DS/P_EN����~�0OBPROC�3ܷ�JOGV�1S�_�@��8�?р';ZO'??0CPO�SREO�KANJI_�Ϡu�A#��3T ���E�O�ECL_LM B2e?�@�EYLOGGINʭ������LA�NGUAGE ,_�=� }Q���LG�2U�����J �x�����PC �� �'0������MC:\RS�CH\00\˝L�N_DISP �V�������TOYC�4Dz\A�S�OGBOOK W+��o���o�o���Xi�o�o�o�o�o�~}	x(y��	�ne�i�ekElG_BUFF 1X�	��}2����Ӣ ������'�T� K�]�����������ɏ ۏ���#�P��Ëq�DCS Zxm =���%|d1h`�ฟʟܟ�g�IO ;1[+ �?'����'�7�I�[�o�� ������ǯٯ���� !�3�G�W�i�{�����б�ÿ׿�El TM  ��d��#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g��yߋߝ߈t�SEVt�0m�TYP΁� ��$�}�AR�S"�(_�s�2FL 31\��0�������������5�T�P<P���DmNGNAM�4�U�f�7UPS`GI�5�A��5s�_LOAD�@G %j%@_MOV�u�����MAXUALRM B7�P8��y���3�0Q]&q��Ca]s�@3�~�� 8@=@^+� طv	���V0+�P�A5d�1r���U�� ����E(i Ty������ �/ /A/,/Q/w/b/ �/~/�/�/�/�/�/? ?)?O?:?s?V?�?�? �?�?�?�?�?O'OO KO.OoOZOlO�O�O�O �O�O�O�O#__G_2_ D_}_`_�_�_�_�_�_ �_�_o
ooUo8oyo do�o�o�o�o�o�o�o��o-��D_LDX�DISA^�� �M�EMO_APX�E� ?��
  �0y�����������ISC 1_�� �O�� ��W�i�����Ə�� ���}��ߏD�/�h� z�a����������� ���@���O�a�5� �����������u�� ׯ<�'�`�r�Y���� ��y�޿�ۿ���8� ��G�Y�-ϒ�}϶ϝ� ����m�����4��X��j�#�_MSTR �`��}�SCD 1as}�R���N��� �����8�#�5�n�Y� ��}���������� ��4��X�C�|�g��� ������������	 B-Rxc��� ����>) bM�q���� �/�(//L/7/p/ [/m/�/�/�/�/�/�/ ?�/"?H?3?l?W?�?�{?�?�?�?n�MKC_FG b���?~��LTARM_�2�cRuB ��3WpTNBpMETsPUOp�2�����NDSP_CMN�TnE@F�E�� 	d���N�2A�O�D��EPOSCF�G��NPSTOL 1�e-�4@�<#�
;Q�1;UK_YW7_Y_ [_m_�_�_�_�_�_�_ o�_oQo3oEo�oio�{o�o�a�ASING_CHK  �M^AqODAQ2CfO��7J�eDEV }	Rz	MC:'|�HSIZEn@�����eTASK %�<z%$123456789 ��u�gTRIG 1g�� l<u%���3`���>svvYPaq���kEM_INF� 1h9G �`)AT&�FV0E0(���)���E0V1&A�3&B1&D2&�S0&C1S0=>��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ߏP� �t�������]�ί�� ���(�۟�^�� #�5�����k�ܿ� � ��ů6��Z�A�~ϐ� C���g�y�������� 2�i�C�h�ό�G߰� �ߩ��ߙϫ������ ��d�v�)ߚ��߾�y� ��������<�N�� r�%�7�I�[������ 9�&��J[��g��>ONITO�R�@G ?;{  � 	EXEC�1�3�2�3�4��5��p�7�8
�9�3�n�R� R�RRR R(R4R@RL�R2Y2e2q2�}2�2�2�2��2�2�3Y3�e3��aR_GRP_SV 1it���q(�5�
�4w-8��"�۵MO~q_DCd~�1�PL_NAME �!<u� �!�Default �Personal�ity (fro�m FD) �4R�R2k! 1j)T?EX)TH��!�AX d�?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O�Ox2-?�O�O�O_�_0_B_T_f_x_�b< �O�_�_�_�_�_�_o@ o2oDoVoho&xRj"g 1o�)&0\�bO, �9��b�a� @D�  �a?���c�a?�`�a�aA�'�6�ew;��	l�b	 �xJp���`�`	p �<� �(p� ��.r� K�K ���K=*�J����J���JV���kq`q�P��x�|� @j�@wT;f�r�f�qx�acrs�I�� ��p���p�r�ph}��3��´  ��>��ph�`z��꜖"g�Jm�q� H��N��ac��$�dw�� � �  P� Q� �� |  �а�m�Əi}	'�� � �I�� �  �����:�È���=���(��#�a�	���I  �n @H�i~�ab��Ӌ�b�$w���"N<0��  'Ж�q��p@2��@�����r�q5�C�pC>0C�@ C��z��`
�A1�q   @�B�V~X�
nwBD0h�A��p�ӊ�p�`���aDz���֏࿯�Я	�pv�(� �� -���I��-�=��A�a��we_q�`�p �??�ff ��m�|�� �����Ƽ�!1!ݿ�>1�  P�apv(�`ţ�� �=�qst��?˙��`x`�� <
�6b<߈;����<�ê<�? <�&P�ς��AO��c1��ƍ�?offf?O�?&���qt@�.�J<?�`��wi4� ���dly�e߾g;ߪ� t��p�[ߔ�߸ߣ� ���� ����6�wh�F0%�r�!�����1ى����E��� E�O�G+� F�!���/���?�e�`P���t���lyBL�cB��Enw4������� +��R��s���������h�yÔ�>���I�mXj���A�y�weC��������#/*/c/�N/wi�����v/C�`� CHs/`
=$��p�<!�!��ܼ�'��3A�A�AR�1AO�^?��$�?������
=ç>�����3�W
=�s#�]�;e�׬a�@����{�����<�>�(�B�u���=B0�������	R��zH��F�G���G���H�U`E����C�+��}I�#�I��H�D�F��E��RC�j=�>�
I��@H��!H�( E?<YD0w/O *OONO9OrO]O�O�O �O�O�O�O�O_�O8_ #_\_G_�_�_}_�_�_ �_�_�_�_"oooXo Co|ogo�o�o�o�o�o �o�o	B-fQ �u������ �,��P�b�M���q� ����Ώ���ݏ�(� �L�7�p�[������ ʟ���ٟ���6�!��Z�E�W���#1( �3�9�K���ĥ ������Ư!3ǭ8���!4M�gs��,�IB+�8�J��a���{�d�d�����ȿ��(�ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ�������,���  %�� �� h�Vߌ�z߰�&�g�/ 9�$�������7�����A�S�e�w�  ������������~�2 F�$�&'Gb������,��!C���@����8�����F� D�zN�� F�P D�������)#B�'9K]o#�?���@@v
J4$8�8��8�.
 v�� �!3EWi{�����:� ���ۨ�1��$�MSKCFMAP�  ��� ���(.��ONREL  ��!9��EX_CFENBE'
#�7%^!FNCe/W$JOGOVLIME'�dO S"d�KEY�E'�%�RUN�,�%�SFSPDTY0g&P%9#�SIGNE/W$T1�MOT�/T!�_�CE_GRP 1-p��#\x��? p��?�?�?�?�?O �?OBO�?fOO[O�O SO�O�O�O�O�O_,_ �OP__I_�_=_�_�_ �_�_�_oo�_:o��TCOM_CF/G 1q	-�vo�o�o
Va_ARC�_b"�p)UAP�_CPL�ot$NO�CHECK ?	+ �x� %7I[m�� ������!�.+�NO_WAIT_�L 7%S2NT^a�r	+�s�_ER�R_12s	)9�� A,ȍޏ��x��x�&��dT_MO��}t��, Gq*o|q�9�PARAM��u	+��a�ß�'g{�� =?�345678901� �,��K�]�9�i��������ɯۯ��&g������C��cUM_?RSPACE/��|����$ODRD�SP�c#6p(OFF�SET_CART��o��DISƿ��PEN_FILE��!�ai��`OPTI�ON_IO�/��PWORK ve7s# ��V�ؤ��p�4�p�	 �М�p��<���RG�_DSBL  Đ�P#��ϸ�RI_ENTTOD ?��C�� !l�UT�_SIM_D$��"���V��LCT w}�h�iĜa[�>1�_PEXE�j�RATvШ&p%� ���2^3j)TEX)�TH�)�X d3�������%�7� I�[�m������� �������!�3�E���2��u����������� ����c�<d�A Sew���������Ǎ�^0OU�a0o(��(�����u2, ���O H @D7�  [?�aG1?��cc�D][<�Z�;�	ls���xJƵ��������< ��� ���2�H(��H�3k7HSM5G��22G���G�p
͜�'f�X/-,2�CR�>��D!�M#{Z/��37�����4y H �"�c/u/�/0B_�����jc��gt�!�/ �/��"t32����/6�  ��P%�Q*%��%�|T��S62��q?'e	'� �� �2I� ��  ��+==�C�ͳ?�;	�h	�0��I  �n @�2�.��Ov;�ٟ?&gN�]O C ''�uD@!� C�C�@F#H!�/�O�O� sb
���@��@��@�e`0B��QA�0Yv: �13Uwz$oV_�/�z_e_�_�_	��(� �� -��2�1�1ta�Ua�c����:A-���.  �?�ff���[o"oB�_U�`oXÜQ8��t�o�j>�1  Po�V(���eF0�f�Y�x��L�?�����xb�P<
6b<�߈;܍�<��ê<� <G�&�,/aA�;�r�@Ov0P?fff�?�0?&ip�T@��.{r�J<?�`�u#	�Bdqt�Y c�a�Mw�Bo� �7�"�[�F��j��� ����ُ����3�����,���(�E��� E��3G+� F��a��ҟ��� ��,��P�;���B�pAZ�>��B��6� <OίD���P��t�=����a�s�����6j�h���7o��>� S��O�����Fϑ�#A�a�_��C3Ϙ�x/�%?��?����P�����#	Ę��P �N||CH�����������@I��_�'�3A�A��AR1AO�^?�$�?���� �±
=ç>�����3�W
�=�#� U��e����B��@��{����<����(�B�u�����=B0�������	�b�H��F�G���G���H�U`E���C�+���I#�I���HD�F���E��RC�j=�[�
I��@�H�!H�( E<YD0� ���������� �9� $�]�H�Z���~����� ��������#5 Y D}h����� ��
C.gR �������	/ �-//*/c/N/�/r/ �/�/�/�/�/?�/)? ?M?8?q?\?�?�?�? �?�?�?�?O�?7O"O [OmOXO�O|O�O�O�O@�O�O�O�O3_Q(��g����b��gUU��W_i_2я3�8��_�_2�4�Mgs�_�_�RIB�+�_�_�a���{�miGo5okoPYo�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�uX���  �p�� �o��/��S��z
u@үܠ�������ڱ������������  /�M�w�e���������l2 F�$N��Gb��t��a�X`�p�S�C�y�@p��5�G�Y�۠F� �Dz�� F�P D��]��������ʯܯ� ��~~�?���@@��?�K�K���:K���
 �|� ������Ŀֿ���π�0�B�T�fϽ�V� ����{��1���$PARAM_M�ENU ?3���  �DEFPUL�SEr�	WAI�TTMOUT���RCV�� S�HELL_WRK�.$CUR_ST�YL��	�OP9T��PTB4�.��C�R_DECSN���e��ߑߣ��� ��������!�3�\��W�i�{���USE�_PROG %��%�����CCR����e����_HO�ST !��!��:���T�`�V���/�X����_TI�ME��^��  ~��GDEBUG\���˴�GINP_FOLMSK����Tfp\����PGA  �����)CH����TWYPE������ ������  -?hcu��� ����//@/;/ M/_/�/�/�/�/�/�/ �/�/??%?7?`?��WORD ?	=�	RSfu	�PNSUԜ2J9OK�DRTEy�]�TRACECTL� 1x3���� �`B C&�`�`�>�6DT �Qy3�%@�0D� �  %�T�2@&6D'6D(�6D)6D*6D`8B,�6D-6D.6D/6D0�6D16A�c2@2L��H�`8BV�8BR��8BM 8BJ�8BF�8B�6D6D	6D
6D�6D6D6D6D�6D^�8B6D6D�6D6D6D�8B*6D6D6D6DV�(8Bj�8B6D6DҀ�8B�8B!6D"6D# 6D�8B5OGOYOkO}O�O�O�O�O�O�O_ Y�H�mMo_oqo�o�o �o�o�o�o�o#5 GYk}��_-_ ?_�I]_o_�I�_�_�I �_�_�I�_�_�Io/o ����	��-�?� A_S_u�w_�_���_Ϗ.A:m~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n����� ���������"�4�F� X�j�|����������� ����0BTf x��r����� ,>Pbt� ������// (/:/L/^/p/�/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�& 8J\n���� �����"�4�F� X�j�|�������ď֏ �����0�B�T�f� x���������ҟ��� ��,�>�P�b�t��� ������ί���� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ����������� �*��$�PGTRACEL�EN  )�  ��(���>�_UP z/���m�u�Y��n�>�_CFG7 {m�W�(�En���PЬ� ���DEFSPD e|���aP��>��IN��TRL �}��(�8��IPE_CONFI��}~m��m����Ԛ�>�LID����=�GRP� 1��W���)�A ���&f�f(�A+33D��� D]� C�O� A@1��Ѭ(��d�Ԭ��0�0�� 	 1��1���G ´�����B� 9����O�9�s�(��>�T?�
5�������� =��=#�
���� P;t_��������  Dz (�
H�X ~i������ /�/D///h/S/�/���
V7.10�beta1��  A�E�"�ӻ�A (�� ?�!G��!>��r�"����!���!oBQ��!A\� P�!���!2p����Ț/8?J?\?n?};� ���/��/�?}/ �?�?OO:O%O7OpO [O�OO�O�O�O�O�O _�O6_!_Z_E_~_i_ �_�_�_�_�_�_'o 2o�_VoAoSo�owo�o �o�o�o�o�o.�R=v1�/�#F@ �y�}��{m��y =��1�'�O�a��? �?�?������ߏʏ� �'��K�6�H���l� ����ɟ���؟�#� �G�2�k�V���z��� �����o��ίC� .�g�R�d��������� �п	���-�?�*�c� ����Ϯ���� ��B�;�f�x����� ��DϹ��߶������ ��7�"�[�F�X��|� �����������!�3� �W�B�{�f������� �� �����/S >wbt���� ��=Ozό� �ψ����ϼ� / .�'/R�d�v߈߁/0 �/�/�/�/�/�/�/#? ?G?2?k?V?h?�?�? �?�?�?�?O�?1OCO .OgORO�OvO�O�O�� �O�O�O__?_*_c_ N_�_r_�_�_�_�_�_ o�_)oTfx�to ���/�o/ >/P/b/t/mo�| �������3� �W�B�{�f�x����� Տ�������A�S� >�w�b����O��џ�� ����+��O�:�s� ^�������ͯ���ܯ �@oRodo�o`��o�o �o��ƿ�o���*< N�Y��}�hϡό� �ϰ��������
�C� .�g�Rߋ�v߈��߬� ����	���-��Q�c� N�ﲟ���l����� ���;�&�_�J��� n�����������,� >�P�:L������� �����(�:�3 ��0iT�x�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?a?s? ��?�?X?�?�?�?�? O'OOKO6OoOZO�O ~O�O�O�O�O*\ &_8_r���_�_���$PLID_K�NOW_M  ~�� Q��TSV ��]�P��? o"o4o�OXoCoUo�o� R�SM_GRP� 1��Z'0{`J�@�`uf�e�`
�5� �gpk 'Pe]o�� ��������S+MR�c��mT�EyQ}? yR�������� ��폯���ӏ�G�!� �-������������ ����ϟ�C���)� ����������寧����QST�a1 1�j�)���P0� A 4��E2�D�V� h�������߿¿Կ� ��9��.�o�R�d�v�@���ϬϾ����2�90� Q�<3��A3�/�A�S��4l�~ߐߢ��5���������6
��.�@��A7Y�k�}���8���������MAD � )��P�ARNUM  �!�}o+��SCH
E� S�
��f���S��UPDf�x�|�_CMP_�`�H�� �'�UE�R_CHK-�a��ZE*<RSr��_�Q_MOG����_�X�_RES_G��!���D� >1bU�y�� ���/�	/����+/�k�H/g/ l/��Ї/�/�/�	� �/�/�/�X�?$?)? ���D?c?h?����?x�?�?�V 1��U��ax�@c]�@t�@(@c\�@��@D@c[�*@���THR_INR�r�J�b�Ud2FMA�SS?O ZSGMN�>OqCMON_QU?EUE ��U�V� P~P X�N$ U�hN�FV�@END8�A��IEXE�O�E���BE�@�O�COP�TIO�G��@PR�OGRAM %��J%�@�?���BT�ASK_IG�6^O?CFG ��Oz���_�PDATA�c�.�[@Ц2=�Do Vohozo�j2o�o�o�o �o�o);M j�INFO[��m� �D������ ��1�C�U�g�y��� ������ӏ���	�dwpt�l )�QE ?DIT ��_i�>�^WERFLX	C��RGADJ M�tZA�����?נ�ʕFA��IORIT�Y�GW���MPD�SPNQ����U�G�D��OTOE@1��X� (!A�F:@E� c�Ч!�tcpn���!�ud����!i�cm���?<�XY_��Q�X���Q)�� *�1�5��P��]�@�L���p��� �����ʿ��+�=Ϡ$�a�Hυϗ�*��P�ORT)QH��P��E��_CART�REPPX��SK�STA�H�
SSA�V�@�tZ	25?00H863���_�x�
�'��X�@�swPtS�ߕߧ���/URGE�@B��x	WF��DO�F"[�W\�������WRU�P_DELAY ��X���R_HO�TqX	B%�c���R_NORMALq^xR��v�SEMI�������9�QSKIP�'��tUr�x 	7�1�1��X�j�|� ?�tU������������ ��$J\n4 ������� �4FX|j� ������/0/ B//R/x/f/�/�/�/�tU�$RCVTM�$��D�� DCR�'���Ў!Cq��C�2AC���u?�A!>��R�<|�{:���p�� ������ʿ��Ҿ����|��:��o?�� <
6b�<߈;܍��>u.�?!<�&�?h?�?�? �@>��?O O2ODOVO hOzO�O�O�O�O�O�? �O�O__@_+_=_v_ Y_�_�_�?�_�_�_o o*o<oNo`oro�o�o �o�_�o�o�o�o�o 8J-n��_�� �����"�4�F� X�j�U������ď�� �ӏ���B�T�� x���������ҟ��� ��,�>�)�b�M��� ���������ïկ� Y�:�L�^�p������� ��ʿܿ� ����6� !�Z�E�~ϐ�{ϴϗ� ����-�� �2�D�V� h�zߌߞ߰������� ��
���.��R�=�v� ��k��������� �*�<�N�`�r����� �����������& J\?���� ����"4F�Xj|��!GN_�ATC 1�	;� AT&F�V0E0�A�TDP/6/9/�2/9�ATA��,AT%G1%B960�_+++�,��H/,�!IO_T?YPE  �%�#�t�REFPO�S1 1�V+ 'x�u/�n�/ j�/
=�/�/�/Q?<? u??�?4?�?X?�?�?^�+2 1�V+�/��?�?\O�?�O�?�!3 1�O*O<OvO�O��O_�OS4 1� �O�O�O_�_t_�_+_S5 1�B_T_f_�_o	oBo�_S6 1��_�_�_5o�o�o|�oUoS7 1�lo�~o�o�oH3l�oS8 1�%_����SMAS�K 1�V/  
8?�M��XNOS/�r�������!MOT�E  n��$��_CFG ����q����"PL_RANG������POWER� �����S�M_DRYPRG %o�%�P��TART ���^�UME_PRO�-�?����$_EXE�C_ENB  <���GSPD��Ր8ݘ��TDB��
�sRM�
�MT_'��T����OBO�T_NAME �o����OB_�ORD_NUM �?�b!H863  ��կ���PC�_TIMEOUT��� x�S232�Ă1�� L�TEACH PENDAN��w���-��Ma�intenanc?e Cons����s�"���KCLC/Cm��

���t��ҿ No U�se-��Ϝ�0�N�PO�򁋁z��.�CH_L��3����q	��s�?MAVAIL����糅��SPAC�E1 2��, j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��� ���ߚ� �2�D��� hߊ�|��`������ ����� �2�D�� h��|���`�������(��y���2���� 0�B���f�����{ ���3) ;M_����@��/� /44 FXj|*/���/��/�/?(??=?5 Q/c/u/�/�/G?�/�/ �?O�?$OEO,OZO6n?�?�?�?�?dO�? �?_,_�OA_b_I_w_7�O�O�O�O�O�_ �O_(oIoo^oofo�o8�_�_�_�_�_ �oo6oEf){�x��G �o�� ���
M� ���*�<�N�`� r�������w���o�収���d.��%� S�e�w����������� Ǐَ���Θ8�+�=� k�}�������ůׯ͟ ����%�'�X�K�]� ��������ӿ�������#�E�W� `� @�������x�����\�e����� ������R�d߂�8� j߬߾߈ߒߤ���� ������0�r���X� ������������8�����
�ύ�_M?ODE  �{��/S ��{|�2ς0�����3�	�S|)CWORKw_AD��x�*/R  �{�`� ��� _INTVA�L���d���R_O�PTION� ���H VAT_G�RP 2��up(N�k|��_�� ���/0/B/��h� u/T� }/�/�/�/�/ �/�/?!?�/E?W?i? {?�?�?5?�?�?�?�? �?O/OAOOeOwO�O �O�O�OUO�O�O__ �O=_O_a_s_5_�_�_ �_�_�_�_�_o'o9o �_Iooo�o�oUo�o�o �o�o�o�o5GY k-���u�� ���1�C��g�y� ��M�����ӏ叧�	� �-�?�Q�c������� ��������ǟ��;�M�_����$SC?AN_TIM��_%�}�R �(�#((�<04_d d 	
!D�ʣ���u�/������U��25���@�dD5�P�g��]	����������dd�x� � P���� ��  8� ҿ�<!���D��$�M� _�qσϕϧϹ���������ƿv���F�X��/� ;��ob��pm��t�_DiQ|̡  � l� |�̡ĥ�������!� 3�E�W�i�{���� ����������/�A� S�e�]�Ӈ������� ������);M _q������ �r���j�Tf x������� //,/>/P/b/t/�/��/�/�/�/�%�/  0��6��!?3?E?W? i?{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O*�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o 9oKo�O�OJ�o�o�o �o�o�o�o 2D Vhz�����`��
�7?  ;� >�P�b�t��������� Ǐُ����!�3�E��W�i�{�������ß �ş3�ܟ��&� 8�J�\�n�������������ɯ�����,� �+�	�12345678^�� 	� =5���f�x�������������
��.�@� R�d�vψϚ�៾��� ������*�<�N�`� r߄߳Ϩߺ������� ��&�8�J�\�n�� ������������� "�4�F�u�j�|����� ����������0 _�Tfx���� ���I>P bt������ �!/(/:/L/^/p/��/�/�/�/�/�/� 2�/?�#/9?K?]?��iCz  Bp�˚   ��h2���*�$SCR_�GRP 1�(��U8(�\x�d�@ >� �'��	  �3�1�2�4(1*�&�I�3�F1OOXO}m��D�@�0ʛ)����HUK�LM-�10iA 890�?�90;��F;�M61C D�:�CP�*�1
\&V�1	��6F��CW�9)A7Y	�(R�_�_�_�_�_�\���0i^�oO UO>oPo#G�/���o�'o�o�o�o�oB�B0�rtAA�0*  @�Bu&Xw?��ju�bH0{Uz�AF@ F�` �r��o����� +��O�:�s��mBqrr`����������B�͏ b����7�"�[�F�X� ��|�����ٟğ���N����AO�0�B�CU
�L���E�jqBq>m󙵔�$G@�@pϯ B���G�I
E��0EL_DEFA�ULT  �T�_�E���MIPOWERFL  
E*��7�oWFDO� *���1ERVENT �1���`(��� L!DUM_�EIP��>��j!AF_INE�<¿C�!FT�������!o:� ���a�!RPC�_MAINb�DȺ8Pϭ�t�VIS}�C�y�����!TP���PU�ϫ�d��E�!�
PMON_PR'OXYF߮�e4ߑ���_ߧ�f����!RDM_SRV��r��g��)�!R�dIﰴh�u�!
v��M�ߨ�id���!?RLSYNC��>��8���!ROS��4��4��Y�(� }���J�\��������� ����7��["4 F�j|�����!�Eio�ICE_KL ?%�� (%SVCPRG1n>���3D��3���4/D/�5./3/�6V/[/�7~/�/��D�/�9�/�+�@��/ ��#?��K?�� s?� /�?�H/�?� p/�?��/O��/;O ��/cO�?�O�9? �O�a?�O��?_� �?+_��?S_�O{_ �)O�_�QO�_�yO �_��Os���� >o�o}1�o�o�o�o�o �o�o;M8q \������� ��7�"�[�F��j� ������ُď���!� �E�0�W�{�f����� ß���ҟ���A� ,�e�P���t���������ί�y_DEV� ��M{C:��_!�OUT��2��?REC 1�`e��j� �� 	 �����ȿ����׿��!�
 �PJ�%6 (޷�&�!�a�}���,���0�  Z� �3��3��Ge3�c ���V��˒��� ��� $��H�6�l�~�`ߢ� ���ߴ������� �� �V�D�z�h����� ��������
��R� @�v���j��������� ����*N<^ �r����� �&J8Z�b �������"/ 4//X/F/|/j/�/�/ �/�/��2��/�/�/? :?(?^?L?�?�?v?�? �?�?�?�?�? O6OO FOlOZO�O~O�O�O�O �O�O_�O2_ _B_h_ V_�_n_�_�_�_�_�_ 
o�_.o@o"odoRoto vo�o�o�o�o�o�o <*`Np�x �������8� J�,�n�\��������� Ə�Ώ�����F�4��j�X���`�p�V 1-�}� P��1��ܺ�  7 y��TYPE\���HELL_CF�G �.�F��� � 	�����RSR������ӯ���� ���?�*�<�u�`�������������_�  ��!%Ϡ3�E��Q�\����M�o�p�����2���d]�K�:�HK ;1�H� u��� ����A�<�N�`߉� �ߖߨ������������&�8��=�OMM� �H���9�FT?OV_ENB&��!�1�OW_REG_�UI��8�IMWA�IT��a���OU�T������TIM������VAL|����_UNIT���K�1�MON_AL�IAS ?ew� ( he������ ������і��); M��q����d ��%�I[ m�<���� ��!/3/E/W//{/ �/�/�/�/n/�/�/? ?/?�/S?e?w?�?�? F?�?�?�?�?�?O+O =OOOaOO�O�O�O�O �OxO�O__'_9_�O ]_o_�_�_>_�_�_�_ �_�_�_#o5oGoYoko o�o�o�o�o�o�o�o 1C�ogy� �H����	�� -�?�Q�c�u� ����� ��ϏᏌ���)�;� �L�q�������R�˟ ݟ�����7�I�[� m��*�����ǯٯ� ���!�3�E��i�{� ������\�տ���� �ȿA�S�e�wω�4� �Ͽ����ώ����+� =�O���s߅ߗߩ߻� f�������'���K� ]�o���>������ ����#�5�G�Y���}���������n��$�SMON_DEF�PRO ������ �*SYSTEM*  d=���RECALL ?�}�� ( �}�/xcopy f�r:\*.* v�irt:\tmp�back7=>i�nspiron:?11828 Yb�t�� }0.a 6HZ_���4/s:orde�rfil.dat��Mbt�� }=+/mdb:�M Z��/�-�Q b/t/�/�/�</�a/ �/??);��/p? �?�?���]?�? O O%/�/�/[/lO~O�O �/�/FO�/�O�O_!? 3?�?W?h_z_�_�?�? L_�?�_�_
oO/O�O SOdovo�oo�O>o�O �o�o+_=_�_�o r���_D�__� ��'o�o�o]on��� ���o6�H��o�������
xyzrate 61 ��ˏݏ�n�������.�M�3304 H�Z�������3.@��a�s�������*�I���Y�������..�A��� ݯn�����%���G�Y� _����'�9�¯]� nπϒϥ���ɯ[��� ���#�5�ȿY�j�|� �ߡ���D�׿����� �1Ϻ�U�f�x��� ��J����������-� ��Q�b�t�������<� �ߚ���)��������p����N�6368ǟY��!� 3��as���� E�Y��/!�3� F��n/�/�/��6/ H/� ^/�/??&8 ��m??�?����Z?�?�?O!w�$S�NPX_ASG �1����9A�� P 0� '%R[?1]@1.1O y?�#s%dO�OsO�O �O�O�O�O�O __D_ '_9_z_]_�_�_�_�_ �_�_
o�_o@o#odo GoYo�o}o�o�o�o�o �o�o*4`C� gy������ �	�J�-�T���c��� ����ڏ�����4� �)�j�M�t�����ğ ������ݟ�0��T� 7�I���m�������� ǯٯ���$�P�3�t� W�i��������ÿ� ���:��D�p�Sϔ� wω��ϭ��� ���$� ��Z�=�dߐ�sߴ� �ߩ������� ��D� '�9�z�]������ ����
����@�#�d� G�Y���}��������� ����*4`C� gy����� �	J-T�c� �����/�4/ /)/j/M/t/�/�/�/ �/�/�/�/?0?4,D�PARAM ��9ECA �	U��:P�4�0$H�OFT_KB_CFG  p3?E�4�PIN_SIM  9K�6�?�?�?��0,@RVQSTP/_DSB�>�21O|n8J0SR ��;�� & MUL�TIROBOTTgASK=Op3�6�TOP_ON_ERR  �F�8�A�PTN �5��@A�BRI�NG_PRM�O �J0VDT_GR�P 1�Y9�@  	�7n8_(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2Dkhz� ������
�1� .�@�R�d�v������� ��Џ�����*�<� N�`�r���������̟ ޟ���&�8�J�\� ����������ȯگ� ���"�I�F�X�j�|� ������Ŀֿ��� �0�B�T�f�xϊϜ� ������������,� >�P�b�tߛߘߪ߼� ��������(�:�a� ^�p��������� �� �'�$�6�H�Z�l� ~��������������3�VPRG_COUNT�6��A�5'ENB�OM=�4�J_UPD 1�>�;8  
p2 ������ ) $6Hql~�� ���/�/ /I/ D/V/h/�/�/�/�/�/ �/�/�/!??.?@?i? d?v?�?�?�?�?�?�? �?OOAO<ONO`O�O �O�O�O�O�O�O�O_ _&_8_a_\_n_�_�_��_YSDEBU)G" � �Pdk	�PSP_PASS"�B?�[LOG [��m�P9�X�_  �g�Q?
MC:\d�_b_MPCm��o$�o�Qa�o �vf�SAV �m�:dUb�U\gSV��\TEM_TIM�E 1�� (�) �%��o	T1?SVGUNS} #�'k�spASK_OPTION" �gospBCC�FG ��| q�b�{�}`� ���a&��#�\�G��� k�����ȏ������ "��F�1�j�U���y� ��ğ���ӟ���0��T�f��UR���S� ��ƯA������ �� D��nd��t9�l����� ����ڿȿ����� "�X�F�|�jϠώ��� ����������B�0� f�T�v�xߊ��ߦؑ� ������(��L�:� \��p�������� ��� �6�$�F�H�Z� ��~������������� 2 VDzh� �������� 4Fdv��� ���//*/�N/ </r/`/�/�/�/�/�/ �/�/??8?&?\?J? l?�?�?�?�?�?�?�? �?OO"OXOFO|O2 �O�O�O�O�OfO_�O _B_0_f_x_�_X_�_ �_�_�_�_�_ooo Po>otobo�o�o�o�o �o�o�o:(^ Lnp�����O ��$�6�H��l�Z� |�����Ə؏ꏸ�� ��2� �V�D�f�h�z� ����ԟ����
� ,�R�@�v�d������� ��ίЯ���<�� T�f�������&�̿�� ܿ��&�8�J��n� \ϒπ϶Ϥ������� ���4�"�X�F�|�j� �߲ߠ���������� �.�0�B�x�f��R� �����������,�� <�b�P�������x��� ������&(: p^������ � 6$ZH~ l�������� /&/D/V/h/��/z/��/�/�/�/�&0�$�TBCSG_GR�P 2��%��  �1 
 ?�  /? A?+?e?O?�?s?�?�?��?�?�;23�<_d, �$A?1�	 HC���6>���@E�5CL � B�'2^OjH4J���B\)LFY�  A�jO�MB���?�IBl�O�O�@��JG_�@�  D	 �15_ __$YC-P{_HF_`_j\��_�]@0 �>�X�Uo�_�_6oSo@o0o~o�o�k�h�0�	V3.00~'2	m61c�c	*�`�d2�o�e�>�JC0(�a�i q,p�m-  �0�����omvu1J�CFG ��%e 1 #0vz��r�Brv�x� ���z� �%��I� 4�m�X���|������� �֏���3��W�B� g���x�����՟���� ����S�>�w�b� ����'2A ��ʯܯ�� ����E�0�i�T��� x���ÿտ翢���� /��?�e�1�/���/ �ϜϮ��������,� �P�>�`߆�tߪߘ� �߼��������L� :�p�^������� ����� �6�H�>/`� r�������������� �� 0Vhz8 ������
 .�R@vd�� �����//</ */L/r/`/�/�/�/�/ �/�/�/�/?8?&?\? J?�?n?�?�?�?�?�� �?OO�?FO4OVOXO jO�O�O�O�O�O�O_ _�OB_0_f_T_v_�_ �_�_z_�_�_�_oo >o,oboPoroto�o�o �o�o�o�o(8 ^L�p���� ���$��H�6�l� ~�(O����f�d��؏ ���2� �B�D�V��� ����n����ԟ
��� .�@�R�d����v��� �����Я���*�� N�<�^�`�r�����̿ ���޿��$�J�8� n�\ϒπ϶Ϥ����� ��ߊ�(�:�L���|� jߌ߲ߠ��������� �0�B�T��x�f�� ������������,� �P�>�t�b������� ��������:( JL^����� � �6$ZH ~l��^���d� � //D/2/h/V/x/ �/�/�/�/�/�/�/? 
?@?.?d?v?�?�?T? �?�?�?�?�?OO<O *O`ONO�OrO�O�O�O �O�O_�O&__6_8_ J_�_n_�_�_�_�_�_ �_�_"ooFo��po �o,oZo�o�o�o�o �o0Tfx�H �������,� >��b�P���t����� ����Ώ��(��L� :�p�^�������ʟ�� �ܟ� �"�$�6�l� Z���~�����دꯔo ��&�ЯV�D�z�h� ������Կ¿��
�� .��R�@�v�dϚτ��  ���� ��������$TBJ�OP_GRP 2�ǌ�� � ?������������_xJBЌ���9� �< ��X���� @����	 �C��} t�b  C��<��>��͘Ր���>̚йѳ33�=�CLj�f�ff?��?�ff�BG��ь�����t��ކ�>�(�\�)�ߖ�E噙�;���hCYj�� � @h��B�  �A����f��C�  Dhъ�1���O�4�N����
:���Bl^���j�i�l�l����A�ə�A�"��D9��֊=qH����нp�h�Q�;�A�j��o��@L��D	2��������$�6�>B��\��T���Q�ts>x�@33@���C���y�1�����>��Dh�����x�����<{�h�@i� ��t ��	���K& �j�n|��� p�/�/:/k/������!��	V�3.00J�m61cI�*� IԿ���/�' Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I�!CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;��;Q�T,8�4`� *�ϴ?�2����3\�X/O��ESTPARS  ���	���HR@ABL/E 1����0�É
H�7 8��9
GB
H
H����
G	
HE

H
HYE��
H�
H
H6FRD	IAO�XOjO|O�O�O�ETO"_4[>_P_�b_t_�^:BS _�  �JGoYoko}o�o�o�o �o�o�o�o1C Ugy����`#o RL�y�_�_�_�_�O�O��O�O�OX:B�rNUoM  ���P��� V@P:B_CFG ˭��Z�h�@��IMEBF_TT%AU��2@��VERS�q���R 1���
 �(�/����b�  ����J�\���j�|��� ǟ��ȟ֟����� 0�B�T���x�������R2�_���@�
��MI_CHAN��� � ��DBGL�V���������E�THERAD ?U��O������h�����ROUT6�!��!����~��SNMASKD�|�U�255.���#�����OOLO_FS_DI%@�u�.�ORQCTRL �����}ϛ3r� �Ϲ���������%� 7�I�[�:���h�z߯��APE_DETA�I"�G�PON_S�VOFF=���P_?MON �֍��2��STRTCH/K �^������VTCOMPAT���O�����FPRO�G %^�%M�ULTIROBO�TTݱ���9�PL�AY&H��_INSWT_Mް �������US�q��LC�K���QUICK�ME�=���SCR�EZ�G�tps� ���u�z���_��@@n�.�SR_GRP 1�^�_ �O�� ��
��+O=sa�쀚�
m��� ���L/C1 gU�y���� �	/�-//Q/?/a/��/	12345C67�0�/�/@Xt��1���
 �}�ipnl/� gen.htm�? ?�2?D?V?`Pa�nel setupZ<}P�?�?�?�?�?�? �??,O>O PObOtO�O�?�O!O�O �O�O__(_�O�O^_ p_�_�_�_�_/_]_S_  oo$o6oHoZo�_~o �_�o�o�o�o�o�oso �o2DVhz� 1'���
��.� �R��v����������ЏG���UALRM���G ?9�  �1�#�5�f�Y���}� ������џן���,���P��SEV  �����ECFG ��롽���A��   B���
 Q���^�� ��	��-�?�Q�c�u��������������� �����I��?���(%D�6� �$� ]�Hρ�lϥϐ��ϴ� ������#��G����c �߿U�I_Y�HIST 1���  (�� ���4/SOFT�PART/GEN�LINK?cur�rent=edi�tpage,��,�5ӷ��+�;��y ����menu��962,1;������M�_�,936 u�
��.�@���W�i� {���������R����� /A��ew� ���N�� +=O�s��������f��f/ /'/9/K/]/`�/�/ �/�/�/�/j/�/?#? 5?G?Y?�/�/�?�?�? �?�?�?x?OO1OCO UOgO�?�O�O�O�O�O �OtO�O_-_?_Q_c_ u__�_�_�_�_�_�_ ��)o;oMo_oqo�o �_�o�o�o�o�o�o %7I[m�  �������3� E�W�i�{������Ï Տ�������A�S� e�w�����*���џ� ����ooO�a�s� ��������ͯ߯�� �'���K�]�o����� ����F�ۿ����#� 5�ĿY�k�}Ϗϡϳ� B���������1�C� ��g�yߋߝ߯���P� ����	��-�?�*�<� u����������� ��)�;�M������ ����������l� %7I[���� ���hz!3 EWi����� ��v////A/S/�e/P���$UI_�PANEDATA 1�����!�  	�}w/�/�/�/�/?? )?>?��/i? {?�?�?�?�?*?�?�? OOOAO(OeOLO�O �O�O�O�O�O�O�O_.&Y� b�>RQ? V_h_z_�_�_�__�_ G?�_
oo.o@oRodo �_�ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_ ��!�3�E�W��{� �_����ÏՏ���`� �/��S�:�w���p� ����џ������+� �O�a��������� ͯ߯�D����9�K� ]�o��������ɿ�� �Կ�#�
�G�.�k� }�dϡψ����Ͼ��� n���1�C�U�g�yߋ� �ϯ���4�����	�� -�?��c�J���� ������������;� M�4�q�X������� ����%7��[ �������@ ��3WiP �t�����/ �//A/����w/�/�/ �/�/�/$/�/h?+? =?O?a?s?�?�/�?�? �?�?�?O�?'OOKO ]ODO�OhO�O�O�O�O N/`/_#_5_G_Y_k_ �O�_�_?�_�_�_�_ oo�_Co*ogoyo`o �o�o�o�o�o�o�o�-Q8u�O�O}��������)�>��U-�j�|��� ����ď+��Ϗ�� �B�)�f�M������� �������ݟ�&�S��K�$UI_PA�NELINK 1��U  ��  ���}1234567890s��������� ͯդ�Rq����!�3� E�W��{�������ÿ�տm�m�&����Qo�  �0�B�T�f� x��v�&ϲ������� ��ߤ�0�B�T�f�x� ��"ߘ���������� �߲�>�P�b�t��� 0������������ $�L�^�p�����,�>�������� $�0,&�[gI�m� ������> P3t�i��� �� -n��'/9/K/ ]/o/�/t�/�/�/�/ �/�/?�/)?;?M?_? q?�?�UQ�=�2"� �?�?�?OO%O7O�� OOaOsO�O�O�O�OJO �O�O__'_9_�O]_ o_�_�_�_�_F_�_�_ �_o#o5oGo�_ko}o �o�o�o�oTo�o�o 1C�ogy�� ���B�	��-� �Q�c�F�����|��� ����֏�)��M� ��=�?��?/ȟڟ ����"�?F�X�j� |�����/�į֯��� ��0��?�?�?x��� ������ҿY���� ,�>�P�b��ϘϪ� ������o���(�:� L�^��ςߔߦ߸��� ����}��$�6�H�Z� l��ߐ��������� y�� �2�D�V�h�z� ���-���������
 ��.RdG�� }����c��� <��`r���� ����//&/8/J/ �n/�/�/�/�/�/7� I�[�	�"?4?F?X?j? |?��?�?�?�?�?�? �?O0OBOTOfOxO�O O�O�O�O�O�O_�O ,_>_P_b_t_�__�_ �_�_�_�_oo�_:o Lo^opo�o�o#o�o�o �o�o ��6H� l~a����� ���2��V�h�K� ������1�U
� �.�@�R�d�W/���� ����П������*� <�N�`�r��/�/?�� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��+������:� L�/�p���e������� ���� ��6����ۏ��$UI_�QUICKMEN�  ����}��REST�ORE 1٩��  �A
�8m3 \n���G�� ��/�4/F/X/j/ |/'�/�/�//�/�/ ??0?�/T?f?x?�? �?�?Q?�?�?�?OO �/'O9OKO�?�O�O�O �O�OqO�O__(_:_ �O^_p_�_�_�_QO[_ �_�_I_�_$o6oHoZo loo�o�o�o�o�o{o �o 2D�_Qc u�o������ �.�@�R�d�v����ଏ��Џ⏜SCR�E� ?��u1sc� u2��3�4�5�6��7�8��US#ER����T���Sks'���4��5���6��7��8��� N�DO_CFG mڱ  �  � PDATE h���None��SEUFRAM/E  ϖ���RTOL_ABRqT����ENB(�~�GRP 1��	��Cz  A� ~�|�%|�������įB֦��X�� UH��X�7�MSK  hK�S�7�N�%u�T�%�����VIS�CAND_MAX�I�I�3���FA?IL_IMGI�z ��% #S���IMR_EGNUMI�
����SIZI�� ��ϔ,�ONTM�OU'�K�Ε��&����a��a���s�FR�:\�� � �MC:\(�\L�OGh�B@Ԕ �!{��Ϡ�����z MCV�����UD1 �EX�	�z ��PO6�4_�Q��nm6��PO!�LI��Oڞ�e�V�N�fy@`�I�� =	_�wSZVmޘ��`��WAImߠ�STAOT �k�% @��4�F�T�$#�x ��2DWP  ���P G��=���͎���_J�MPERR 1��
  �p2345678901�� ��	�:�-�?�]�c� ��������������<��$�MLOW�ޘ������_TI/�˘'���MPHASE'  k�ԓ� ���SHIFT%�1 Ǚ��<z�� _����F /|Se���� ���0///?/x/ O/a/�/�/�/�/�/�����k�	VSF�T1\�	V��MN+3 �5�Ք p�����A�  B8*[0[0�Πpg3a1bY2�_3Y�7ME���K�͗	6e���&%���M���b���	��$��TDINGEND3�4��4OH�+�G1�OS2OIV �I���]LREL�EvI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�Y?BOX �ǝf_V\��b�2�TI�190.0.��P83p\�V2�54p^�Ԓ	 ��S�_�[b��?robot84q_   p�<9o\�pc�PZo Mh�]Hm�_Jk@1�o�ZABCd��k�, ���P\�Xo}�o0 );M�q���������>��aZ�b��_V