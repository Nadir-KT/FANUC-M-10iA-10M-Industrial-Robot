��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  �(��ALRM_R�ECOV1  � $ALMOEkNB��]ONi��APCOUPL�ED1 $[P�P_PROCES_0  �1��  |UREQ�1 � $S�OFT; T_ID��TOTAL_E�Q� $� � NO��PS_SPI_oINDE��$��X�SCREEN�_NAME ��SIGN���� PK_FI�L	$THKY�MPANE� � 	$DUMMYR � u3|4|~�RG_STR1� � $TI}TP$I��1�{�����U5�6�7�8�9�0��z������1�1�1� '1
'2"GSB�N_CFG1 � 8 $CNV�_JNT_* |�$DATA_CM�NT�!$FLA�GS�*CHEC�K�!�AT_CE�LLSETUP � P $H�OME_IO,G��%�#MACRO��"REPR�(-DWRUN� D|3�SM5� UTOB�ACKU0 � $ENAB�ު!EVIC�TI� � D� DMX!2ST� ?0B�#�$INTERVA�L!2DISP_U�NIT!20_DO�n6ERR�9FR_�F!2IN,GRkES�!0Q_;3!4C_WA�471�8ҰW+0�$Y $sDB� 6COM�W!2MO� H.�	 \rVE�1�$F�RA{$O�UDcB]CTMP1k_FtE2}G1_�3T�B�2�GXD�#�
 d $C�ARD_EXIS�T4$FSSB�_TYP!AHK�BD_SNB�1AG�N Gn $SLOT_NUM��APREV4DE�BU� g1� ;1_E�DIT1 � U1G=� S�0�%$EP��$OP�U0L�ETE_OK�BU�S�P_CR�A�$;4AV� 0LACIw1�R�@k �1�$@MEN�@$D�V�Q`PvVA{�QL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�08� <za�q;�G0 � 
$WARNM�0f�!p�@� -s�pNST� �CORN�"a1FL{TR{uTRAT� �T}p  $ACCa1�p��|{�r�ORI�P�C�kRT�0_S~B� CHG�,I1 [ Th�`�"3I�pTYD(�@*2 3`#@� X�!�B*HDDcJ* TCd�2_�3_�4_�U5_�6_�7_�8_��94�ACO�$ <� �o�o�hK3 1#`�O_Mc@AC t� � E#6NGPvABA� �c1�Q 8��`,��@nr1�� d�P�0e��� cvnpUP&Pb26h���p�"J�p_R�r�PBC��J�rĘߜJV�@U� B��s}�g1��"Q@��P_*0OF�S&R @� RO1_K8T��aIT�3T�ONOM_�0�1p��3�P�D !�� Ќ@��hPV��mCEX�p� �0g0ۤ<�p�r
$TF�2Co$MD3i�TO�3��0U� F� R��Hw2tC1(�Ez�g0#E{"F�"F�F40CP@�a2 �@$�PPU�3N�)ύRևAXd�!DU��AI�3�BUF�F��@1c |pp���pPIT�� PP�M�M��y��F�SIMQSI�"ܢVAڤT�9��x T�`(z�M��P�B�qFAC5Tb�@EW�P1��BTur�MC�k �$*1JB`p�*1DEC��F���x����� �H0�CHNS_EMP�1�$G��8��@_�4�3�p|@P��3�TCc�(r/�0-sx���ܐ� MBi��!����J�R� i�SEGFRR��Iv �aR�Tp9N�C��PVF4r�>bx &��f {uJc!�Ja��� !28�pץ�AJ���SIZ�3S�c�B�TM���g��>JaRSINFȑb� ��q�۽�н�����L�3�B���CRC�e�3CCp���� c��mcҞb�1J�cѿ��.����D$ICb�C q�5r�ե��@v�'���SEV���zF��_�եF,pN��ܫ�p?�4�0A�! �r ���h�Ϩ��p�2��@�a�� �د�@�	�>�Cx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�IM��UR��QUA1w  $@TITO1�/S@S�!����"0�?DBPXWO��B0=!5�$SK���2M@DBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z�s��L�)$�/PAt���� %�/PAC�PEC�!&?��WPE�q�.'*?�#� RE|�p2(H ���O�0#$L|3$�$�#�B[�;���FO�_D��ROS�r�#������3RIoGGER�6PApS|����ETURN�2n�cMR_8�TUw���0EWM���M�GN�P���BLA�H�<E���P��&$P� �'P@�Q3�CkD{��DQ���4��11��FGO_AWAY�BMO�ѱQ#!�� CS_�)  �PIS� I g�b {s�C��A��[  �B$�S��AbP�@�E9W-�TNTVճ�BV�Q[C�(c`�UWr��P�J��P�$0��SAsFE���V_SV�b�EXCLU��NnONL2��SY��*a&�OT�a'�HI�_V�4��B���_G *P0� 9�_z���p ��ASG�� +nrr�@6A@cc*b��G�#@E�V.i|Hb?fANNUN$0,.$fdID�U�2�SC@�`�i�a��j�f�p�z��@I$2,O�c$FibW$}�OT9@��1 $DUM�MYT��da��dn��� � �E- ` ͑HE4(sg�*b�S|AB��SUFFIW�[�@CA=�c�5�g6�a�bMSW��E. 8̀KEYI5���TM�10s�qA�vIN���ї!��/ D��HOST_P!�rT��ta�`�tn��tsp�pEMӰ�V��� SBLc U}LI�0  8	8=ȳ�r�DTk0�!?1 � $S��ESAMPL��j�۰f璱f���I�0��[ $SUB�k�#0��C��T�r#a�SAV ʅ��c���C��P��fP$n0E�w YwN_B#2 0�`DI{dlpO(��9#�$�R_I��� �ENC2_S� 3  5�C߰�f�- �SpU���B�!4�"g�޲�1T���5X�j`ȷg���0�0K�4�AaŔA�VER�qĕ9g�D3SP�v��PC���r"��(���ƓVALMUߗHE�ԕM+�sIPճ��OPP ��TH��֤��P��S� �۰F��dpf�J� ��~(T�{ET+6 H�bLL_DUs�~a3@`{��3:���OTX"����s����0N_OAUTO�!7�pC$)�$�*��c4�*(�C�8�C, �"�p�&�L�� 8/H *8�LH < 6����c"�`, `Ĭ� kª�q��q��sq��T~q��7��8��9���0����1��1̺1�ٺ1�1�1 �1*�1�2(�2����U2̺2ٺ2�2�U2 �2�2�3(ʥ3��3��̺3ٺ3��3�3 �3�3��4(�ɢT�?��!9� <�9�&�z��I�1���M�TR��FE@'@� : ,<6��Q? �@P�?9��5�9�E@�@A��a�A� ;p�$TP�$V�ARI:�Z���UP�2�P< ���TD�e���K`Q�����BAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�H  ��P�Y�@`>�!>t ;E��sC�ST�D�@ D���c�<� 	C� �{��_���l���R�  ���FORCE�UP?b��FLUS
�`H�N>�F ���R/D_CM�@E������� ��@vMP��REMr F�Q��1k@��(�7Q
K4	NJ�5�EFFۓ:�@IN�2Q��OVO�OV=A�	TROV����DTՀ�DTMX � ��@�
ے_P�H"p��CL��_ TpE�@�pK	_(�Y�_T��v(��@A;QD� ������!00tܑ0RQ����_�a����M�7�C9L�dρRIV'�{�n�EARۑIOH#PC�@����B�B��cCM9@���R ��GCLF�e!DY�k(M�ap#5TuD�G��� �%|ʠFsSSD �s? P�a(�!�1���P_�!�(J�!1��E�3�!3�+=5�&�GRA��7��@��;�PW��OyNn��EBUG_S�D2H�P{�_E �A`�_�TERM`5Bi9'ORI#e0Ci5=���SM_�P��e0DVi5��s0A�9Ei5��qUP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1젎4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ3Q�E�p %B`�'EC����AR$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"�r�A��?���ERV��XQ�Y�� mG>@�BN��U\���R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`�!�GRSMT6�G�3�GR��13�aPA�L@���`�q�uH �� ���TOC�A�`P	P�`$O�P����p�ѡ�`�0O��RE�`R�4C�AO�p낎Be��`R�Eu�h�A��eo$PWR�IMu��RR_�cN��q=B �I&2H���p_A�DDR��H_LE�NG�B�q�q�qz�Rj��S�JڢSS��SKN��u\��u̳�u�ٳSE�A����HmS��MN�!K������b����OL�X��p����`ACRO3pJ�@��X�+�p�Q��6�OUP3��b_�IX��a�a1 ��}򚃳���(��H ��D��ٰ��氋�+IO2S�D���𯅣`�7�L $xd��`Y!_OFFr��PRM_��^�aTTP_+�H:�wM (|pOBJ]"l�p��$��LE~C�d���N � \��֑AB_�Tq�b��S�`H�LVh��KR"uHITC�OU��BG�LO�q���h�����`���`SS� ���HQW�#A:�Oڠ<`�INCPU2VISIOW�͑��n��t�o��to�ٲ�IO�LN��P 8��R���p$SLob� PUT_n�$$p��P& ¢ ��Y �F_AS�"Q���$L������Q  U�0	P4A��^���ZP�HY��-��x��U9OI �#R `�K�����$�u�0pP pk���$������p��UJ5�S-���N�E6WJOGKG̲DIS��Z�Kp���#T (�uAVF�+`��CTR�C
�FLA�G2Z�LG�dU ����؜�13LG_SIZ����b�4�a�,�a�FDl�I`�w�  m�_�{0a�^��cg� ��4�����Ǝ���{0<��� SCH_���aR7�N�d�VW���AE�"����4��UM��Aљ`LJ�@�DAUf�EAU�p��d|�r��GH�ba���BOO>��WL ?�6 �IT��y0�REC��SCR ܓ��D
�\���MARG m�!��զ ��d%�����S����W���U�� �JGM[�MNC�HJ���FNKEY�\�K��PRG��UqF��7P��FWD��HL��STP��V`��=@��А�RS��HO`����C9T��b ��7�[�UL���6� (RD� ����Gt��@CPO��������MD��FOCU��RGE]X��TUI��I��4�@�L��� ��P����`��P��9NE��CANA��B�j�VAILI�CL� !�UDCS_HII4��s�O�(!��S���S�����_BUFF�!Xj�?PTH$m�@��v`��D���AtrY�?P��j�3��`WOS1Z2Z3Z��1�� � Z � ���[aEȤ��ȤIKDX�dPSRrO�X��zA�STL�R}��Y&�� Y$E�C���K�&&8��п![ LQ�� +00�	P���`#qdt
��U�dw<���_ \ ?�4Г�\��Ѩ#�\0C4�] ��C�LDPL��UTRQ�LI��dڰ�)�$F�LG&�� 1�#�D���'B�LD�%�$�%ORGڰ5�2�PVŀ�VY8�s�T�r�$}d^� ���$6��$�%SB�`T� �B0�4�6RCLMC�4]?o?��9��MI�p}d_� d=њRQ���DSTB�p� �;F�HHAX�R �JHdLEXCESHr1!BM!p�a`�@/B�TyB��`a�p=F_A7Ji��KbOttH� K�db \Q����v$MBC�LI�|�)SREQUIR�R�a.\o�AXDEB�UZ��ALt M��c@�b�{P����2�A#NDRѧ`�`d;�2��ȺSDC��N�IN@l�K�x`��X� N&���aZ�����RPS�T� ezrLO�C�RIrp�EX�<fA�p�9A�AOD�AQ��f XY�OND�rMF,Łf �s"��}%�e/� �9�FX3@IGG�� g ��t"��ܓhs#N�s$R�a%���iL��hL�v�@�D'ATA#?pE�%��tR��Y�Nh t_ $MD`qI}�A)nv� ytq�ytHP`��Pxu��(�zsANSAW)�yt@��yuD+��)\b���0o�i �@CUw�V�p 0XewRR2��j Du��{Q��7Bd$CALIIA@��G��2���RIN��"�<OL��INTE��Ck��r^�آXb]���_N�qlk���9�*����B�m��DIV��DH�@���qnI$V�,��S�$��$AZ�X�o�*�����oH �$B�ELT�u!ACC�EL�.�~�=�ICRC�� ���D�T��8�$PS�@�"L�@�r��#^�S�E�<� T�PATH3���DI���3x�p�A_W ��ڐ���2nC��4��_MG�$DDx��T���$FW��Rp9��I�4��DE�7�PPABN��R?OTSPEE�[g�� J��[�C@4�~�@$USE_+�2VPi��SYY��Z�1 qYN!@A��ǦOFF�qǡMO�U��NG���OL����INC�tMa6���HB��0HBENCS+�8q9Bp�4�FDm�IN�Ix�]��BƉ�VE��#�y�23�_UP񕋳LOWL���p� B���Du�9B#P`�x ���ByCv�r�MOSI���BMOU��@�7PE�RCH  ȳOV ��â
ǝ����D �ScF�@MP����� !Vݡ�@y�j�LUk��Gj�p�UP=ó����ĶTRK��AYLOA�Qe��A��x������N`�F�RTI�A$��MOUІ�HB@�BS0�p7D5����x��Z�DUM2ԓ�S_BCKLSH_Cx�k����ϣ����=���ޡ �	ACLAL"q��1м@N��CHK� �S�RTY��^�%E1rQq_�޴_UM�@r�C#��SCL0��r�LMT_J1_�L��9@H�qU�E�O�p�b�_�e�k�e�S�PC��u���N�P	C�N�Hz \P��C�0~"XT��C�N_:�N9��I�S	F!�?�V���U�/����x�T���CB!�SH�:��E�E1T�T�����y���T��PAL ��_P��_� �=������!����Jb6 L�@��OG��G�TORQU��ONֹ��E�R��H�E�&g_W2���_郅P���I�I�%I��Ff`xJ�1�,~1�VC3�0BD:B��1�@SBJ�RKF9�0DBOL_SM��2M�P�_DL2GRV�����fH_p��d���COS���LNH�� ������!*,�baZ���fMY��_(�TH��)TH�ET0��NK23����"��CB�&CB�CAA�B�"��!��!�&SB� 2�%'GTS�Ar�CIMa������,4#97#$DU���H\1� ��:Bk62�:AQ(rSf$NE�D�`I��B$+5��$̀�!A�%�5p�7���LPH�E�2���2SC%C�%�2-&FC0JM&̀V��8V�8߀LVJV�!KV/KV=KVKKV
YKVgIH�8FRM���#X!KH/KH=KH�KKHYKHgIO�<OR�8O�YNOJO!KUO/KO=KOKKOYKOM&F�2�!+i%0d��7SPBALANgCE_o![cLE0H_�%SPc� &�b�&�b&PFULC��h�b�g�b%p�1k�%�UTO_��Tg1T2�i/�2N�� "�{�t#�Ѱ`�0�*�.�T��OÀ<�v �INSEG"�ͱR�EV4vͰl�DIF��ŕ�1lzw��1m���OBpq�я?�M�I{���nLCHW3ARY�_�AB��!�?$MECH�!o X��q�AX��P��p��7Ђ�`n 
��d(�U�ROB��C�Rr�H���c(��MSK_f`�p WP �`_��R/�k�z�����1S�~�|�`z�{���z��qINUq��MTCOM_�C� �q  ����pO�$NOR�En����pЂr� 8p GRe�uS�D�0AB�$XYZ_DA�1a���DEBUUq�������s z`$��COD��� L���p��$BUFIN�DX|�  <�M{ORm�t $فUA��֐���r��<��rG��u � $SIMUL  �S�*�Y�̑a�OBJ�E�`̖ADJUS<�ݐAY_IS��D�3����_FI�=��Tu 7�~� 6�'��p} =�C�}p�@:b�D��FRIr��MT��RO@ \�E}z��y�OPWOY�q�v0Y�SYS�BU/@v�$SOP�ġd���ϪUΫ}pPgRUN����PA���D���rɡL�_OUbo顢q�$)�/IMAG��w��0�P_qIM��L�IN�v�K�RGOVR!Dt��X�(�P*�J�|��0L_�`]��0�RB1�0��ML��ED}��p ��%N�PMֲ��Hc�w��SL�`q�w x �$OVSL4vS;DI��DEX�� ��#���-�V} *�N4�\#�B�2�G�B�2_�M�x� �q�>E� x Hw��p^��ATUSW����C�0o�s���BTMT�ǌ�I�k�4��x�԰q�y Dw�E&���@E�r��7�8�жЗ�EXE�����������f q�z �@w���UP'��$�pQ�XN�����x����� �PG΅�{ h $SUB����0_���!�_MPWAIv�P7�&��LOR���F\p˕�$RCVFAI�L_C���BWD�΁�v�DEFSP>!p | Lw����Я�\���UNI+�����H�R�+�}K_L\pP��t�P��p�}H�> �*�j�(�ts`~�N�`KETB�J%�J�PE Ѓ~��=J0SIZE����hX�'���S�OR��?FORMAT�`�Ӱc ��WrEM�t���%�UX��G��P�LI��p�  �$ˀP_SWI��pq�J_PL��A�L_ �����AR��B��� C��D��$E��.�C�_�U�� � �� ���*�J3xK0����TIA4��u5��6��MOM��@������ˀB�ЃAD����������PU� NR�������m��� A$PI�6q��	� ����K4�)6��U��w`��SPEEDgPG������� �Ի�4T�� � 8@��SAMr`��p\�]��MOV_� _$�npt5��5���	1���2��������Ȣ'�S�Hp�IN �'�@�+�����4($4+T+GAMM�Wf�1'�$GETH`�p���Da���

pOLIBR>�II2�$HI=�_g�t��2�&E;��(A�.� �&LW�-6<�)56�&�]��v�p��V��?$PDCK���q"��_?�����q� &���7��4���9+�� �$IM_SR�pD�s�rF��r&�rLE���Om0H�]��0�-�pq���PJqUR_SC�RN�FA���S_SAVE_D��dE@�NOa�CAA�b�d@ �$q�Z�Iǡs	�I�  �J�K� ����H�L� �>�"hq����� �ɢ�� bW^UST�A�F��M4��� a��)q`��3�WW�I@�v�_�=���MUAo�� � $PY+�θ�$W�P�vNG �{��P:��RA��RH��RO�PL�����q� (��s'�X;�OI�&��Zxe ���m�� p��ˀ�3s�O�O�O��O�O�aa�_т� |��q�d@��.v��.v@��d@��[wFv��E��F�% ,r;B�w��|�tP���PMvA�QUa ��qQ8��1�QTH��HOLG�QHYSf��ES��qUE�ptZB��Oτ�  ـPܐ(�A����v�!�%t�O`�q��u�"�p��FA��IROG�����Q2���o�"���p��INFOҁ��׃V����R�H�OI� (�0SLEQ������Y�3���$�Á��P0Ow0�j��!E0NU���AUT�A�CO�PY�=�/�'��@Mg�N��=�}1������M ��RG��Á���3X_�P�$;ख�`��W��P��@��������EXT_CYC bHᝡRpÁ��r��_NAe1!А���ROv`	�?� � ��ЇPOR_�1�E2�S�RV �)_�I�DI��T_�k�}�'���PdЇ�����5��6��%7��8i�H�SdB��-�2�$��F�p���GPLeAdA
�TAR�Б@���P��2�裔d� ,�0F1L`�o@YN��K��M��Ck��PWR�+�9ᘐ��DELiA}�dY�pAD�a�p�QSKIPN4� �A�$�OB`�NT�} ��P_ $�M�ƷF@\bIpݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q����TQ������ ���`�#�RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�d"�REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"�������2�Қ�߼���P������3�қ'�@9�K�]�o���4���������������5�ҝ!�3�E�W�i�{��6�Ҟ������P�������7�ҟ@-?Qcu�8����������SMSKÁ�l��a��EkA��MOT-E6�����@��݂TQ�IO}5�I8STP��POW@��� �pJ����p�����E�"$DS?B_SIGN�1UQ��x�C\��S23�2���R�iDEVICEUS�XRSR�PARIT��4!O�PBIT�QI�O?WCONTR+�TQX��?SRCU� MpS�UXTASK�3Nx�p�0p$TATU�P��qRS�0������p_XPC)�$�FREEFROMqS	pna�GET�0.��UPD�A�2E#�P� :��� !>$USAN�na8&����ERI�0�&RpRYq5*"_j@�qPm1�!�6WRK9�KD���6��QFR�IEND�Q�RUFxg�҃�0TOOL�6�MY�t$LEN�GTH_VT\�FCIR�pC�@ˀE> �+IUFIN-RM�ΕRGI�1ÐAITI�$GXñ3IvFG2v7G1���p3��B�GPR�p�1F�Oa_n 0��!RE��0p�53҅U�TC��3A�A�F �G(��":���e1n!��J�8 �%���%]��%�� 74��X O0�L
��T�3H&��8���%�b453GE�W�0�WsR�TD����T��M�����Q�T]�$V �2����1�а91T�8�02�;2k3�;3�:ifa�9-i�aQ0��NS��ZR$V��2B�VwEV�	V�B;�����&�S�`��F�"��k�@�2a�PS�E���$r1C��_3$Aܠ6wPR��7vMU�cS�t '�/89�G� 0G�aV`��p�d`���50�@��-��
25S�� �"�aRW����B�&�MN�AX�!�A:@�LAh��rTHIC¤1I���X�d1TF�Ej��q�uIF_C	H�3�qI܇7�Q�pG1RxV���]��:��u�_JF~�PR|ԀƱ�RVAT��� ��`���0R�榀DOfE��COU�Ա��AXI���O�FFSE׆TRIGNS���c����h������H�Y��IG#MA0PA�pJ�E��ORG_UNEV��J� �S������d �$CА��J�GROU����TqOށ�!��DSP���JOGӐ�#��_Pӱ�"O�q����@�&7KEP�IR��ܔ2�@M}R��AP�Q^��Eh0��K�SYS��q"K�PG2�BRAK�B��߄�pY�0=�d����`AD_������BSOC���N���DUMMY14�p�0SV�PDE_�OP�#SFSPD�_OVR-���C���ˢΓOR٧3N�]0ڦF�ڦ��OV���SF��p���F�+�r!���CC��1q"L�CHDL��REC�OVʤc0��Wq@M������RO�#��Ȑ9_+��� @0�e@�VER�$OF�Se@CV/ �2WD��}��Z2���T�R�!���E_F�DO�MB_CM4���B��BL�bܒ#��adtVQR�$0pd���G$�7�AM5�`�� eŤ��_M;��"'����8$CA�'�E�8�8$HB�K(1���IO<�8����QPPA�������
��Ŋ����DVC_DBhC;��#"<Ѝ�r!S�1[ڤ�S�y3[֪�ATIOq 1q� ʡU�3���CABŐ�2�CvP���9P^�B���_� �S�UBCPU�ƐS �P �M�)0NS�c�M�"r�$HW_AC��U��S@��SA�A~�pl$UNITm�l_�AT���e�Ɛ�CYCLq�NEC�A���FLTR_2_FIO�7(��)&�B�LPқ/�.�_S[CT�CF_`�Fb�l���|�FS(!E�e�CHA�1��4�D°"3�RSD��$"}�����_Tb�PROX����� EMi_��ra�8!�a !�̹a��DIR0�RAOILACI�)RMr�CLO��C���Qq���#q�դ�PR=�S��AC/�c 	���FUNCq�0rRINP�Q�0��2�!3RAC �B ��[8���[WARn���#BL�Aq�A�����DAk�\���LD0���Q��q2eq�TI"r8��K�hPRIA�!r"AF��Pz!=�;���?,`�RK���MǀI�!�DF_@B�%1�n�LM�FAq@H�RDY�4_�P@R�S�A�0� �MUL�SE@���a ���ưt��m�m$�1$�1$1�o����� x*�EG00����!cAR���Ӧ�09�2�,%� 7�AXE��RKOB��WpA��_l-���SY[�W!‎&S&�'WRU�/-1��@��STR������Eb� 	�%��J��A�B� ���&9�����O�To0 	$��A�RY�s#2��Ԓ�	�ёFI@��$LGINK|�qC1�aI_�#���%kqj2XYZ��t;rq�3�RC1j2^8'0B���'�4����+ �3FI���7�q����'���_Jˑ���O3�QO�P_�$;5���AT�BA�QBC��&�D�Uβ�&6��TURN߁"r�E11:�p��9GFL�`_���* �@�5�*7��Ʊ 1��� KŐM��&8����"r��ORQ ��a�(@#p=�j��g�#qXU�����mTOVEtQ:�M��i�� �U��U��VW�Z�A �Wb��T{�, ��@;� uQ���P\�i��UuQ�W`e�e�SERʑ
e	��E� O���UdAas��4S�/7����AX��B�'q ��E1�e��i��irp �jJ@�j�@�j�@�jP �j@ �j�!�f��i� �i��i��i��i� y�y�'y�7yTq�HyDEBU8�$ 32���qͲf2G �+ AB����رnSVS�7� 
#�d�� L�#�L��1W��1W�JA W��AW��AW�QW�@!�E@?D2�3LAB��29U4�Aӏ��C 7 o�ERf�5�� � $�@_ A6��!�PO��à��0#�
�_MRA�t�� d � T��ٔERR����;STY&���I��V�0��cz�TOQ�d�PL�[ �d�"��	��C�! � pp`T8)0���_V1Vr�a(Ӕ����2ٛ2�E�ĺ��@�H�E���$QW�����V!��$�P��o�cI��a�Σ	I�SHEL�L_CFG!�� 5��B_BA�Sq�SR3���� a#Sb���1��%��2��3��4���5��6��7��8���RO����I0�03NL�\CAB+�����ACK4�����,��\@2@�&�?�_PUf�CO. U�OUG�P~ ����m�������{TPհ_KAR�Ll�_�RE*��P���|�QUE���uP�����CSTOPI_AL7�l�k0��h�8�]�l0SEM�4Ĳ(�M4�6�TYN�SO���DIZ�~�AӸ����m_TM�MOANRQ��k0E�����$KEYSWITCH���m���{HE��BEAT��|�E- LE~����ȅU��F!Ĳ���B�O�_HOM=OGREFUPPR&��y!�� [�C��O��-E�COC��Ԯ0_IO�CMWD
�a�(qk��� � Dh1$���UX���M�β<gPgCFORC������OM.  � Q@�5(�U�#P, Q1��, 3��45� �SNPX_A�St�� 0��AD�D���$SIZ>��$VAR����TIP/�.��A�ҹM�ǐ��/�1�+ �U"S�U!Cz���F'RIF��J�S���5Ԓ�NF�Ѝ� �� xp`SI��TqE�C���CSGL��	TQ2�@&����� ���STMT��,�P� �&BWuP��SHsOW4���SV��$�� �Q�A00�@Ma}���� ������&���5��6���7��8��9��A ��O ���Ѕ�Ӂ���0��F��� G��0G ���0G���@G��PTG��1	1	1	U1+	18	1E	2��U2��2��2��2��U2��2��2��2��U2��2	2	2	U2+	28	2E	3��U3��3��3��3��U3��3��3��3��U3��3	3	3	U3+	38	3E	4�U4��4��4��4��U4��4��4��4��U4��4	4	4	U4+	48	4E	5�U5��5��5��5��U5��5��5��5��U5��5	5	5	U5+	58	5E	6�U6��6��6��6��U6��6��6��6��U6��6	6	6	U6+	68	6E	7�U7��7��7��7��U7��7��7��7��U7��7	7	7	�7+	78	7E��V�P��UPDs� � �`NЦ�5�Y�SLOt�� � �L��d���A�aT�A�0d��|�ALU�:ed�~�CUѰjgF�!aID_L�ÑeH�I�jI��$FILcE_���d��$2�vfSA>�� hO�~�`E_BLCK���b$��hD_CPU yM�yA��c�o�d��yY����R �Đg
PW��!� oqLA��S=�ts�q~tRUN�qst�q~t����qst�q~t ��T��ACCs���X -$�qLE�N;��tH��ph�_�I���ǀLOW_AXMI�F1�q�d2*�AMZ���ă��W�Im�8ւ�aR�TOR��p�g�D�Y���LAC�Ek�ւ�pV�ւ~�_�MA2�v�������T#CV��؁��T��ي �����t��������IJj�R�MA���J���m�u�b����q2�j�#�f�{�t�K�JK���VK;���H���3f��J0����JJ��;JJ��AAL��ڐ(��ڐԖ4Օ5����N1���ʋƀW�LP�_(�g�,��pr��� `�`GRO�Uw`��B��NF�LIC��f�REQ�UIRE3�EBU`��qB���w�2�����p���q5�p�� �\��APPR��C�}�Y�
ްEN٨CsLO7��S_M���H���u�
�qu�� ���MC�����N9�_MG��C�Co���`M�в�N�BRK�L�NOL|�N�[�R��_LINђ�|�=�	J����Pܔ������@�����������6ɵ��̲8k�D���ď� ��
��qx)��7�PATH3ǀL�B�L��H�wࡠ�6J�CN�CA�Ғ�lڢB�IN�rUCV��4a��C!�UM��Y,���aE�p�����ʴ���PAYLO�A��J2L`R_AN�q�Lpp����$�M�R_F2LgSHR��N�LO���Rׯ�`ׯ�ACRL_G�ŒЛ� ��9Hj`߂$HM��үFLEXܣ�qJ>�u� :�� �����������1�F1�V�j�@�R� d�v�������E���� ȏڏ����"�4�q� ��6�M���~��U�g�Hy�ယT��o�X�� w����藕?��� ��ǟِݕ�ԕ�����%�7��P��J�� � V�h�z���`cAT�採@�EL��S S��J|�Ŝ�;JEy�CTR��~��TN��FQ��HA_ND_VB-����v`�� $��F20M����ebSW�q��'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aDM)F�AW�Z`i�Aw�AA��X X�'pi�Dw��D��Pf�G�p�)S�Tk��!x��!N��DY�pנM�9$`%Ц� H��H�c�׎���0� ��Pѵڵ����������J��� ���1��R�6��QOASYMvř����v��J���cі�_SH>��ǺĤ�ED����������J�İ%�p�C�IDِ�_VI��!X�2PV_UN!IX�FThP�J��_R �5_Rc�cTz�pT�V�݀@���İ�߷��U $�������Hqpˢ3��aEN�3�SDI����O4d ��`J�� x g"IJAAȱz�aabp�coc��`a�pdq�a� �^�OMME��� h�b�RqT(`PT�@ � S��a7�;�Ƞ�@ȷh�a�iT�@<� �$DUMMY9�Q�$PS_��R�FC�E`$v �� ���Pa� XXƠ���STE����SBRY�M21_�Vu�8$SV_E�RF�O��LsdsCLRJtA��Odb`�O�p � D ?$GLOBj�_LO���u�q�cAp�rܛ@aSYS�qADqR``�`TCH  � ,��ɩb�oW_NA����7�Ac�TSR���l ���
* ?�&Q�0"?�;'?�I) ?�Y)��X���h���x� �����)��Ռ�Ӷ�;� �Ív�?��O�O�O�D>�XSCRE栘p5����ST��s#}y`���Ea/u_HA�q� TơgpTYP�b���PG�aG���Od0�IS_䓀d�UEMd� ����ppyS�qaRSM_�q�*eUNEXCEP)fW�`S_}pM�x����g�z�����ӑCO�U��S�Ԕ 1�!�UE&��Ubwr���PROGM�FL�@$CUgpPOX�Q��5�I_�`H�� � 8�� �_�HE�PS�#��`RY ?�qp�b�t�dp�OUS��� � @6p�v_$BUTTp�Rp>R�COLUMq�e���SERV5�P�ANEH�q� �; �@GEU����Fy��)$HELyPõ)BETERv�)ෆ���A � � ��0��0��0ҰSIN簪c�@N���IH�1��_� �֪�LN�rؓ �qpձ_ò=�s$H��TEXl�����FLA@��RELV��D`����j����M��?,�Š��m����"�U�SRVIEW�q�S <6p�`U�`��NFI@;�FOC�U��;�PRI@�m�`�QY�TRIP>�qm�UN<`Md�� #@p�*eWA�RN)e6�SRTO�L%��g��ᴰO�NCORN��RAU䘠��T���w�VI�N�Le� $�גPATH9�גCwACH��LOG�!�LIMKR����v����HOST��!�b�R��OB�OT�d�IM>� �� ���Zq��Zq;�VCPU_A�VAIL�!�EX
	�!AN���q��10r��1r��1 �ѡ�.�p�  #`C����@$TOOL��$��_JMP� ����e$SS����EaVSHIF��Nc�P�`ג��E�ȐR����OSU�R��Wk`RADILѮ��_�a��:�9a���`a�r��LULQ�$OUTPUT_3BM����IM�ABp �@�rTIL'SCO��C7� ������&��3 ��A���q���m�I�2G��V�pLe��}��yDJU��N_�WAIT֖�}Ҵ�{�%! NE�u��YBO�� ��� $`�t�S�B@TPE��NE�Cp�J^FY�nB_T��R�І�a$�H[YĭcB��dM� ��F� �p�$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"�`�"��[���P?� 4�ZABC~%��  $�"�R��
E`�$$C�LAS�������!E`4�� � VI�RT]��/ 0ABS�����1 5�� < �!F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZi{0�-�AXL�pl��!�n63  �{tIN��qztPRE�����v��p�uLARMRECOV 9l�rwtNG�� .;	 A   �|.�0PPLIC���?5�p��Handlin�gTool o� �
V7.50P�/23-�  �P�z��
��_S�Wt� UP�!�� x�F0��t�Qz�A� v� �864�� �it��y�2�2 7DA5��� �� d��@<ϐo�Noneisͅ�˰ ��T����!�Ayx>�_l�V�uT��s9�UTO�"�Њt��y��HGAPON�
0g�1��Uh�D [1581�����̟ޟry����Q 1���p�,� 蘦���;�@��q_���"�" �c�.�H���D�HTTHKYX� �"�-�?�Q���ɯۯ 5����#�A�G�Y�k� }�������ſ׿1��� ��=�C�U�g�yϋ� �ϯ�����-���	�� 9�?�Q�c�u߇ߙ߫� ����)�����5�;� M�_�q������� %�����1�7�I�[� m����������!�� ��-3EWi{ ������ )/ASew�� ��/��/%/+/ =/O/a/s/�/�/�/�/ ?�/�/?!?'?9?K? ]?o?�?�?�?�?O�?��?�?O#O]���TO��E�W�DO_CL�EAN��7��CNMw  � ��__/_A_S_�DS�PDRYR�O��H	Ic��M@�O�_�_�_ �_oo+o=oOoaoso��o�o���pB��v �u���aX�t������>9�PLUGG���G\��U�PRCvPB�@E��_�orOr�_7�SEGF}�K [mwxq�O�O���p��?rqLAP�_ �~q�[�m�������� Ǐُ����!�3�x�TOTAL�f yx�_USENU�p��� �H���B��RG_�STRING 1�u�
�M�n�S5�
ȑ_I�TEM1Җ  n 5�� ��$�6�H�Z� l�~�������Ưد����� �2�D�I�/O SIGNA�L̕Tryout Modeӕ�Inp��Sim�ulatedב�Out��OV�ERR�P = 1�00֒In c�ycl��בProg Abor���ב��Statu�sՓ	Heart�beatїMH� Faul��Aler'�W�E�W�iπ{ύϟϱ������� �CΛ�A����8� J�\�n߀ߒߤ߶��� �������"�4�F�X�8j�|���WOR{pΛ ��(ߎ����� ��$� 6�H�Z�l�~���������������� 2PƠ�X ��A{ ������� /ASew��p���SDEV[ �o�#/5/G/Y/k/ }/�/�/�/�/�/�/�/�??1?C?U?g?y?PALTݠ1��z? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�Op�O�O_�?GRI�` ΛDQ�?_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o2_l�R��a\_�o" 4FXj|��� ������0�B�<T��oPREG�>��  f���Ə؏����  �2�D�V�h�z��������ԟ���Z��$�ARG_��D ?�	���;���  	�$Z�	[O�]�O��Z�p�.�SBN�_CONFIG S;��������CII_SAVE  Z�����.��TCELLSET�UP ;�%HOME_IOZ�~Z�%MOV_��
�REP�lU�(�UTOBACKܠ���FRwA:\z� \�,z�Ǡ'`�z����n�INI�0z����n�MESSA�G���ǡC���OD�E_D������%�Ox�4�n�PAUSX�!�;� ((O>��ϞˈϾϬ��� �������*�`�N����rߨ߶�g�l TSK  w�Կ׿q��UPDT+��d�!�A�WSM_CF��;���'�-�GRP 2:�?�� N�BŰA��%�XoSCRD1�1
7�' �ĥĢ���� ������*������� r�����������7��� [�&8J\n���*�t�GROUN��UϩUP_NA��:�	t��_�ED�17�
 ��%-BCKEDT-�2�'K�`���-t�z�eq�q�z���A2t1�����q��k�(/��ED3 /��/�.a/�/;/M/ED4�/t/)?�/�.?p?�/�/ED5 `??�?<?.�?O�?�?ED6O�?qO�?�.MO�O'O9OED7 �O`O_�O.�O\_�O�OED8L_,�_�^�-�_ oo_�_ECD9�_�_]o�_	-09o�oo%oCR_  9]�oF�o�k� ~� NO_DEL���GE_UNUS�E��LAL_OUT ����WD_ABOR���~��pITR_R�TN��|NON�Sk���˥CA�M_PARAM �1;�!�
 8�
SONY XC�-56 2345�67890 �ਡ@���?�>�( А\�
�Ԫ�{����^�HR�5q�̹��ŏR57�ڏ�Aff���KOWA SC3W10M
�x�̆�d @<�
�� �e�^��П\�����*�<��`�r�g�CE_RIA_I��!�=�F���}�z� ��_LI�U�]�����<z��FB�GP 1��Ǯ�M�_�<q�0�C*  �����C1��9��@��G����CR�C]��d*��l��s��R��翪��[Դm��v���������� C�����(�����=�H=E�`ONFIǰ��B�G_PRI 1�{V���ߖϨ�������������CH�KPAUS�� 1K� ,!uD�V� @�z�dߞ߈ߚ��߾� �����.��R�<�b�4���O������^��_MOR��� �6��� 	  �����*��N�<���D����?��q?;��;����K��9�P��ça�A-:���	�

�� M���pU�ð��<��Y,~��DB�������)
mc:cpmidbg�f�3:��p��:¥��p�/�  Y�0�)�� X�s>��p��pa�U�?�� \Ug�/�+��p�Uf�M/�w�O/�
DEF �l��s)�< b?uf.txts/��t/��ާ�)�	`z�����=L���*[MC��1����X?43��1��t�~īCz  BHH��Co�C|���CqD���C���C�{i�Y
K�D��F.���F��E����F,E��ٟ�K�F�N�I�U��I?O�I�<#I6�I�Y	��H�$w�K1���s���U.�p������BDLw�M@x8��1Ҩ�����g@D�p@�0E�YK�EX�E�Q�EJP F��E�F� G���>^F E��� FB� H�,- Ge��H�3Y��:�  >�33 ���N~  n8�~@��#5Y�E>�ðA��Yo<#�
"Q ����+_�'RSMOF�S�p�.8��)T1>��DE ��C�
Q��;�(P  QB_<_��R����,	op6C4P�Y
s@E ]AQ�2s@C�0)B3�MaC{@@*cw���UT�pFPROG %�z�o�oig�I�q���v��ldKEY_TBL  �&�S�#� �	
��� !"#$�%&'()*+,�-./01i�:;�<=>?@ABC�� GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����vq���͓��������������������������������������������������?�������p`�LCK�l4�p`�`S�TAT ��S_AU_TO_DO����5�INDT_EN�B!���R�Q?�1�Ty2}�^�STOPb����TRLr`LET�E��Ċ_SCR�EEN �Z_kcsc��U���MMENU 1 ~�Y  <�l �oR�Y1�[���v�m� ��̟�����ٟ�8� �!�G���W�i����� ���ïկ��4��� j�A�S���w������ ��ѿ����T�+�=� cϜ�sυ��ϩϻ�� �����P�'�9߆�]� o߼ߓߥ�������� :��#�p�G�Y��� ���������$���� 3�l�C�U���y����� ������ ��	VY)��_MANUAL���t�DBCO[�R�IGڇ
�DBNUIM� ��B1 e
��PXWORK 1!�[�_U/4�FX�_AWAYz�i�GCP  b9=�Pj_AL� #��j�Y��܅ `�_�  1"�[ , 
�mg�&/~&JlMZ�IdPx@P�@#ONTIMهM� d�`&�
�e��MOTNEND��o�RECORD 1(�[g2�/{�O��!�/ky"? 4?F?X?�(`?�?�/�? ?�?�?�?�?�?)O�? MO�?qO�O�O�OBO�O :O�O^O_%_7_I_�O m_�O�_ _�_�_�_�_ Z_o~_3o�_Woio{o �o�_�o o�oDo�o /�oS�oL�o� ���@���+� yV,�c�u������ ��Ϗ>�P�����;� &���q���򏧟��P� ȟ�^������I�[� ���� ���$�6��������jTOLEoRENCwB���L�͖ CS_?CFG )�/'dMC:\U��L%04d.CS�V�� c��/#A V��CH��z� /�/.ɿ��(S�RC_�OUT *���1/V�SGN �+��"��#�1�9-FEB-20� 16:0001�7l�9:09+? PQ�8�ɞ��/.��f�pa�m��PJPѲ���VERSION� Y�V2�.0.84,EFLOGIC 1,�/ 	:ޠ=��ޠL��PROG_�ENB��"p�UL�Sk' ����_WRSTJNK ��"�fEMO_OPT?_SL ?	�#�
 	R575/#=�����0�B�|���TO  ��صϗ��V_F EX�d�%��PAT�H AY�A\p�����5+ICT�-Fu-�j�#�egS�,�STBF_TTS�(@�	d���l#!w�� �MAU��z�^"MS%WX�.�<�4,#�
Y�/�
!J�6�%ZI~m��$SBL_FAUL(�y0�9'TDIA[��1<�<� ����1234567G890
��P�� HZl~���� ���/ /2/D/V/hh/�� P� ѩ�yƽ/��6�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�,�/�UMP���� �ATR���1OC@�PMEl�OOY_T�EMP?�È�3pF���G�|DUNI���.�YN_BRK �2_�/�EMGDI_STA��]��E�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�a�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��aDzr�A W�_BWD�p��xf�́t�_DI�� 9�5�d�T�asRֆSTEP��:P��OP_DOv��f�PFACTOR_Y_TUNwdM��EATURE �:�5̀rQ�Handling�Tool �� \�sfmEng�lish Dictionary���roduAA� Vis�� Ma�ster����
�EN̐nalog� I/O����g.�fd̐uto S�oftware �Update  �F OR�mat�ic Backu�p��H596�,�ground �Editޒ  1� H5Cam�era�F��OP;LGX�ell𜩐�II) X�omm�Րshw���com揭co���\tp����pane�� � opl��tyl�e select^��al C��nJ�~Ցonitor��gRDE��tr��?Reliab𠧒�6U�Diagno�s(�푥�552�8�u��heck �Safety U�IF��Enhan�ced Rob �Serv%�q )� "S�r�UserG Fr[�����a���xt. DIO 6�fiG� sŢ��wendx�Err�MLF� pȐĳr�r�� ����  !���FCTN Men�u`�v-�ݡ���T�P Inېfac��  ER J�GC�pבk E�xct�g��H55�8��igh-Sp�ex�Ski1�  �2
P��?���m�munic'�on1s��&�l�ur�ې���ST Ǡ��c�onn��2��TX�PL��ncr�s�tru����"FA�TKAREL Cmd. LE�{uaG�545\�ſRun-Ti��E{nv��d
!����ؠ++�s)�S/�W��[�Lic�enseZ��� 4�T�0�ogBook�(Syڐm)��H�54O�MACRO�s,\�/Offs�e��Loa�MH�������r, k�M�echStop �Prot���� l�ic/�MiвSh�if����ɒMixpx��)���,e�S��Mode Swiwtch�� R5W��Mo�:�.�� 7#4 ���g��K��2h�ulti-T�=�M���LN (�Pos�Reg�iڑ������d�ݐtO Fun�ǩ�.�����Num~����Ï lne��ᝰ Adjup������  - W��ta�tuw᧒T��RDMz�ot��s�cove U�9����3Ѓ�uesOt 492�*�o������62;�SNP�X b ���8 Jy7`���Libr��FJ�48���ӗ� ����
�6O�� Pa�rts in VCCMt�32���x	�{Ѥ�J990��{/I� 2 P���TMILIB��Ht���P�AccD��L�
TE$TX܍ۨ�ap1S�Te<����pkey���wգ�d��Un�exceptx�motnZ��������3є�� O��΄� 90J�єSP CSXC<�f�l�Ҟ� Py�We}�Β�PRI�>vr\�t�men�� ��/iPɰa������vGrid�play��v��0�)��H1�M-10iA(B201 ��2\� 0\k/�A/scii�l�Т��ɐ/�Col��ԑG7uar� 
�� /�P-�ޠ"K��stN{Pat ��!S��Cyc�҂�or�ie��IF8�ata- quҐ�� ƶ���mH574��RML��am���Pb�HMI De3�(�b����PCϺ�P�asswo+!��"PE? Sp$�[���stp��� ven���Tw�N�p�YEL?LOW BOE	k$wArc��vis���3*�n0WeldW�cial�7�V#Mt�Op����1y�֠ 2F�a�pocrtN�(�p�T1�`T� �� ��xy]ֹ&TX��tw�ig�j�1� b� ct\��JPN ARC?PSU PR��ovݲOL� Sup�2fil� &PAɰא�cro�� "PM�(����O$SS� enвtex�� r����=�t�ssag$T��P��P@�Ȱ�锱�rtW��H'�>r�dpn��n1#
t�!� z ���ascbin4p�syn��+Aj�M� HEL�NCL� VIS PKG�S PLOA`�McB �,�4VW��RIPE GET_VAR FIEo 3\t��FL[��OOL: ADD� R729.FD/ \j8'�CsQ�Q�E��DVvQ�sQNO WTWTE��>}PD  Dp��b�iRFOR ��EC�Tn�`��ALSE� ALAfPCPM�O-130  M�" #h�D: H�ANG FROM�mP�AQfr��R7�09 DRAM �AVAILCHE�CKSO!��sQVP�CS SU�@LIMCHK Q +P~d�FF POS��F��Q R593�8-12 CHA�RY�0�PROGR�A W�SAVE�N`AME�P.SV2��7��$En*��p�?FU�{�TRC|� �SHADV0UPD�AT KCJўRS�TATI�`�P M�UCH y�1��I�MQ MOTN-�003��}�ROB�OGUIDE DAUGH�a���*�Gtou����I� Š�hd�ATH�PepM�OVET�ǔVM�XPACK MA�Y ASSERT��D��YCLfqTA��rBE COR �vr*Q3rAN�pR�C OPTION�SJ1vr̐PSH�-171Z@x�tcǠSU1�1Hp^9R!�Q�`_T�P��'��j�d{tby app wa 5IҌ~d�PHI���p�aT�EL�MXSPD' TB5bLu 1��U�B6@�qENJ`CEV2�61��p��s	�may n�0� �R6{�R� �Rtr�aff)�� 40�*�p��fr��sy�svar scr� J7��cj`DJ�U��bH V��Q/��PSET ERR�`J` 68��PN�DANT SCR�EEN UNRE�A��'�J`D�pPA��pR`IO 1����PFI�pB�pG/ROUN�PD��G���R�P�QnRSVIP� !p�a�PDIGI?T VERS�r}B�Lo�UEWϕ P�06  �!��MA�Gp�abZV�DIx�`� SSUE��ܰ�EPLAN {JOT` DEL�p�ݡ#Z�@D͐CAsLLOb�Q ph���R�QIPND��I{MG�R719���MNT/�PES ��pVL�c��Holp�0Cq���tPG:�`:C�M�canΠ���pg.v�S: 3�D mK�view� d�` �p��eat7У�b� of �P�y���ANNOT �ACCESS M���Ɓ*�t4s a��lok��Fle�x/:�Rw!mo?�PA?�-�����`~n�pa SNBPJ AUTO-�0�6f����TB��PIA�BLE1q 636>��PLN: RG$��pl;pNWFMD�B�VI���tWIT� 9x�0@o��Qu�i#0�ҺPN RR�S?pUSB�� t� & removb�@ )�_��&AxEP7FT_=� 7<`�p�P:�OS-14;4 ��h s�g���@OST� � C�RASH DU �9��$P�pW�� .$��LOGI�N��8&�J��6b0�46 issue� 6 Jg��: �Slow �st~��c (Hos`��c���`IL`IMP�RWtSPOT:Wqh:0�T�STYW =./�VMGR�h��T0CAT��hosB��E�q��� �uO�S:+pRTU' �k�-S� ����E:���pv@�2�� t\�hߐ��m ��al�l��0�  $�H� �WA͐��3 CN�T0 T�� Wr}oU�alarm���0s�d � �0SE1����r R{�OMEpBp���K� 55��REàSEst��g�     �KoANJI�no����INISITA�LIZ-p�dn1we�ρ<��dr�� l�x`�SCII L��fails w��� ��`�YSTE�a���o��Pv� IItH���1W�Gro>P�m ol\wpSh�@�P��Ϡn cfslxL@АWRI ЏOF Lq��p?�F��up��de-r�ela�d "A�Po SY�ch�Ab�etwe:0INDc t0$gbDO����r� `�Gig�E�#operab[ilf  PAbHi�xH`��c�lead�\etf�Ps�r��OS 030�&: f{ig��GLA )P� ��i��7Np t�pswx�B��If��g������5aE>�a EXCE#dU��_�tPCLOS��"�rob�NTdpF�aU�c�!���PNIO V750�Q�1��Qa��DB Ė�P M�+P�QED��DET��-� \�rk��ONLINEhSBUGIQ ߔXĠi`Z�IB�S a�pABC JAR�KYFq� ���0MSIL�`� R�pNД� �p0GAR��D�*pR��P�"! jK�0cT�P�Hl#n��a�ZE V�� TwASK�$VP2(��4`
�!�$�P�`WI[BPK05�!FȐ�B/��BUSY oRUNN�� "��ȁ����R-p�LO��N�DIVY�CU9L��fsfoaBW�p���30	�V��ˠIT`�a5�05.�@OF�UGNEX�P1b�af�@��E��SVEMGN� NMLq� D0pCC_SAFEX �0c�08"qD �PE�T�`N@�#J87�����RsP�A'�M��K�`K�H G�UNCHG۔MEKCH�pMc� T� � y, g@�$ ORY LEAKA8�;�ޢSPEm�Ja:��V�tGRIܱ��@�CTLN�T�Rk�FpepR�j506�EN-`IN������p �`�Ǒk!��Tq3/dqo�STO�0)A�#�L�p �0�@�Q�АY�&�;pb1CTO8pP�s���FB�0@Yp`�`DU��a!O�supk�t4 � PЙF� Bnf�Q�PSVGN-1��V�S'RSR)J�UP��a2�Q�#D�q l �O��QBRKCTR5Ұ�|"-�r�<p�c�j!INVP�D ZO� ��T`h#�Q�cHset,|D��"DUAL� w�2*B�RVO117 A�]�TNѫt�+bTa2�473��q.?��r��{1 009.fd|8�y`j604.\P�-�`hanc�U�� F��e8�� 	 ��npJtPd!q��`���� 5h596p�!5d�� "p�P�P�Q�0�P2�p�A� \P���R(}\\Pe� aʰI���E��1��p�� j  �� ,e�D'p� �A�A\P�q\ 5 sig��a��"AC;a��
�b�Ce\Pb_p��.p�c]l<bHbcb_c�irc~h<n�`tl 1�~`\P`o�d\P�b]o2�� �cb�c�i\P>�jupfrm�d\P�o�`exe�a�oFd\Ptped}o��u`>�cptlibxz\P�lcr�xr\P\�b�lsazEd\P_fm �}gc\P�x���o|sp��o�mc(��ob_jDzop�u6�wf���t��wms�1q��s1ld�)��jmc�o\��n��nuhЕ��|st�e��>�pl�qp�iwcck���uvf0uxߒ��lvisn��CgaculwQ
E  `RFciV\PqiP���Data Acq/uisi��nZU�SOR631`��TR�Q_DMCM �2�P�75H�1�P583�\P1��71��59`�5�P57<P\P�Q����(���Q��o� p\P!daq\b�oA��@�� ge�/�etdms�"D�MER"؟,�pgdD���.�m���-���qaq.<᡾\Pm�o��h���f{�oR5�03��MACRO�s, SksaffP�@lR���03�SR�QT(��Q6��1�Q9ӡ��R�ZSh��P\PJ6+43�@7ؠ6�P�@�PRS�@���e �Q��UС PIK�Q5?2 PTLC�W���\P3 (��p/O ��!�Pn �\P5���03\sfmn�mc "MNMCPq�<��Q��\$AcX�FM���ci,Ҥ�X�����cdpq+�
�sk��SK�\P�SH5�60,P��,�y�r�efp "REF�p�d�A�j\P	�of��OFc�<gy�to��TO_����ٺ����+je�u��caxis2�\PE�\�}e�q"ISDTc�|�]�prax ���MN��u�b�is�de܃h�\�iR\P!� isbasic���B� P]��QA7xes�R6�������.�(Ba�Q�ess��\P���2�pD�@�z�atis�� ��(�{�����~��m��FMc�u�{�
���MNIS��ݝ�� ��x����ٺ��jW�75��Devic��� Interf�ac�RȔQJ75a4��� \P�Ne` ��\P�ϐ2�б�����dn� "DN�E���
tpdnui5UI��ݝ	�bd�bP�q_r�sofOb
dv_aro��u��|���stchkc���z	 �(}on1l��G!ffL+H��J(��"l"/�n��b��z�hamp���T�C�!i�a"�5�9��S�q��0 (��+P�o�u�!2��xp}c_2pcchm�ЏCHMP_�|8бp�evws��2쳌p�csF��#C Se=n\Pacro�U���-�R6�Pd�\Pk�����p��gT�L��1d M�2`��8�1c4�ԡ�3 qem��G�EM,\i(��Dgesnd�5���H{�}H�a�@sy���c�Is1u�xD��Fmd��I���7�4���u���AccuCal�P�4t@���ɢ7ޠB0��6j+6f�6��99\aFF q�S(�U��2�
�X�p�!Bd��cb�_�SaUL��  ��t@?�ܖto��o�tplus\tsCrnغ�qb�Wp���t���1��Tool� (N. A.)0�[K�7�Z�(P�m� ���bfclst@k94�"K4p��q�tpap� "P�S9H�stpsw�o��p�L7��t\ �q����D�yt5�4�q���w�q��t@�M�uk��rkey����s���}t�sfeatu6�EA��t@cf)t�\Xq�����d�h5���LRC0�md��!�587���aR�( ����2V��8c?u3l\�pa3}H�&r-�Xu���t,�t@�q "�q�Ot��~,����{�/��1c�}����y �p�r��5���S�XA�g�-�y���Wj87�4�- iRViys���Queu� t@Ƒ�-�6�1���	(����u���tӑ�����
�tpvtsn "VTSN�3�C�+�t@v\pRDVx����*�prdq\�yQ�&�vstk=P0������nm&_����clrqν���get�TX��Bd��aoQϿ�0qst!r�D[t@��t�p'Z�����npv��@�enlIP0��D!x�'��|���sc ߸��tvo/��2�q���vb����q���!����h]��(� Co�ntrol�PR�AX�P5��556l�A@59�P56.@�56@5A�J6�9$@982 J552 IDVR7� hqA���16�H���La�� ��Xe��frlparm.�f�FRL�am0��C9�@(F�����w6{���A��QJg643�t@50�0�LSE
_pVA�R $SGSYS�C��RS_UNITS �P�2�4tA��TX.$VNUM?_OLD 5�1�| {�50+�"�`? Funct���5@tA� }��`#@�`3�a0�cڂ��9���@�H5נt@�P���( �A����۶}����0ֻ}��bPRb�߶�~ppr4�TPSP`I�3�}�r�10�#@;A� t�
`���1����96�����%C��� Aف��J�bIncr�	����\���1�o5qni4�MNINp	�t@���!���Hour  �� 2�2�1 �AAV1M���0 ���TUP ��J�545 ��61�62�VCAM�  (�CL�IO ��R6x�N2�MSC �"P �ST�YL�C�28~ 1�3\�NRE "�FHRM SCH~^�DCSU%�ORSR {b�0�4 �EIO�C�1 j 542� � os| � egist������7�1�MA�SK�934"7 <��OCO ��"%3�8��2����� 0 HB��� 4v�"39N� Re��� �LCHK
%O�PLG%��3"%M7HCR.%MC  ; �4? ��6 dPI��54�s� DSW�%MD� pQ�K!6C37�0�0p"�1��֠"4 �6<27 �CTN K � 5 J���"7��<25�%z/�T�%FRDM� �Sg!��9309 FB( NBA�P� �( HLB  Me�n�SM$@jB( PgVC ��20v�α2HTC�C�TMIL��\@PA�C 16U�hAJ`S9AI \@ELN��<2�9s�UECKy �b�@FRM �b��OR���IPL���Rk0CSXC \���VVFnaTg@�HTTP �!2�6 ��G�@ob�IGUI"%IP�GS�r� H863� qb�!�07r�!34� �r�84 \s`o`! Qx`CC3 Fbr�21�!96 rb�!51 ���!53R% 1!s3!��~��.p"9js VATFUJ775"��pLRu6^RP�WSMjU'CTO�@xT58 F�!80���1XY <ta3!770 ��7885�UOL  GT�So
�{` LCM9 �r| TSS�EfP�6 W�\@CPE `��0VR� l�Q�NL"��@001 oimrb�c3 =�`�b�0���0�`6 w�b-P- R-�b8nn@5EW�b9 �Ҁ�a� ���b�`ׁ�b2� 2000��`3$��`4*5�`5!�c��#$�`7.%�`8 oh605? U0�@�B6E"aRp7� !Pr8 t�a@�>tr2 iB/�1vp�3�vp5 Ȃtr9�Σ�a4@-p�r3 F��r5&�re`Lu��r7 ��r8�U��p9 \h738|�a�R2D7"�)1f��2&�7� �O3 7iC��4>wq5Ip�Or60 CҲL�1bEN�4 I�p�yL�uP��@N�-PJ�8�N�8NeN�9 PH�r`�E�b7]��|���8�Вࠂ9 �2��a`0�qЂ5~�%U097 0��@1�0���1 (<�q�3 5R��� �0���mpU��0�0�7*�H@(q�\P�"RB6�q124��b;��@���@06l� x�3 pB/x��u ��x�6 H60�6�a1� ��7 �6 ���p�b1�55 ����7jUU�162 �3 �g��4*�65 2�e "_��P�4U1H`���B1���`0'�174 �q��P�E?186 R ��P��7 ��P�8&�3 }(�90 B/�s�191����@202��6 3���A��RU2� d��2 �b2h`��4�᪂2��4���19v Q�2T��u2d�Tpt2� ���H�a2hP�$�5����!U2�p�p
�2�p��@5�0-@��i8 @�9��TX@�t� �e5�`rb26Af�2^R�a�2Kp��1Dy�b5Hp�`
�5��0@�gqGA���a52hѐ�Ḳ6�60ہ)5� ׁ2��8�E��M9�EU5@ٰ\�qQ5hQ`S�2ޖ5�p\w�۲�pJ �-P��M5�p1\t�H�4���PCH�7j��phi�w�@��P�x��559 ldu� P�D��@�Q�@������� �`�.��P>��8�58�1�"�q58�!AM�۲T�A iC�a5�89��@�x����5 �a��12׀0.�1���,�2����,�!P'\h8��Lp ��,��7��6�0840\�t� "T20C�}A��p��{��ran��FRA��Д� �е���A%���ѹ� �Ҁ�����(����� ����З�������� �р����$�G��1�Čը���������� ,e�`q� c �����`64���M��iC/50T-H������*��)p46��� C��N�����m75s֐� 1Sp�ѯb46��v�x���ГM-71?�a7�З����42������C��-�а�7�0�r�E��/h ����O$��rD���c7c7C�q�䈀Ѕ���L��/��2\imm7c7�@g������`��� (��e�����"�������a r��c�T	,�Ѿ�"��,�� ���x�Ex�m77t ���k���5������)�iC��-HS -� B
_�>���+�Т�7U�]���TMh7�s��7�������-9?�/260L_������Q�������]�9pA/@���q�S�х���h�621��c��92�������.�)92c0�g$�@������)$��5$���pylH"O"
�21���t?�350�����p��$�
�� �350!���0��9��U/0\m9��M9�A3��4%� s"�3M$��X%u���"him98J3����� i d�"m4~�10�3p�� �Ӏ�h79!4̂�&R���H�0�� ��\���g�5A���� ���0���*2��00��#06�АՃ�,�է!07{r ��� �����kЙ@����EP�#�������?��#!�;&07\;!�B1P�߀A��/ЁCBׂ2�!�:/�p�?�ҽCD25L�����0�"l�2�BL
#��B��\20 �2_�r�re���X���1��N����A@��z��`C�pU��`F�04��DyA�\�`fQ��sU����\�5  ���; p�Dp���<$�85���+P=�ab;1l�1LT��lA8�!uDnE(�2�0T��J�1 e�bHC85���b�Հ�5[�16Bs���������d2��x��m6t!`Q����bˀ��8�b#�(�6iB;S�p �!��3� ��b�s ��-`�_�W8�_�L���6I	$�X5�1��U85��R�p6S ����/�/+q�!�q��`�6o��5m[o)�m6sW��Q�?��set06p ��3%H�5��10p$�����g/�JrH���  ��A�85!6����F�� ���p/2��� ��܅�✐)�5��̑v��(�&�m6��Y�H�ѝD̑m�6�Ҝ��a6�DM����-S�+��H2�����Ҽ�� �r ̑��✐��l���p1���F���2��\t6h T6H ����Ҝ�'Vl�� �ᜐ�V7ᜐ/����
;3A7��p~S��������4�`圐�V����!3��2�PM�[��%ܖO�chn��vel5����Vq���_arp#��̑��.���2l_hempq$�.�'�6415� ��5���?����F�����5g�L�ј[���!1��𙋹1����M7NU�М��e(ʾ����uq$D;��B-�4��3&H�f�c�� ��h������u� ��㜐��ZS�!ܑL4���M-����S�$ ̑�ք �� 0��<�p����07shJ�H�v�À�sF��S*� ������̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(U L�&�(�,���0�\�?����̑�a�� ,e����a�e�w��2��(�	�2�C��A/���\�+p������21 (ܱ�CL S����B̺��7FГ��?�<�lơ1L@����c� ���u9�0����e/q��O���q9�K��r9 (�� ,�Rs�ז�5�G�m20c��i��w�2��:�0`�$��2 �2l�0�k�X�S� ,�Bι2��O���1!�41w���2T@� _std��G�y� ��x��H� jdgm�� ��w0\� �1L���	� P�~�W*�b��t �5������3�,���E{�������L��5\L��3 �L�|#~���~!���4�#��O����h�LA6A�������2�����44�����>[6\j4s��·����#��ol�E"w�8 Pk�����?0xj�H1��1Rr�>��]�2aF�2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l���0�&�"��|�`Am1��2��ػ��3�HqB ��K�R��ˑb� W���Fs���)�ѐ�@!���a�1����5��;16�16C��xC����0\imBQ@��d����b��\B5�-���DiL���O� _�<ѠPEtL�E�R�H�ZǠPgω�am1l��u���̑�b�<����<�$�T�̑�F ����Ȋ�Dpb��X�"��hr��p� .��Dp���9�0\�� j971\kc/krcfJ�F�s������c��e "CTME�r���ɛ��a�`main.[��g��`run}�_vc �#0�w�1Oܕ_u��<��bctme��Ӧx�`ܑ�j735��- KAREL /Use {�U���AJ��1���p� Ȗ�9�B@��L�9���7j[�atk208 "K��Kя�
�\��9��a��̹8����cKRC�a�o ��kc�qJ�&s�� ���Grſ�fsD��:`y��s��A1X\j|�&�rdtB�, ��`.v�q�� �sǑIf\�Wfj52�TKQuto Set���J� H5K53M6(�932���91�K58(�9�BA�1(��74O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v����! conre�;a#�Contro�l Re�ble��CNRE(�T�<р4�2���D�)���S�5�52��q(g�� (�򭂯4X�cOux�\�sfuts�UTAS`�i�栜���t�棂��? 6�T�!�GSA OO+D6� ��������,!���6c+� igt�t6�i��I0�TW8` ���la��vo58�o��bFå򬡯i�Xh���!Xk�0Y!8\m;6e�!6EC���v��6���������B<16�A���A�6s� ���U�g�T|ώ����r1�qR��˔Z4 �T�����,#�eZp)g����<ONO0���uJ��tCR;��F�a�� ,e��f��pr?dsuchk �1"��2&&?���t��*D%$�r(�✑�娟:r��'�s�qO��<�scrc�C�\At�trldJ"o�\��V����Paylo>�nfirm�l�!�87��7��A�3ad�! �?ވIЯ?plQ��3��3"0�q��x pl�`��p�d7��l�calC��uDu���;��mo�v�����initX�:s8O��a�r4 ���r67A4|�e �Generati�ڲ���7g2q$��g{ R� (Sh��$�c ,|�bE��$Ԃ�\�:�"��4b��4�4�. sg��A5�F$d6"e;Qp "SHAP��TQ ngcr pG�C�a(�&"� ��"gGDA¶��r6��"aW�/�$dat�aX:s�"tpadx��[q�%tput;a __O7;a�o8�1�yl+s�r�?�:�#�?�5Ix�?�:c O�:y O��:�IO�s`O%g �qǒ�?�@0\��"o��j92;!�Ppl.�Collis�QSkip#��@5��@J� �D��@\ވ�C@XJ�7��7�|s2���ptcls�LS��DU�k?�\_ ects�`�< \�Q ��@���`dcKqQ�FC;��J,�n��`# (��4eN����T�{���'j(�c �����/IӸaȁ��̠�H�����зa��e\mcclm?t "CLM�/�¾� mate\��lmpALM�?>p�7qmc?����2vm��q��%�3s��_svx90�_x_msu�2�L^v_� K�o�{i�n�8(3r<�c_l�ogr��rtr)cW� �v_3��~yc��d�<�te���der$cCeN� Fiρ�R���Q�?�l�ent�er߄|��(Sd���1�TX�+fK�r�a99sQ9+�5��r\tq\� "F�NDR����STDn$LA�NG�Pgui��D�⠓�S������sp�!ğ֙uf�ҝ�s ����$�����e+�=� ��������������<w�H�r\fn_�ϣ���$`x�tcpma>��- TCP���~��R638 R�X�Ҡ��38��M7p,���Ӡ�$Ӡ�8p0а��VS,�>�tk��99�a��B3���PզԠ`��D�2�����UI�� t���hqB���8�����0���p���re�ȿ��exe@4φ�B�ࠓe38�ԡG�rmp8WXφ�var@�π��3N�����vx�!�ҡ��q�RBT� $cOPTN? ask E0�Ӿ1�R MAS0�H�593/�96 HY50�i�480�5�!H0��m�Q�K��7�
0�g�Pl�h0ԧ�<2Ҧ�DP��@"���t\mas��0��a��"�ԧ�����k@�գR����ӹ`m�՘b��7�.f��u�d���r��spla�yD�E���1w�UP�DT Ub��887� (��Di{���v �Ӛ�Ԛ⧔��#�B���㟳��o  �@���a�䣣��60q���B����qscaan��B���ad@�������q`�䗣��#��К�`2�� vlv��Ù�$�>�b����! S��Ea�sy/К�Util���룙�511 JȘ����R7 ��No�r֠��inc),(<6Q�� �`c��"84�[���986FVR�x So����q�nd6����P��4�a\ �(��
  �������d���K�bdZ���meyn7���- Me`CtyFњ�Fb�0�8TUa�577?Ai3R��\�5�u?��!� n���f�x�����l\mh����űE|hmn�	��<\O����e�1�� l!��y(��Ù�\|p����0�B���Ћmh�@�� :.aG!���/� t�55�6�!X�l�.�us��Y/k)ensSubL���eK�h��  �B\1;5g?y?�?0�?D��?*rm�p�?Ktbox O2K|`?�G��C?A%ds��0�?�P"�!� �TR ��/��P�T6@�`�U�P(�V�P�Ue�P0�U�PO��\3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?�Ă�Q3t.�P׀al���P+OP51�7��IN0a��Q(8}g��PESTf3u�a�PB�l�ig�h�6��aq��P � s,e��`  n��0mbumpP�Q969g�69�Qq��P�0�baAp�@Q� �BOX��,>vchqe�s�>vetu㒼�=wffse�3� ��]�;u`aW��:z#ol�sm<ub�a-��]D�K�ibQ�c���p�Q<twaǂ tp�Q�҄Taror ROecov�b�O�P�642����a�0q��a⁠QErǃ�QCry��`�P'�T�`��aar������	{'�p�ak971��71���m���>��`jo@t��PXc��C�1�adb� -�ail��na�g���b�QR629��a�Q��b�P  ?�
  �P���$$CL[q O����������$�PS_DI�GIT���"�!�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����*�璬1:PROD�UCT�Q0\PGSTK�bV,n��99�����$FEAT_I�NDEX��~������I�LECOMP ;��)��"���SETUP2 �<��� � N !�_AP2BCK 1=�?  �)}6/"E+%,/i/��W/ �/~+/�/O/�/s/�/ ?�/>?�/b?t??�? '?�?�?]?�?�?O(O �?LO�?pO�?}O�O5O �OYO�O _�O$_�OH_ Z_�O~__�_�_C_�_ g_�_�_	o2o�_Vo�_ zo�oo�o?o�o�ouo 
�o.@�od�o� ��M�q�� �<��`�r����%� ��̏[�������!� J�ُn�������3�ȟ W������"���F�X� �|����/���֯e� �����0���T��x� �����=�ҿ�s�π��,ϻ�9�b�� P�/ 2) *.cVRiϳ�!�*�����������PC��7�!�FR6:D"�c��χ��T� �߽�Lը��ܮx���*.F��>� �	N�,�k��ߏ��STM �����Q������!�iPe�ndant Pa'nel���H��F����4������GIF�������u����JPG&P��<�����	PAN?EL1.DT�́������2 �Y�G��
3w�����//�
4�a/�O///��/�
TPEIN�S.XML�/����\�/�/�!Cus�tom Tool�bar?�PA?SSWORD/�?FRS:\R??� %Passw�ord Config�?��?k?�?O H�6O�?ZOlO�?�OO �O�OUO�OyO_�O�O D_�Oh_�Oa_�_-_�_ Q_�_�_�_o�_@oRo �_voo�o)o;o�o_o �o�o�o*�oN�or ��7��m� �&���\����� y���E�ڏi������ 4�ÏX�j�������� A�S��w�����B� џf�������+���O� ��������>�ͯ߯ t����'���ο]�� ���(Ϸ�L�ۿpς� Ϧ�5���Y�k� ߏ� $߳��Z���~�ߢ� ��C���g�����2� ��V����ߌ���?� ����u�
���.�@��� d������)���M��� q�����<��5r �%��[� &�J�n� �3�W���"/ �F/X/�|//�/�/ A/�/e/�/�/�/0?�/ T?�/M?�??�?=?�? �?s?O�?,O>O�?bO �?�OO'O�OKO�OoO �O_�O:_�O^_p_�O �_#_�_�_Y_�_}_o�_�_Ho)f�$FI�LE_DGBCK� 1=��5`��� (� �)
SUMM?ARY.DGRo�\OMD:�o�o
`�Diag Su�mmary�o�Z
CONSLOG�o��o�a
J�aCo�nsole lo�gK�[�`MEMCHECK@'�o��^qMemor?y Data��W߁)�qHADOW���P��s�Shadow ChangesS��-c-��)	F�TP=��9����w�`qmment T�BD׏�W0<�)�ETHERNE�T̏�^�q�Z��a�Ethernet� bpfigura�tion[��P��DCSVRFˏ��Ï�ܟ�q%�� v�erify alylߟ-c1PY���DIFFԟ��̟a���p%��dif!fc���q��1X�?�Q�� ����{X��CHGD��¯ԯi��px��� �¤�2`�G�Y�� 1��� �GD��ʿ�ܿq��p���Ϥ�F�Y3h�O�a��� 1��(�GD���ψ��y��p�ϡ�0��UPDATES.��Ц��[FRS:�\�����aUpd�ates Lis�t���kPSRBW�LD.CM.��\���B��_pPS_R?OBOWEL���_ ����o��,o!�3��� W���{�
�t���@��� d�����/��Se �����N�r � =�a�r �&�J���/ �9/K/�o/��/"/ �/�/X/�/|/�/#?�/ G?�/k?}??�?0?�? �?f?�?�?O�?OUO �?yOO�O�O>O�ObO �O	_�O-_�OQ_c_�O �__�_:_�_�_p_o �_o;o�__o�_�o�o $o�oHo�o�o~o�o 7�o0m�o� � �V�z�!��E� �i�{�
���.�ÏR� ���������.�S�� w������<�џ`��� ���+���O�ޟH��� ���8���߯n����$FILE_��{PR��������� ��MDONLY 1�=4�� 
 ���w�į��诨�ѿ �������+Ϻ�O�޿ sυ�ϩ�8�����n� ߒ�'߶�4�]��ρ� ߥ߷�F���j���� ��5���Y�k��ߏ�� ��B�����x����1� C���g������,��� P���������?���Lu�VISBC�KR�<�a�*.V�D|�4 FR:�\��4 Vi�sion VD file� :L bpZ�#��Y �}/$/�H/�l/ �/�/1/�/�/�/�/ �/ ?�/1?V?�/z?	? �?�???�?c?�?�?�? .O�?ROdOO�OO�O ;O�O�OqO_�O*_<_ �O`_�O�__%_�_��MR_GRP 1�>4�L�UC4�  B�P	 �]�ol`�*u����RHB� ��2 ���� ��� ��� He�Y�Q`orkbIh�o�Jd�o�Sc�o�oL�ЊJe?JI��9F�5U�a�Q���o�o �D�	�G��aE�9��o9cݨ>���F}@MZ}@Q�۸lr?7T@N�I�@O؁}E�� F@ �r��d�a}J��NJ�k�H9�H�u��F!��IP�s}?�`�.�9�<9��896C'�6<,6\b��}A+~�BS/��B� JA���?B#�VA�4�. �"7�A��_B|EDA����A�a�A������,.��PA� ����|�ݏx���%������4,AX4�P@#x�@ICm4���j�����ǟ ���֟��!��E�`�r�UBH�P p�a`�M�H��o"K�豯ï�T
6�PS@�PS�d˯�o�o�B��P5���@�33@���4�m�T��UUU��U�~w�>u.�?!x��^��ֿ���3��=�[z�=�̽=�V6<�=�=�=$q��~���@8�i7�G��8�D�8@9!�7���@Ϣ���:t�@ ?D�� Cϫo��+C��P��P'�6� �_V� m�o��To��xo �ߜo������A�,� e�P�b������� ������=�(�a�L� ��p���������.��� ����*��N9r] ������� �8#\nY�} �������/ԭ //A/�e/P/�/p/�/ �/�/�/�/?�/+?? ;?a?L?�?p?�?�?�? �?�?�?�?'OOKO6O oO�OHߢOl��ߐߢ� �O�� _��G_bOk_V_ �_z_�_�_�_�_�_o �_1ooUo@oyodovo �o�o�o�o�o�o Nu��� ������;�&� _�J���n�������ݏ ȏ��%�7�I�[�"/ �描�����ٟ���� ���3��W�B�{�f� ������կ������ �A�,�e�P�b����� ���O�O�O��O�O L�_p�:_�����Ϧ� �������'��7�]� H߁�lߥߐ��ߴ��� ����#��G�2�k�2 ��Vw��������� ��1��U�@�R���v� ������������- Q�u���r� �6��)M 4q\n���� ��/�#/I/4/m/ X/�/|/�/�/�/�/�/ ?ֿ�B?�f?0�B� �?f��?���/�?�?�? /OOSO>OwObO�O�O �O�O�O�O�O__=_ (_a_L_^_�_�_�_�� �_��o�_o9o$o]o Ho�olo�o�o�o�o�o �o�o#G2kV {�h����� ��C�.�g�y�`��� �������Џ��� ?�*�c�N���r����� ���̟��)��M� _�&?H?���?���?�? �?����?@�I�4�m� X�j�����ǿ���ֿ ����E�0�i�Tύ� xϱϜ���������_ ,��_S���w�b߇߭� ���߼�������=� (�:�s�^����� �����'�9� �]� o����~��������� ����5 YDV �z������ 1U@yd� �v�����/Я*/ ��
/�u/��/�/�/ �/�/�/�/??;?&? _?J?�?n?�?�?�?�? �?O�?%OOIO4O"� |OBO�O>O�O�O�O�O �O!__E_0_i_T_�_ x_�_�_�_�_�_o�_ /o��?oeowo�oP��o o�o�o�o�o+= $aL�p��� ����'��K�6� o�Z������ɏ��� �� ��D�/ /z� D/��h/ş���ԟ� ��1��U�@�R���v� ����ӯ������-� �Q�<�u�`���`O�O �O���޿��;�&� _�J�oϕπϹϤ��� �����%��"�[�F� �Fo�ߵ����ߠo�� d�!���W�>�{�b� ������������� �A�,�>�w�b����� ����������=���$FNO ����\�
F0l} q  FLAG>��(RRM_CHKTYP  ] ���d �] ���OM� _MIN܍ 	���� � � XT SSB_�CFG ?\? �����OTP_�DEF_OW  �	��,IRC�OM� >�$GE�NOVRD_DO��<�lTHR֮ d�dq_E�NB] qRA�VC_GRP 19@�I X(/  %/7//[/B//�/ x/�/�/�/�/�/?�/ 3??C?i?P?�?t?�? �?�?�?�?OOOAO�(OeOLO^O�OoRO�U�F\� ��,�B,�8�?���O�O�O	__>���  DE_�Hly_�\@@m_B�=��vR/��I�O�SMT
�G�SUoo&o�RHOSTC�19H�I� ��zM�SM�l[�bo�	127.�0�`1�o  e �o�o�o#z�oF�Xj|�l60s	a�nonymous��������(ao�&�&��o� x��o������ҏ�3 ��,�>�a�O���� ������Ο�U%�7�I� �]����f�x����� ���ү����+�i� {�P�b�t�������� ����S�(�:�L� ^ϭ�oϔϦϸ���� ��=��$�6�H�Zߩ� ��Ϳs���������� � �2���V�h�z�� �߰���������
�� k�}ߏߡߣ���߬� ��������C�*< Nq�_����� �-�?�Q�c�eJ�� n������ �/"/E�X/j/|/ �/�/�%'/? [0?B?T?f?x?��? �?�?�?�??E/W/,O�>OPObO�KDaENT� 1I�K P!�?�O   ��O�O �O�O�O#_�OG_
_S_ ._|_�_d_�_�_�_�_ o�_1o�_ogo*o�o No�oro�o�o�o	�o -�oQu8n� �������#� �L�q�4���X���|� ݏ���ď֏7���[����B�QUIC�C0��h�z�۟��1 ܟ��ʟ+���2,����{�!ROUT�ER|�X�j�˯!�PCJOG̯���!192.16?8.0.10��}GNAME !�J!ROBOT��vNS_CFG 1�H�I ��Auto-st�arted�$FTP�/���/�?޿ #?��&�8�JϏ?n� �ϒϤ�ǿ��[����� �"�4ߵ&�������� ��濜���������� '�9�K�]�o���� ����������/�/�/ G���k��ߏ������� ������1T��� Py�����"� 4�	H-|�Qcu �VD���� /�;/M/_/q/�/� ���/
/�/>?%? 7?I?[?*/?�?�?�? �/�?l?�?O!O3OEO �/�/�/�/�?�O ?�O �O�O__�?A_S_e_ w_�O4_._�_�_�_�_ oVOhOzO�O�_so�O �o�o�o�o�o�_ '9Kno�o��� ��o*o<oNoP5� �oY�k�}�����pŏ ׏����0���C�U��g�y���_�T_ER�R J;�����P�DUSIZ  j��^P����>ٕ?WRD ?z����  guest���+�=��O�a�s�*�SCDMNGRP 2Kz�wÐ���۠\��K�� 	�P01.14 8~�q   y���B   � ;����{ ������������������?�����~ �ǟ�I�4�m�X�|���  i  ��  
���� �����+�������
���l��.x����"�l�ڲ۰s�d����|���_GROU��]L�� ��	���۠07K�QUPD'  ���PČ��TYg�����T�TP_AUTH �1M�� <!iPendan����<�_�!K?AREL:*�����KC%�5�G���VISION �SETZ���|�� Ҽߪ��������� 
�W�.�@��d�v���CTRL N��軡���
�F�FF9E3����FRS:DEFA�ULT�FA�NUC Web �Server�
 ������q��������������WR_CONFIG O��� ���IDL_CPU_PC"���B��= �BH#MIN.�B?GNR_IO���� ���% NPT_S_IM_DOs}�TPMODNTO�Ls �_PRT�Y�=!OLNK 1P����'9K]o�MA�STEr �����O�_CFG��UO�����CYCLE����_ASG s1Q���
 q 2/D/V/h/z/�/�/�/ �/�/�/�/
??y"NUM���Q��IPCH��£R?TRY_CN"�u<���SCRN��擊��� ����R����?��$J�23_DSP_E�N�����0OB�PROC�3��J[OGV�1S_�@��?8�?�';ZO�'??0CPOSRE�O�KANJI_@�Ϡu�A#��3T ����E�O�ECL_�LM B2e?�@EYL_OGGIN��������LANGU�AGE _�=e� }Q��LG�2YU����� �x������PC � �'�0�����M�C:\RSCH\�00\˝LN_D?ISP V���0����TOC�4�Dz\A�SOGB?OOK W+��`o���o�o���Xi��o�o�o�o�o~}	x(y��	ne�i��ekElG_BUF/F 1X���}2����Ӣ��� ���'�T�K�]��� ��������ɏۏ����#�P��ËqDCS� Zxm =���%|d1h`���ʟܟ|�g�IO 1[+G �?'����'� 7�I�[�o�������� ǯٯ����!�3�G� W�i�{�������ÿ׿z�El TM  ��d��#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝߜ�t�SEV�0m.�TYP�� �0�$�}�ARS"�(_|�s�2FL 1\��0���������0�����5�TP<P����DmNGNA�M�4�U�f�UPSF`GI�5�A�5s��_LOAD@G �%j%@_M�OV�u����MAXUALRMB7�P8 ��y���3�0]&q
��Ca]s�3�~��� 8@=@^+ �Z�v	��V0+�P1�A5d�r���U����� �E(iTy� ������/ / A/,/Q/w/b/�/~/�/ �/�/�/�/??)?O? :?s?V?�?�?�?�?�? �?�?O'OOKO.OoO ZOlO�O�O�O�O�O�O �O#__G_2_D_}_`_ �_�_�_�_�_�_�_o 
ooUo8oyodo�o�o �o�o�o�o�o�o-���D_LDXDIS�A^�� �MEMO�_APX�E ?��
 �0y� ���������ISC 1_�� �O����W�i� ����Ə�����}� �ߏD�/�h�z�a��� ����������� @���O�a�5������� �����u��ׯ<�'� `�r�Y������y�޿ �ۿ���8Ϲ�G�Y� -ϒ�}϶ϝ�����mπ����4��X�j�#�_MSTR `��~}�SCD 1as}�R���N�������� 8�#�5�n�Y��}�� �����������4�� X�C�|�g��������� ������	B-R xc������ �>)bM� q�����/� (//L/7/p/[/m/�/ �/�/�/�/�/?�/"? H?3?l?W?�?{?�?�?��?n�MKCFG �b���?��LT�ARM_�2cRu;B �3Wp|TNBpMETPUOp��2����NDS?P_CMNTnE@8F�E�� d���N��2A�O�D�EPO�SCF�G�NPS�TOL 1e-�4=@�<#�
;Q�1 ;UK_YW7_Y_[_m_�_ �_�_�_�_�_o�_o Qo3oEo�oio{o�o�a��ASING_CH�K  �MAqODAQ2CfO�7J�e�DEV 	Rz	�MC:'|HSI�ZEn@����eTA�SK %<z%$�12345678�9 ��u�gTRI�G 1g�� l<u%���3����>svvYPaq��kE�M_INF 1h�9G `�)AT&FV0�E0(���)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ���ڄH�� ����G�ֈAO�w� 2�������џ ���� ����͏ߏP��t��� ����]�ί����� (�۟�^��#�5��� ��k�ܿ� ϻ�ů6� �Z�A�~ϐ�C���g� y��������2�i�C� h�ό�G߰��ߩ��� �ϫ��������d�v� )ߚ��߾�y����� ���<�N��r�%�7� I�[������9�& ��J[�g��>�ONITOR�@G� ?;{   	?EXEC1�3�U2�3�4�5�T�p�7�8�9�3�n�R�R�R RRR(R@4R@RLR2YU2e2q2}2�U2�2�2�2�U2�3Y3e3���aR_GRP_SOV 1it��q(�a���C?BPR��A4�>%���gYw>rﳌ"}~q_DCd~�1P�L_NAME �!<u� �!D�efault P�ersonali�ty (from� FD) �4RR�2k! 1j)TE�X)TH��!�AX d�?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�Ox2-?�O�O�O__@0_B_T_f_x_�b<�O �_�_�_�_�_�_o o�2oDoVoho&xRj" �1o�)&0\�b,� �9��b�a �@D�  �a?�ľc�a?�`�a�aA'�6�ew;�	�l�b	 ��xJp���`�`	p �<w �(p� �.r�� K�K ���K=*�J����J���JV�`�kq`q�P�x��|� @j�@T;;f�r�f�q�a�crs�I�����p���p�r�p�h}�3��´  � �>��ph��`z��ꜞ�a��Jm�q� H�N��ac���dw���  �  �P� Q� �� |  а�m�Əi}	'� � ��I� �  �����:�È~�È=���(��ts�a	���I  ?�n @H�i~�ab�Ӌ�b�w���urN0��  '�Ж�q�p@2��@Ǔ���r�q5�C��pC0C�@ C�����`
��A1q) " � @B�V~X�
nwB0h�A��p�ӊa�p�`���aDz����֏���Я	�pv��( �� -��I��-�=��A&�a�we_q�`�p� �?�ff ���m��� �����Ƽuq@ݿ�>N1�  P�apv(�` ţ� �=�qst��/?���`x`�� �<
6b<߈�;܍�<�ê�<� <�&P�ό�AO��c1��ƾ��?fff?O�?y&��qt@�.���J<?�`�� wi4����dly�e߾g ;ߪ�t��p�[ߔ�� �ߣ����� ����6�wh�F0%�r�!�߷�1ى����E��� E�O�G+� F�!���/���?�e�P���t���lyBL�cB��Enw4��� ����+��R��s���������h�Ô�>��I�mXj�F��A�y�weC�p�������#/�*/c/N/wi�����fv/C�`� CHs/�`
=$�p�<!�!������'�3A�A��AR1AO�^?�$�?���5p±
=ç>�����3�W
�=�#�]�;e��׬a@����{�����<��>(�B�u���=B0��?����	R��z�H�F�G����G��H�U`�E���C�+���}I#�I���HD�F���E��RC�j�=�>
I���@H�!H�(� E<YD0 w/O*OONO9OrO]O �O�O�O�O�O�O�O_ �O8_#_\_G_�_�_}_ �_�_�_�_�_�_"oo oXoCo|ogo�o�o�o �o�o�o�o	B- fQ�u���� ���,��P�b�M� ��q�����Ώ���ݏ �(��L�7�p�[��� ���ʟ���ٟ����6�!�Z�E�W���#1(�$1��9�K���<ĥ%����Ư!3�8���!�4Mgs��,�I�B+8�J��a���{�d�d������ȿ���ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ��ϰ�������  %��  ��h�Vߌ�z߰�&ڀg�/9�$������� 7����A�S�e�w�  ��������������2 F��$�&Gb��������!C���@����$����F�� DzN�� F?�P D�������)#B�'9K]�o#?���@@*v
��8�8��u8�.
 v ���!3EW i{����:�� ��ۨ�1���$MSKCFM�AP  ��� ����(.�ONREL  �!9��EXCFENBE'q
#7%^!FNCe/�W$JOGOVLI�ME'dO S"d�K�EYE'�%�R�UN�,�%�S?FSPDTY0g&<P%9#SIGNE/W$�T1MOT�/T!��_CE_GRP� 1p��#\ x��?p��?�?�?�? �?O�?OBO�?fOO [O�OSO�O�O�O�O�O _,_�OP__I_�_=_ �_�_�_�_�_oo�_�:o�TCOM_�CFG 1q	-оvo�o�o
Va_A�RC_b"�p)U?AP_CPL�ot$�NOCHECK {?	+ � x�%7I[m ���������!�.+NO_WAI�T_L 7%S2NT�^ar	+�s�_7ERR_12s	)9�� ,ȍޏ��x����&��dT_M�O��t��, 	��*oq�9�PARAuM��u	+��`a�ß'g{�� =?��345678901��,��K�]�9� i�������ɯۯ��&g������C��cU�M_RSPACE�/�|����$OD�RDSP�c#6p(O�FFSET_CAsRT�o��DISƿ���PEN_FIL�E尨!�ai��`OPTION_IO�/���PWORK 5ve7s# ��V���8� "�ep�4�p��	 ���p��<����RG_DSBL'  ��P#������RIENTTOD ?�C�� !l����UT_SIM_ED$�"���V��?LCT w}���6��a[�1�_PEX9E�j�RATvШ&�p%� ��2^3j)T�EX)TH�)�X d3������ �%�7�I�[�m��� ������������!�3�E���2��u����� ����������c�<d�ASew�� ������Ǎ��^0OUa0o(��_�(����u2, ���O H� @D�  [?��aG?��cc�D�][�Z�;�	�ls��x7J���������< ���� ��ڐH(���H3k7HS�M5G�22G�?��Gp
͜��'f�/-,ڐCR�>�D!�M#{Z/���3�����4y H "�c/u/�/�0B_����=jc��t�!�/ �/�"t32���~�/6  ��UP%�Q%��%�|T���S62�q?'e	'�� � �2I�� �  ��+==��ͳ?�;	��h	�0�I  �n @�2�.���Ov;��ٟ?&gN�]O  ''�uD@!:� C�C�@F#H!��/�O�O sb
�T��@�@��@$�e0@B�QA�0Y�v: �13Uwz $oV_�/z_e_�_�_	���( �� -�2�1�1ta�UDa�c���:A-���~.  �?�ff���[o"o�_U�`oXâ0A8���o�j>�1  Po�V(���eF0��f�Y���L�?˙���xb0@<
�6b<߈;����<�ê<�? <�&�,�/aA�;r�@Ov0P?offf?�0?&ipޘT@�.{r�J<?�`�u#	�B dqt�Yc�a�Mw �Bo��7�"�[�F� �j�������ُ� ���3����,���~(�E�� E��3?G+� F��a�� ҟ�����,��P�(;���B�pAZ�>� �B��6�<OίD���P� �t�=���a�s������6j�h��7o��>�S��O�����Fϑ�A�a�_���C3Ϙ�/�%?��?Ƀ��������#	���P �N||CH����Ŀ������@�I�_�'�3A��A�AR1A�O�^?�$�?������±
=�ç>����3�W
=�#� U���e���B��@���{����<����(�B��u��=B0�������	��b�H�F�G����G��H��U`E���C��+��I#�I���HD�F���E��RC��j=[�
I���@H�!H��( E<YD0߻�������� � �9�$�]�H�Z��� ~�������������# 5 YD}h�� �����
C .gR����� ��	/�-//*/c/ N/�/r/�/�/�/�/�/ ?�/)??M?8?q?\? �?�?�?�?�?�?�?O �?7O"O[OmOXO�O|O �O�O�O�O�O�O�O3_:Q(������b���gUU��xW_i_2�3�8��_<�_2�4Mgs�_�_��RIB+�_�_�a?���{�mi�Go5okoYo�o}l��P'rP�nܡݯ�o=_`�o�_�[R?�Q�u���  �p���o��/�� S��z
uүܠ�������ڱ�����������  /�M�w��e��������l2 wF�$��Gb���t��a�`�p�S�C��y�@p�5�G�Y�۠F�� Dz��� F�P D��]����پ��ʯܯ�� ��~�?��ͫ@@�?�K��K���K���
 �|�������Ŀֿ �����0�B�T�f�ܽ�V� ���{���1��$PARA�M_MENU ?�3�� � DEF�PULSEr�	�WAITTMOU�T��RCV�� �SHELL_�WRK.$CUR�_STYL���	�OPT��PT�B4�.�C�R_DECSN���e��� �ߣ����������� !�3�\�W�i�{����USE_PROG %��%�����CCR���e�����_HOST !F��!��:���T�`�V��/�X����_TIME��^���  ��GDEB�UG\�˴�GINP_FLMSK�����Tfp����PGA�  ����)CH�����TYPE���������� � -?hcu �������/ /@/;/M/_/�/�/�/ �/�/�/�/�/??%?�7?`?��WORD �?	=	RS�fu	PNSU�Ԝ2JOK�DRT�Ey�]TRACE�CTL 1x3���� �`� &�`�`�>�6_DT Qy3�%@~�0D � �co�a:@V�@BR�2ODOVOhOzO�B�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofox`|d�b�h�o�g �m�a�o�o�o�ouJ� }�`M �b5GY~�`F��b�J�tr� ��O�ol���t� #�5��xZ�l�~�P���D\vR��d��N�qf 
��.�@�R�d�v��� ������П����� *�<�N�`�.Iv����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p��j��� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o��o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*���$PGTRACELEN  )��  ���(��>�_UP �z���m��u�Y�n�>�_C�FG {m�W�(�n���PК����DEFSPD �|��'�P���>�IN��TRL +}��(�8�����PE_CONFI���~m���mњ��ղ�LID����=�GRP� 1��W���)�A ���&f�f(�A+33D��� D]� C�O� A@1��Ѭ(��d�Ԭ��0�0�� 	 1�ح֚Ҏ�� ´�����B �9����O�9�s��(�>�T?�
�5�������� =?��=#�
�� ��P;t_�������  Dz (�
H� X~i����� �/�/D///h/S/��/��
V7.1�0beta1���  A�E>�"ӻ�A (�� �?!G��!>���"����!����!BQ��!A\�� �!���!2p����Ț/8?J?\?n?};!� ���/��/�? }/�?�?OO:O%O7O pO[O�OO�O�O�O�O �O_�O6_!_Z_E_~_ i_�_�_�_�_�_�_' o2o�_VoAoSo�owo �o�o�o�o�o�o.�R=v1�/�#F@ �y�}��{m� �y=��1�'�O�a� �?�?�?������ߏʏ ��'��K�6�H��� l�����ɟ���؟� #��G�2�k�V���z� �������o��ί C�.�g�R�d������� ���п	���-�?�*� cώ���Ϯ��� ���B�;�f�x��� ����DϹ��߶����� ���7�"�[�F�X�� |�����������!� 3��W�B�{�f����� ���� �����/ S>wbt��� ���=Oz� �Ͼψ����ϼ�  /.�'/R�d�v߈߁/ 0�/�/�/�/�/�/�/ #??G?2?k?V?h?�? �?�?�?�?�?O�?1O CO.OgORO�OvO�O�O ���O�O�O__?_*_ c_N_�_r_�_�_�_�_ �_o�_)oTfx� to���/�o/ >/P/b/t/mo� |������� 3��W�B�{�f�x��� ��Տ�������A� S�>�w�b����O��џ ������+��O�:� s�^�������ͯ��� ܯ�@oRodo�o`��o �o�o��ƿ�o���* <N�Y��}�hϡ� ���ϰ��������
� C�.�g�Rߋ�v߈��� ������	���-��Q� c�N�ﲟ���l��� �����;�&�_�J� ��n����������� ,�>�P�:L������ ������(�:� 3��0iT�x� ����/�/// S/>/w/b/�/�/�/�/ �/�/�/??=?(?a? s?��?�?X?�?�?�? �?O'OOKO6OoOZO �O~O�O�O�O�O* \&_8_r���_�_���$PLID_�KNOW_M  ���| Q�TSV ����P� �?o"o4o�OXoCoUo��o R�SM_GROP 1��Z'0{`��@�`uf�e�`
�5� �gpk 'Pe]o� ��������V�SMR�c��mT�EyQ}? yR������ ����폯���ӏ�G� !��-����������� 韫���ϟ�C��� )�����������寧����QST�a1 1Ն�)���P0� A 4��E2�D� V�h�������߿¿Կ ���9��.�o�R�dπvψ��ϬϾ����2r�0� Q�<3߂�3�/�A�S��4 l�~ߐߢ��5���������6
��.�@��7Y�k�}���8��������MAD  )���PARNUM  �!�}o+��SCHE� S�
��f���S��UPDf�x���_CMP_0�`H�� �'�U�ER_CHK-����ZE*<RS8r��_�Q_MOG���_�X�_RES_G��!���D� >1bU�y� ����/�	/����+/�k�H/ g/l/��Ї/�/�/� 	��/�/�/�X�?$? )?���D?c?h?�����?�?�?�V 1�x�U�ax�@c]�@}t@(@c\�@}�@D@c[�*@���THR_IN�Rr�J�b�Ud2FM�ASS?O ZSGM�N>OqCMON_QUEUE ��UX�V P~P X�N$ �UhN�FV�@ENqD�A��IEXE�O��E��BE�@�O�CO�PTIO�G��@P�ROGRAM %�J%�@�?���B?TASK_IG�6^OCFG ��Oxz��_�PDATA�c]��[@Ц2=� DoVohozo�j2o�o�o �o�o�o);M^ jINFO[��m��D����� ���1�C�U�g�y� ��������ӏ���	�4dwpt�l )�Q~E DIT ��_|i��^WERFLX�	C�RGADJ ��tZA�����?�נʕFA��IORI�TY�GW���MPGDSPNQ����U�GyD��OTOE@�1�X� (!�AF:@E� c�Ч�!tcpn����!ud����!�icm���?<�XYm_�Q�X���Q)� *�1�5��P��]�@�L���p� �������ʿ��+�@=�$�a�Hυϗ�*��OPORT)QH��P��E��_CAR�TREPPX��S�KSTA�H�
SS�AV�@�tZ	2500H863��P�_x�
�'��X�@�swPtS�ߕߧ�^��URGE�@B��6x	WF��DO�F"�[W\�������WR�UP_DELAY� �X���R_HOTqX	B%�c����R_NORMAL�q^R��v�SEMI������9�QSKI�P'��tUr�x 	7�1�1��X�j� |�?�tU���������� ����$J\n 4������� �4FX|j �������/ 0/B//R/x/f/�/�/��/tU�$RCVT�M$��D�� DC�R'���Ў!?��1�C�k�>��>5F=��� �0r�������A����i�:�o?2? �<
6b<���;܍�>u.��?!<�&�?h?�?�?�@>��? O O2ODOVOhOzO�O �O�O�O�O�?�O�O_ _@_+_=_v_Y_�_�_ �?�_�_�_oo*o<o No`oro�o�o�o�_�o �o�o�o�o8J- n��_����� ��"�4�F�X�j�U ������ď���ӏ� ��B�T��x����� ����ҟ�����,� >�)�b�M��������� ���ïկ�Y�:�L� ^�p���������ʿܿ � ����6�!�Z�E� ~ϐ�{ϴϗ�����-� � �2�D�V�h�zߌ� �߰���������
��� .��R�=�v��k�� ���������*�<� N�`�r���������� ������&J\ ?������� �"4FXj|���!GN_ATC� 1�	; �AT&FV0E�0�ATDP�/6/9/2/9��ATA�,�AT%G1%�B960�+�++�,�H/,��!IO_TYPE'  �%�#t��REFPOS1 �1�V+ x�u/�n�/j�/
= �/�/�/Q?<?u??�?�4?�?X?�?�?�+2 1�V+�/�?�?\O��?�O�?�!3 1� O*O<OvO�O�O_�OS4 1��O�O�O�_�_t_�_+_S5 1�B_T_f_�_o	o|Bo�_S6 1��_��_�_5o�o�o�oUoS7 1�lo~o�o�o�H3l�oS8 1�%_����SMASK 1�V/  
?�M��'XNOS/�r�������!MOTE  �n��$��_CFG �����q���"PL_RANG������POWER �����SM_D�RYPRG %�o�%�P��TAR�T ��^�UME_PRO-�?�����$_EXEC_E�NB  ���GSPD��Րݘ��gTDB��
�RM�.
�MT_'�T�����OBOT_N�AME o�����OB_ORD_NUM ?��b!H863  �կ�����PC_TI�MEOUT�� xޚS232Ă1��� LTE�ACH PENDcAN��w��-���Maint�enance CGons���s�"��~�KCL/Cm�Ț

���t�ҿ No Use-p��Ϝ�0�NPO�\򁋁��.�oCH_L�������q	��s�MAVGAIL�����糅���SPACE1 ;2��, j�߂ �D��s�߂� �{~S�8�?�k� v�k�Z߬��ߤ��ߚ � �2�D���hߊ�|� ��`��������� � �2�D��h��|� ��`���������y���2����0�B��� f�����{���3);M_ ������/� /44FXj |*/���/�/�/?(??=?5Q/c/u/ �/�/G?�/�/�?O�? $OEO,OZO6n?�? �?�?�?dO�?�?_,_@�OA_b_I_w_7�O �O�O�O�O�_�O_(o�Ioo^oofo�o8 �_�_�_�_�_�oo6o Ef){����G �o� t���
M� � ��*�<�N�`�r����� ��w���o�収���d.��%�S�e�w� ����������Ǐَ�� �Θ8�+�=�k�}��� ����ůׯ͟���� %�'�X�K�]������� ��ӿ������#��E�W� `� @�������x�����\�e���������� �R�d߂�8�j߬߾� �ߒߤ���������� 0�r���X�����������8����
��ύ�_MODE�  �{��S E��{|�2�0�����3�	S|)�CWORK_AD޳���+R  �{�`� �� _INTVAL����d���R_OPT�ION� ���H VAT_GRPw 2��upG(N�k |��_���� �/0/B/��h�u/T�  }/�/�/�/�/�/�/ ?!?�/E?W?i?{?�? �?5?�?�?�?�?�?O /OAOOeOwO�O�O�O �OUO�O�O__�O=_ O_a_s_5_�_�_�_�_ �_�_�_o'o9o�_Io oo�o�oUo�o�o�o�o �o�o5GYk- ���u���� �1�C��g�y���M� ����ӏ叧�	��-� ?�Q�c����������� ����ǟ�;�M��_����$SCAN�_TIM��_%�}�R �(�#�((�<04Wd d 
�!D�ʣ��u��/�����U�"�25���@�d5�P�g��]	����������dd�x�  P~���� ��  8� ҿ�!���D��$�M�_�q� �ϕϧϹ��������8ƿv��F��X��/� ;�o�b��pm��t�_DiQ̡  � l�|�̡ ĥ�������!�3�E� W�i�{�������� ������/�A�S�e� ]�Ӈ����������� ��);M_q ������� r���j�Tfx� ������// ,/>/P/b/t/�/�/�/p�/�/�%�/  0�� 6��!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O *�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo �O�OJ�o�o�o�o�o �o�o 2DVh z�������
�7?  ;�>�P� b�t���������Ǐُ ����!�3�E�W�i��{�������ß � ş3�ܟ��&�8�J��\�n�������������ɯ����,�� �+�	12�345678��W 	� =5���@f�x���������� ���
��.�@�R�d� vψϚ�៾������� ��*�<�N�`�r߄� �Ϩߺ��������� &�8�J�\�n�ߒ�� �����������"�4� F�u�j�|��������� ������0_�T fx������ �I>Pbt �������! /(/:/L/^/p/�/�/ �/�/�/�/�2�/�?�#/9?K?]?�i�Cz  Bp˚ /  ��h2��*��$SCR_GR�P 1�(�U8�(�\x�d�@ � ��'�	 ?�3�1 �2�4(1*�&�I3�Fp1OOXO}m��CD�@�0ʛ)���H�UK�LM-10�iA 890?�9�0;��F;�M61�C D�:�CP��1

\&V�1	�6F� �CW�9)A7Y	(R�_��_�_�_�_�\���0i^�oOUO>o Po#G�/���o'o�o��o�o�oB�0ƐrtAA�0* C @�Bu&Xw?���ju�bH0{UzAF?@ F�`�r� �o�����+�� O�:�s��mBqrr����������B�͏b�� ��7�"�[�F�X���|� ����ٟğ���N��� AO�0�B�CU
L���xE�jqBq>7�����$G@�@pϯ BȆ��G�I
E�0E�L_DEFAUL�T  �T���E��MI�POWERFL � 
E*��7�WF�DO� *��1E�RVENT 1����`(�� L�!DUM_EI�P��>��j!AF_INE�¿C�O!FT�����r�!o:� ���a�!RPC_M'AINb�DȺPϭ�Nt�VIS}�Cɻ�����!TP��PU��ϫ�d��E�!
P�MON_PROX	YF߮�e4ߑ��_��f����!RD�M_SRV�߫�g��)�!R�IﰴYh�u�!
v�M���id���!RL�SYNC��>�8|���!ROS��4��4��Y�(�}��� J�\����������� ��7��["4F� j|����!��Eio�ICE_�KL ?%� �(%SVCPRG1n>���3��3���4//�5./3/�6V/[/��7~/�/��D�/�9�/�+�@��/�� #?��K?��s?�  /�?�H/�?�p/�? ��/O��/;O��/ cO�?�O�9?�O� a?�O��?_��?+_ ��?S_�O{_�)O �_�QO�_�yO�_� �Os����>o�o }1�o�o�o�o�o�o�o ;M8q\� �������� 7�"�[�F��j����� ��ُď���!��E� 0�W�{�f�����ß�� �ҟ���A�,�e� P���t��������ί��y_DEV ���MC:����_!�OU�T��2��RE�C 1�`e�j�� � 	��  �������Fg �������̿��Ge��������
 �PSD#6 r�����O��������`D�����`e�����堆�0�  +T^�3���I3��3�!3����^Ͽ�_�^`ePSJ;:��U��?��(�ϋ �������RZ������E3�����
�k���Cl:̠��̒���
^��&�2�D�Vߜ�T�ߌ�":���=��*����؆����Y����-�����
��"3����b���*� �������(��L�:� p���d�����������  ��$ZH~ l�������  VDz�n ������/./ /R/@/b/�/v/�/�/�/}�2��/�/�/? :?(?^?L?�?�?v?�? �?�?�?�?�? O6OO FOlOZO�O~O�O�O�O �O�O_�O2_ _B_h_ V_�_n_�_�_�_�_�_ 
o�_.o@o"odoRoto vo�o�o�o�o�o�o <*`Np�x �������8� J�,�n�\��������� Ə�Ώ�����F�4��j�X���`�p�V 1�}� P����ɿ��$ 
�e �y���TYPE\���HELL_CF�G �.�є��8��}��RS-Ѡ� ����֯������	� B�-�f�Q�c���������������ؐ�%�3�E��Q�)�a��M�o�p�����2��d]�K�:�H�K 1�H�  u�������A�<�N� `߉߄ߖߨ������߀����&�8��=�OMM �H���9��FTOV_ENB�&�1�OW_RE�G_UI��8�IM/WAIT��a���OUT������T�IM�����V�AL����_UNI�T��K�1�MON_�ALIAS ?e~w� ( he�� ����������ж�� );M��q��� �d��%� I[m�<�� ����!/3/E/W/ /{/�/�/�/�/n/�/ �/??/?�/S?e?w? �?�?F?�?�?�?�?�? O+O=OOOaOO�O�O �O�O�OxO�O__'_ 9_�O]_o_�_�_>_�_ �_�_�_�_�_#o5oGo Yokoo�o�o�o�o�o �o�o1C�og y��H���� 	��-�?�Q�c�u� � ������ϏᏌ��� )�;��L�q������� R�˟ݟ�����7� I�[�m��*�����ǯ ٯ믖��!�3�E�� i�{�������\�տ� ����ȿA�S�e�w� ��4ϭϿ����ώ��� �+�=�O���s߅ߗ� �߻�f�������'� ��K�]�o���>�� ��������#�5�G� Y��}���������n���$SMON_D�EFPRO ������� *SYS�TEM*  d=���RECALL� ?}�� ( ��}3copy �frs:orde�rfil.dat� virt:\t�mpback\=�>inspiro?n:3648��r؄�n�}*.mdb:*.*CU
Y����	.x.:\�8R�n��
�/.a6H_^��//�
xyz�rate 61 ����n/�/�/�|.'R6044 H/ Z/�/�/?�-?Q	 �"a?s?�?�?�E?�( Y?�?�?O!3F/�# �?nO�O�O�6OHO�  ^O�O__&?8?�?�? m__�_�?�?�?Z_�_ �_o"O4O�OXOio{o �o�O�OCo�O�o�o _0_B_T_ew��_ �_I�_����,o �oPoa�s������o;� �o`����(:� ޏo��������\� ����$���ɏZ�k� }�������E�؏��� � /2/į֯g�y���|�/�/:5076�/ Y�����!�3����� a�sυϗϪ�EϽ�Y� �����!�3�F�³�� n߀ߒߥ�6�H�Ű^� ����&�8�����m� ��϶���Z����� �"�4���X�i�{��� �߲�C�������� 0�����ew������ 4060ǿY� �!�3��as ����E�Y�� /!�3�F��n/�/ �/��6/H/� ^/�/? ?&8��m??�? ���Z?�?�?O!7��$SNPX_A�SG 1�����9A� �P 0 '%�R[1]@1.Y1O 9?�#3%dO �OsO�O�O�O�O�O�O  __D_'_9_z_]_�_ �_�_�_�_�_
o�_o @o#odoGoYo�o}o�o �o�o�o�o�o*4 `C�gy��� ����	�J�-�T� ��c�������ڏ��� ��4��)�j�M�t� ����ğ������ݟ� 0��T�7�I���m��� �����ǯٯ���$� P�3�t�W�i������� �ÿ����:��D� p�Sϔ�wω��ϭ���  ���$���Z�=�d� ��sߴߗߩ�������  ��D�'�9�z�]�� ��������
���� @�#�d�G�Y���}��� ����������*4 `C�gy��� ���	J-T �c������ /�4//)/j/M/t/ �/�/�/�/�/�/�/?�0?4,DPARAM� �9ECA ��	��:P�4��0$HOFT_K�B_CFG  �p3?E�4PIN_S_IM  9K�6��?�?�?�0,@RVQSTP_DSB�>��21On8J0SR ���:� & �CAR=O~N��6TOP_ON_�ERl@�F�8�AP_TN �5�@�A�BRIN�G_PRM�O �J0VDT_GRP� 1�Y9�@  	�7n8_(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2Dkhz�� �����
�1�.� @�R�d�v��������� Џ�����*�<�N� `�r���������̟ޟ ���&�8�J�\��� ��������ȯگ��� �"�I�F�X�j�|��� ����Ŀֿ���� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�tߛߘߪ߼��� ������(�:�a�^� p�����������  �'�$�6�H�Z�l�~���������������3V�PRG_COUN�T�6��A�5ENB�OM=�4J_UPD 1��;8  
p2� ����� )$ 6Hql~��� ��/�/ /I/D/ V/h/�/�/�/�/�/�/ �/�/!??.?@?i?d? v?�?�?�?�?�?�?�? OOAO<ONO`O�O�O �O�O�O�O�O�O__ &_8_a_\_n_�_�_�_�YSDEBUG�" � �Pdk	�PS�P_PASS"�B?�[LOG ���m�P��X�_  �g�Q
MC:\d�_b_MPCm��o�o��Qa�o �vfS_AV �m:dlUb�U\gSV�\�TEM_TIMEw 1�� (�P�ճTԱXfoT1?SVGUNS} #�'k�spASK_OPTION" �gospBCC�FG ��| q�b�{�}`� ���a&��#�\�G��� k�����ȏ������ "��F�1�j�U���y� ��ğ���ӟ���0��T�f��UR���S� ��ƯA������ �� D��nd��t9�l����� ����ڿȿ����� "�X�F�|�jϠώ��� ����������B�0� f�T�v�xߊ��ߦؑ� ������(��L�:� \��p�������� ��� �6�$�F�H�Z� ��~������������� 2 VDzh� �������� 4Fdv��� ���//*/�N/ </r/`/�/�/�/�/�/ �/�/??8?&?\?J? l?�?�?�?�?�?�?�? �?OO"OXOFO|O2 �O�O�O�O�OfO_�O _B_0_f_x_�_X_�_ �_�_�_�_�_ooo Po>otobo�o�o�o�o �o�o�o:(^ Lnp�����O ��$�6�H��l�Z� |�����Ə؏ꏸ�� ��2� �V�D�f�h�z� ����ԟ����
� ,�R�@�v�d������� ��ίЯ���<�� T�f�������&�̿�� ܿ��&�8�J��n� \ϒπ϶Ϥ������� ���4�"�X�F�|�j� �߲ߠ���������� �.�0�B�x�f��R� �����������,�� <�b�P�������x��� ������&(: p^������ � 6$ZH~ l�������� /&/D/V/h/��/z/��/�/�/�/�&0�$�TBCSG_GR�P 2��%��  �1 
 ?�  /? A?+?e?O?�?s?�?�?��?�?�;23�<_d, �$A?1�	 HC���6>���@E�5CL � B�'2^OjH4J���B\)LFY�  A�jO�MB���?�IBl�O�O�@��JG_�@�  D	 �15_ __$YC-P{_HF_`_j\��_�]@0 �>�X�Uo�_�_6oSo@o0o~o�o�k�h�0�	V3.00~'2	m61c�c	*�`�d2�o�e�>�JC0(�a�i q,p�m-  �0�����omvu1J�CFG ��%e 1 #0vz��rqBr�|�|�� ��z� �%��I�4� m�X���|�������� ֏���3��W�B�g� ��x�����՟����� ���S�>�w�b��� ��'2A ��ʯܯ��� ���E�0�i�T���x� ��ÿտ翢����/� �?�e�1�/���/�� �Ϯ��������,�� P�>�`߆�tߪߘ��� ���������L�:� p�^��������� ��� �6�H�>/`�r� ���������������  0Vhz8� �����
. �R@vd��� ����//</*/ L/r/`/�/�/�/�/�/ �/�/�/?8?&?\?J? �?n?�?�?�?�?���? OO�?FO4OVOXOjO �O�O�O�O�O�O__ �OB_0_f_T_v_�_�_ �_z_�_�_�_oo>o ,oboPoroto�o�o�o �o�o�o(8^ L�p����� ��$��H�6�l�~� (O����f�d��؏� ��2� �B�D�V����� ��n����ԟ
���.� @�R�d����v����� ���Я���*��N� <�^�`�r�����̿�� �޿��$�J�8�n� \ϒπ϶Ϥ������� ߊ�(�:�L���|�j� �߲ߠ���������� 0�B�T��x�f��� �����������,�� P�>�t�b��������� ������:(J L^������  �6$ZH~ l��^���dߚ  //D/2/h/V/x/�/ �/�/�/�/�/�/?
? @?.?d?v?�?�?T?�? �?�?�?�?OO<O*O `ONO�OrO�O�O�O�O �O_�O&__6_8_J_ �_n_�_�_�_�_�_�_ �_"ooFo��po�o ,oZo�o�o�o�o�o 0Tfx�H� ������,�>� �b�P���t������� ��Ώ��(��L�:� p�^�������ʟ��� ܟ� �"�$�6�l�Z� ��~�����دꯔo� �&�ЯV�D�z�h��� ����Կ¿��
��.π�R�@�v�dϚτ� s ���� ��������$TBJO�P_GRP 2����� O ?������������x/JBЌ��9�� �< �zX���� @����	 �C�� >t�b  C����>��͘Րդ��>̚йѳ33=��CLj�ff�f?��?�ffB@G��ь�����t�ц��>�(�\)��ߖ�E噙�;���hCYj��  �@h��B�  A�����f��C� � Dhъ�1���O�4�N����
�:���Bl^���j�i�l�l����A�ϙ�A�"��D��֊=qH������p�h�Q�;��A�j�ٙ7�@L��D	2��������$�6�>B�\p��T���Q�tsx�@33@���C����y�1����>G��Dh�������<���<{�h�@i� ��t� �	���K&� j�n|���p��/�/:/k/�ԇ����!��	V3�.00J�m61cI�*� IԿ��/��' Eo��E��E���E�F���F!�F8���FT�Fqe\�F�NaF����F�^lF����F�:
F�)�F��3G��G��G���G,I�!CH`��C�dTDU��?D��D���DE(!/E\��E��E�h��E�ME���sF`F+'�\FD��F`�=F}'�F���F�[
F����F��M;��;WQ�T,8�4` *Q�ϴ?�2���3�\�X/O��ESTP?ARS  ��	����HR@ABLE� 1����0��D
H�7 8��9
G
H�
H����
G	
H
�
H
HYE��
H�
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_Ht_�^:BS _� �J GoYoko}o�o�o�o�o �o�o�o1CU gy����`#oRL �y�_�_�_�_�O�O�O��O�OX:B�rNUM�  ����P��� V@P:B_?CFG ˭�Z��h�@��IMEBF_TT%AU��2@�GVERS�q���R 1���
 (I�/����b� �� ��J�\���j�|���ǟ ��ȟ֟�����0� B�T���x�������2��_���@�
��M�I_CHAN�� �� ��DBGLV����������ET�HERAD ?*��O�������xh�����ROUT�!��!������?SNMASKD��>U�255.���#������OOLOF/S_DI%@�u.��ORQCTRL �����}ϛ3rϧ� ����������%�7� I�[�:���h�z߯�A�PE_DETAI�"�G�PON_SV�OFF=���P_M�ON �֍�2���STRTCHK� �^�����VTCOMPAT���O�����FPROG� %^�%CA������ISPLA�Y&H��_INST+_Mް �������US�q��LCK����QUICKM�E�=���SCRE�Z�G�tps� ���u�z�����_��@@n�.�SR_�GRP 1�^�/ �O���� 
��+O=sa�쀚�
m���� ��L/C1g U�y����� 	/�-//Q/?/a/�/�	123456�7�0�/�/@Xt�1����
 �}i�pnl/� gen.htm�? ?2?�D?V?`Pan�el setupZ<}P�?�?�?�?�?�? �??,O>OPO bOtO�O�?�O!O�O�O �O__(_�O�O^_p_ �_�_�_�_/_]_S_ o o$o6oHoZo�_~o�_ �o�o�o�o�o�oso�o 2DVhz�1 '���
��.�� R��v���������Џ|G���UALRM��oG ?9� � 1�#�5�f�Y���}��� ����џן���,���P��SEV  �����ECFG ��롽�}A��   BȽ�
 Q���^���� 	��-�?�Q�c�u���Й��������� P�����I��?����(%D�6� �$�]� Hρ�lϥϐ��ϴ��π����#��G���� ��߿U�I_Y�H�IST 1�� � (� ���(/SOFTP�ART/GENL�INK?curr�ent=edit�page,��,1`����(�:�'�����menu��71 �߅����J�=��� ����+�=���a�s� ��������J����� '9����o�� ���X��# 5G�k}������f��f// '/9/K/]/`�/�/�/ �/�/�/j/�/?#?5? G?Y?�/�/�?�?�?�? �?�?x?OO1OCOUO gO�?�O�O�O�O�O�O tO�O_-_?_Q_c_u_ _�_�_�_�_�_�_� �)o;oMo_oqo�o�_ �o�o�o�o�o�o% 7I[m� � ������3�E� W�i�{������ÏՏ �������A�S�e� w�����*���џ��� ��ooO�a�s��� ������ͯ߯��� '���K�]�o������� ��F�ۿ����#�5� ĿY�k�}Ϗϡϳ�B� ��������1�C��� g�yߋߝ߯���P��� ��	��-�?�*�<�u� ������������ �)�;�M�������� ��������l�% 7I[����� ��hz!3E Wi������ �v////A/S/e/�P���$UI_P�ANEDATA �1�����!�  	�}w/�/�/�/�/?? )?>?V�/i?{? �?�?�?�?*?�?�?O OOAO(OeOLO�O�O �O�O�O�O�O�O_&Y� b�>RQ?V_ h_z_�_�_�__�_G? �_
oo.o@oRodo�_ �ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_� �!�3�E�W��{��_ ����ÏՏ���`�� /��S�:�w���p��� ��џ������+�� O�a���������ͯ ߯�D����9�K�]� o��������ɿ��� Կ�#�
�G�.�k�}� dϡψ����Ͼ���n� ��1�C�U�g�yߋ��� ����4�����	��-� ?��c�J����� �����������;�M� 4�q�X��������� ��%7��[�� �����@� �3WiP� t�����/� //A/����w/�/�/�/ �/�/$/�/h?+?=? O?a?s?�?�/�?�?�? �?�?O�?'OOKO]O DO�OhO�O�O�O�ON/ `/_#_5_G_Y_k_�O �_�_?�_�_�_�_o o�_Co*ogoyo`o�o �o�o�o�o�o�o-�Q8u�O�O}���������) �>��U-�j�|����� ��ď+��Ϗ��� B�)�f�M��������� �����ݟ��XS�K��$UI_PAN�ELINK 1��U  ��  ��}�1234567890s���������ͯ դ�Rq����!�3�E� W��{�������ÿտDm�m�&����Qo�  �0�B�T�f�x� �v�&ϲ��������� ߤ�0�B�T�f�xߊ� "ߘ����������� ��>�P�b�t���0� ������������$� L�^�p�����,�>�������� $�0, &�[�XI�m�� �����>P 3t�i��Ϻ � -n��'/9/K/]/ o/�/t�/�/�/�/�/ �/?�/)?;?M?_?q? �?�UQ�=�2"��? �?�?OO%O7O��OO aOsO�O�O�O�OJO�O �O__'_9_�O]_o_ �_�_�_�_F_�_�_�_ o#o5oGo�_ko}o�o �o�o�oTo�o�o 1C�ogy��� ��B�	��-�� Q�c�F�����|����� ��֏�)��M�� �=�?��?/ȟڟ� ���"�?F�X�j�|� ����/�į֯���� �0��?�?�?x����� ����ҿY����,� >�P�b��ϘϪϼ� ����o���(�:�L� ^��ςߔߦ߸����� ��}��$�6�H�Z�l� �ߐ���������y� � �2�D�V�h�z�� ��-���������
�� .RdG��} ����c���< ��`r����� ���//&/8/J/� n/�/�/�/�/�/7�I� [�	�"?4?F?X?j?|? ��?�?�?�?�?�?�? O0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�__�_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o ��6H�l ~a������ ��2��V�h�K��� ����1�U
�� .�@�R�d�W/������ ��П������*�<� N�`�r��/�/?��̯ ޯ���&���J�\� n�������3�ȿڿ� ���"ϱ�F�X�j�|� �Ϡϲ�A�������� �0߿�T�f�xߊߜ� ��=���������,� >���b�t����� +������:�L� /�p���e��������� �� ��6����ۏ��$UI_Q�UICKMEN � ����}��RESTO�RE 1٩��  � 
�8m3\ n���G��� �/�4/F/X/j/|/ '�/�/�//�/�/? ?0?�/T?f?x?�?�? �?Q?�?�?�?OO�/ 'O9OKO�?�O�O�O�O �OqO�O__(_:_�O ^_p_�_�_�_QO[_�_ �_I_�_$o6oHoZolo o�o�o�o�o�o{o�o  2D�_Qcu �o������� .�@�R�d�v�������Џ⏜SCRE�� ?�uw1sc� u2�U3�4�5�6��7�8��USE�R����T���k�s'���4��5��6ʆ�7��8��� ND�O_CFG ڶ�  �  � P�DATE h��None��SEUFRAME�  ϖ��R�TOL_ABRT8����ENB(��?GRP 1��	�Cz  A�~� |�%|�������į֦!��X�� UH�X�~7�MSK  K�4S�7�N�%uT��%�����VISCAND_MAXI��I�3���FAI�L_IMGI�z ��% #S���IMRE/GNUMI�
���gSIZI�� �ϔ�,�ONTMOiU'�K�Ε�&�����(��(���s�FR:�\�� � �MC:\(�\LO�Gh�B@Ԕ !�{��Ϡ�����z? MCV����oUD1 �EX	��z ��PO64�_�Q��n66��PO!�LI�O�䞶e�V�N�f@�`�I�� =	_�S�ZVmޘ��`�W�AImߠ�STAT' �k�% @��4�F�T�$#�x �2�DWP  ���P G��=���͎���_JMPERR 1ޱ�
  �p2345?678901�� �	�:�-�?�]�c��� ��������������$�MLOW�ޘ���Ό�_TI/�˘'���MPHASE � k�ԓ� ��SoHIFT%�1 Ǚ��<z��_ ����F/ |Se����� ��0///?/x/O/ a/�/�/�/�/�/�����k�	VSFT]1[�	V��M+3� �5�Ք p��~��A�  B8[0[0�Πpg3a1Y21�_3Y�7ME��K��͗	6e���&%�J�M���b��	���$��TDINE#ND3�4��4OH�+�G1�OS2OIV I����]LRELE�vI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�YBOX �ǝf_[��b�2�TI190.0.�P�83p\�V25�4p^�Ԓ	 ��S�_�[b���robot84q_ ?  p�9o[�pc�PZoMh��]Hm�_Jk@1�o�ZWABCd��k�,�� �P[�Xo}�o0) ;M�q����@����>��aZ�b��_V