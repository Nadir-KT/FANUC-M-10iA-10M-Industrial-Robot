��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �ET�H_FLTR.�� $�  � �FTP_C�TRL. @ ?$LOG_8	��CMO>$DN�LD_FILTE�� � SUBDIR�CAP� �
��HO��NT. �4� H_NAME� !ADD�RTYPA H_?LENGTH'f �z +LS� D $RO�BOTIG PE�ER^� MASKnMRU~OMG�DEV#���RD�M*�DISA�BL&�TCP�IG/ 3 $A�RPSIZ&_�IPF'W_MC���F_IN� F=A~LASSs��HO_� INFO���TELK �PV�b	 W�ORD  $�ACCESS_L�VL?TIMEO{UTuORT � >�ICEUS= ���$#  �����!�� � � V?IRTUAL�/�!�'0 �%
�*��F�����$�%����+ �����$�� �-�2%;�SHARE�D 1�) � P!�!�?���! |?�?�?�?�?O�?%O �?1OOZOOBO�OfO �O�O�O�O_�O�OE_ _i_,_�_P_�_t_�_ �_�_o�_/o�_Soo Lo�oxo�opo�o�o�o �o�o*Os6 �Z�~���� �9��]� ���D�V� ��z�ۏ����#�� �Y�H�}�@���)7z �_LIST 1�=x!1.ܒ0Ȫ�d�ە1�d�2�55.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H� ��	��-�O�5I��@��o�������O�6����8������ �$���-� ���-@��%�%��&!Ò�)�0H!� ����rj3_tp�d���! � �!!KC� e�0ٙ��&W�!Cm ��w����S�!CON� ��1�=�smo	n��W�