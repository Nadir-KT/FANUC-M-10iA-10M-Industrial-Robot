��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �R  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�H UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2F�G1_�3�B�2G�XD�#
 d� $CARD_�EXIST4$�FSSB_TYP�uAHKBD_S��B�1AGN Gn� $SLOT_�NUMJQPREV,DBU� g1G ;1�_EDIT1 W� 1G=� yS�0%$EP��$OP�~AETE_OKR{US�P_CRQ�$;4�V� 0LACIw1�RAPk �1x@ME@$D�V�Q�Pv�A�{oQL� OUzR� ,mA�0�!� B�� LM_O�^eR��"CAM_;1� xr$AT�TR4NP� ANN��@5IMG_HE�IGHQ�cWID�TH4VT� �U�U0F_ASPEC�Q$M�0EXP���@AX�f�CF�T X $GIR� � S�!�@B@�NFLI�`t� U�IRE 3dTuGITSCHC�`N� S�d�_L�`�C�"�`EQDlpE� J�4S�0@� �zsa�!ip;G0� � 
$WARNM�0f�!,P� ܁s�pNST� CO�RN�"a1FLTR^�uTRAT� T�p; H0ACCa1�p��{�ORI
`l"S={RT0_S�BְqHG,I1 E[ Tp�"3I9�CTY�D,P*2 �`�w@� �!R*HD��cJ* C��2��3���4��5��6��7ʳ�8��94���CO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS�`�}Aw��"�tP_*0wOFSzR @� �RO_K8���aIT<�3��NOM_�0�1iĥ3FCPT� �� $���AxP��K}EX�� �0g0�I01��p�
$TF�a��C$MD3��T�O�3�0U� �� K�Hw2�C1|�	EΡg0wE{vF�vF�40CPp@�a2 m
P$A`PU�3N)#�dR*��AX�!sDETAI�3BUFV��p@1� |�p۶�pPIZdT� PP[�MZ��Mg�Ͱj�F[�SIMQSI�"0��A.�p�����lw Tp�|zM��P�B�FAkCTrbHPEW7�`P1Ӡ��v��MCd�� �$*1JB8�p<�*1DECHښ��H��(�c� � �+PNS_EMP���$GP���,P_���3�p�@Pܤ��TC��|r��0�s��b��0�� �B���!
���J�R� ��SEGFRR��Iv �aR�Tkp9N&S,�PVF���>� &k�Bv �u�cu��aE�� !2��p+�MQ��E�SIZ�3����T��P�����>�aRSINF��� ��kq���������LX�����F�CRCMu�3CClpG��p� ��O}���b�1��������2�V�DxIC��C ���r����P��{� SEV �zF_�եF�pNB0�?�p�����A�! �r �Rx����V�lp�2ݠ�aR�t�,�g�qR>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!��$SK��2&p�DB�"�"@�;PR8� 
� ����# >�q1M$��$��+�L9!$?(�V�%@?R4�C&_?R4ENE���'~?(�� R�E�pY2(H v�OS��#$L�3$$3R��;3�MV�Ok_D@!V�RO�Scrr�w�S���CR�IGGER2FPA��S��7�ETURN�0B�cMR_��TUrː[��0EWM%���GN>`��RL�A���Eݡ�P�'&$P�t�'�@4a"��C�DϣV�DXQ���4�1��MVGO_A7WAYRMO#�a�w!� CS_)7  `IS#�  �� �s3S�AQ汯 4Rx�ZSW�AQ�p�@r1UW��cTNTV)�5RV
a���|c�éW�ƃ��JB��x0��S�AFEۥ�V_SV>�bEXCLUU�;���ONL��cY�g�~az�OT�a{�HI_V? ��R, M��_ *�0� ��_�z�2� 	CdSGO  +�rƐm@��A�c~b���w@��V��i�b�fANNUNXx0�$�dIDY�UABc�@Sp�i�a+ �jP�f��ΰAPIx2,���$F�b�$ѐOT��@A $DUMMY��Ft��Ft±�� 6U- ` !�HE�|s��~b�c�B@ SUFFI���4PCA��Gs5Cw6Cq�!M�SWU. 8!�KgEYI��5�TM�10�s�qoA�vINޱ��D, / D��H7OST�P!4����<���<�°<��p<�E�M'���Z�� SBL�� UL��0  ��	����DT��01 � $|��9USAMPL�@��/���決�$ I@|갯 $SUBӄ���w0QS�����#��SAV�����c�S< X9�`�fP$�0E!�� YN_B�#2 M0�`DI�d�pO|��m��#$F�R_I�C� �ENC2s_Sd3  ��< 3�9���� cgp����4�"��2�A9��ޖ5���`ǻ�@Q@K&D-!�a�AVER�q��λ�DSP
���PC�_�q��"�|�ܣ�V7ALU3�HE�(��M�IP)���OP5Pm �TH�*�D�S" T�/�Fb�;�d����d D��q�1�6 H(rLL_DUǀ�a�@��k����֠OT�"U�/���P�R_NO�AUTO70�!$}�x�~�@s��|��C� ��C� 2�iaz�L�� 8H *��L� ��� Բ@sv��`� �� ÿ� ��Xq��cq���q���q���7��8��9��0T���1�1 �1-�U1:�1G�1T�1aʕ1n�2|�2��2� �2-�2:�2G�2�T�2a�2n�3|�3R�3� �3-�3:�U3G�3T�3a�3nʅ4|������9� <���z�ΓKI`����H硵BaFEq@�{@: ,��&a?g P_P?��>�����E�@��v��QQ��;fp$T�P�$VARI�����,�UP2Q`< W�߃TD��g�����`������%���BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P�"r�l@``>�t ;��6����ST����T��M ����0	��i��� F���������kRt �����FORCEUP��b܂FLUS
pH�(N��� ��6bD_CM�@E�7N� p(�v�P��REM� Fa��@j��ʥ
K�	N���EF1F/���@IN�QsOV��OVA�	�TROV DT<)��DTMX:e  �P:/��Pq�v,XpCLN _�p���@ ��	_|��_T�: �|�&PA�QDI���1��L0�Y0RQm�_+qdH���M���CL�d�#�RIV{�ϓN"E�AR/�IO�PC�P��BR��CM؍@N 1b 3GC3LF��!DY�(�l�a�#5T�DG����� �%�'�FSS� )�?��)p1�1�`_1"81�1�EC13D;5�D6�GRA���@������PW�ON<2EBUG�S�2���gϐ_E �A ��?����T�ERM�5B�5����ORIw�0C�9S#M_-`���0D�5p���TA�9E�5$Z� �UP��F�3 -QϒA�P�3>�@B$SEGGJ� �EL�UUSEPNFI��pBx��1@�<�4>DC$UF�P���$���Q�@C����G�0T�����SN;STj�PATۡg���APTHJ�A�E *�Z%qB\`F�{E��F��q�pARxPY�aSH�FT͢qA�AX_SGHOR$�>��6 @�$GqPE���OV�R���aZPI@P@$Uz?r *aAYLO���j�I�"��Aؠ��ؠERV��Qi�[Y )��G�@R��i�e���i�R�!P�uASY1M���uqAWJ�G)��E��Q7i�RD�U�[d�@i�U��C�%UP����P���WOR�@Mv��k0SMT���G��GR��3�aP�A�@��5�'�H ׸ j�A�TO�CjA7pP]Pp$OPd�O��C�%�pe�O!��RE.p�R�C�AO�?��Be5pR�EruIx'QG��e$PWR) IMdu�RR_$s��5��B� Iz2H8�=�_�ADDRH�H_LENG�B�q�q:�x��R��So�J.�SS��SK������ Ì�-�SE*���rS�N�MN1K	�`j�5�@r�֣OL���\�WpW�Q�>pACRO�p���@H ����Q8� ��OUPW3�bE_>�I��!q�a1�� ������|���������-���:���iIOX2S=�D�e��<]���L $��p��!_OFF[r_�P�RM_��aT�TP_�H��M (�pOBJ�"�pG�[$H�LE�C��>ٰN � 9�*��AB_�T��
�S��`�S��LV��KR�W"duHITCOU�?BGi�LO�q ����d� Fpk�GpsSS� ���HWh��wA��O.��`IN�CPUX2VISIO��!��¢.�á<��á-� �IOLN.)�P 87�R'�[p�$SL�bd P7UT_��$dp��Pz �� F_AuS2Q/�$LD���D�aQT U�0]P�Aa������PHYG�d��Z�Ͱ5�UO� 3R `F���H�Y q�Yx�ɱvpP�Sdp����x��ٶBP�UeJ��S����NE�W�JOG�G �DIS���&�KĠ��3T �|��AV��`_�CTyR!S^�FLAGf2v&�LG�dU �n��:��3LG_SIZ��ň��=���FD��I����Z �� ���0�Ʋ�@s��-ֈ� -�=�-���-��0-�I�SCH_��Dq��NT?���V��EE!2�C��n�U�����`�L�Ӕ�DAU��E�A��Ġt����GH�r��I�BOO)�W�L ?`�� ITpV���0\�REC�GSCRf 0�a�D^�<����MARG��`!�P�)�T�/ty�?I�S��H�WW�I���T�J{GM��MNCH��I�FNKEY��Kn��PRG��UF��܋P��FWD��HL.�STP��V��@X�����RSS�H�` �Q�C�T1�ZbT�R ���U�����|R���t�i���G��8PPO���6�F�1�M��FO{CU��RGEXP��TUI��IЈ� c��n��n����eP@f���!p6�eP7�N����CANAI�jB��V7AIL��CLt!;e?DCS_HI�4�D.��O�|!�S �Sn���_�BUFF1XY��PT�$�� �vD��f�LL6q1YY���P �����pOS�1�2�3���_|�0Z �  ��aiE�*��IDX�dP�RhrO�+��AV&ST��R��Yz�~<! Y$EK&CK+���Z&m&KF�1[ L��o�0�� ]PL�6pwq�t^����w���7�_ \ ��`��瀰�7��#�0C��] ��CLD�P��;eTRQLI��jd.�094FLG z�0r1R3�DM�R7Ɩ�LDR5<4R5ORG.���e2(`���V�8�.��T<�4�d^ ��q�<4��-4R5S�`T�00m��0DFRCLMC!D�?�?3I@���MIC��d_ d����RQm�q�DgSTB	�  �Flg�HAX;b �H>�LEXCESZr�RrBMup�a`� �B�;d��rB`��`a��F_A�J��$[�O�H:0K�db \��ӂnS�$MB��LIБ~}SREQUIR�R�>q�\Á�XDEBUT��oAL� MP�c�b�a��P؃ӂ!BKMND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@qt��o��UPST8�w e�rLOC��RI�p�EX�fA��p��AoAODAQnP�f X��ON��[rMF�����f)�"�I��%�e��T���FX�@IGG� g �q��"E�0��#���$R�a%;#7y���Gx��VvCPi�DAT	Aw�pE:�y��RF����NVh t W$MD�qIё)�v+�tń�tH�`�P�ux�|��sANSW}�P�t�?�uD�)�b��	@Ði �@C�U��V�T0�eRR2�j Dɐ�Qނ~�Bd$CALI�@�F�G�s�2�RI�N��v�<��NTE���kE���,��b����_Nl��ڂ���kDׄRm�DIVFiFDH�@ـn��$V��'c!$��$Z������~�[��oH ?�$BELTb��!_ACCEL+��ҡ��IRC�t���T/!��$PS �@#2��Ė83����x��� ��PATH���������3̒Vp�A_@�Q�.�4�B�C�_MGh�$D�DQ���G�$FW�h��p��m�����b�D}E��PPABNԗROTSPEED����00J�Я8��@����$USE_d��P��s�SY���c�A kqYNu@A�g��OFF�q�M�OUN�NGg�K�O9L�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I̒��4��\BݠVEO�w�Ͳ2�3_UPE�߳LOWL���00����D���BwP��� ��1RCʀƶMOSI�V�JRMO���@GP�ERCH  �OV��^��i�<!� ZD<!�c��d@�P��BV1�#P͑��L�0��EW��ĸUP��Ŝ���TRKr�"AYLOA'a�� Q-��(�<�1Ӣ`0 ��RT1I$Qx�0 MO���Ѐ�B R�0J��D��s��H����b�DUM2�(�S_BCKLSH_C(���>�=�q� #�U��ԑ���2�t�]ACLALvŲ�1nМP�CHK00'%SD�RTY4�k��y�1�q_6#2�_UM�$Pj�Cw�_�SCL���ƠLMT_J1_LO��@���q��E�����๕�幘SPC��7������PCo���H� �PU�2m�C/@�"XT_�c�CN_��N��e���SFu���V�&#�� ��9�(���=�C�u�SH6#��c����1�р��o�0�͑
��_�P�At�h�_Ps�W�_ 10��4�R�01D�VG��J� L�@J�OG|W���TORQU��ON*�Mٙ�sRH�L���_W��-�_=���C��I��I�IJ�II�F�`�JLAX.�1[�VC��0�D�BO1U�@i�B\�JRKU��	@D�BL_SMd�BM�%`_DLC�BGR�V��C��I��H�_� �*COS+\�(LN�7+X >$C�9)I�9)u*c,�)�Z2 HƺMY�@!�( "TH&-�)T�HET0�NK2a3I��"=�A CB6CB=�C�A�B(2061C�616SBC�T2N5GTS QơC� �aS$" �4c#�7r#$DUD�EX�1s� t��B�6���AQ|r�f'$NE�DpIB U�H\B5��$!��!A�%�E(G%(!LPH$U�2׵�2SXpCc% pCr%�2�&�C�J�&!�EVAHV6H3�YLVhJUVuKV�KV�KV�KV�KV�IHAHZF`RPXM��wXuKH�KH�KUH�KH�KH�IO2L�OAHO�YWNOhJO�uKO�KO�KO�KO
�KO�&F�2#1ic%��d4GSPBALA�NCE_�!�cLE6k0H_�%SP��T&��bc&�br&PFUL�C�hr�grr%Ċ1=ky�UTO_?�j�T1T2Cy��2N &�v�ϰctw�g�p�0(Ӓ~���T��O���>� INSEGv�!��REV�v!���DI�F��1l�w�1m
�OB�q
�����MIϰ1��LCHgWAR����AB&~u�$MECH,1�� :�@�U�AX:�P���Y�G$�8pn 
pZ��|���ROBR��CR(���N�'��MSK_�`f�p� P Np_��R ����΄ݡ�1��Ұ�Т΀ϳ��΀"�IN��q�MTCOM�_C@j�q  �L��p��$NO�RE³5���$�7r 8� GR�E��SD�0ABF�$?XYZ_DA5A���DEBU�qI���Q�s �`$�COD�� ��k�F��f�$BUFIwNDXР  ���MOR��t $-�U��)��r�B����͓�Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��Ex����OPWO��ŀv0��SYS�BU�@ʐ$SOP�����#�U"��pPgRUN�I�PA��DH�D����_OUb�=��qn�$}�/IMAG��ˀ�0�P�qIM����IN��q���RGOVR!Dȡ:���|�P~���Р�0L_6p���i⦄�RB���0��ML���EDѐF� ��%N`M*������˱�SL�`ŀw x �$OVSL�vS;DI��DEXm�g� e�9w�����V� ~�N���w����Ûǖ���M�H͐�q<�>�� x HˁE�^F�ATUS����C�0àǒ��BTMT����If���4����(�ŀy DˀEz�g���PE�r����8�
���EXE��V���E�Y�$Ժ ŀz �@ˁ��UP{�h�$�p��XN���9x�H� �PG"��{ h $SUB��c�@_��01\�_MPWAI��P��&��LO��<�F�p��$RCVFAI�L_C�f�BWD�"�F���DEFSP>up | Lˀ`��D�� U�UNI��S���R`����_L�pP���P�ā}��� B�~����|��`ҲN�`KET���y���P� $�~z���0SIZE] �ଠ{���S<�OR~��FORMAT/p` � F���rEMR��y�UX������PLI7�ā � $�P_SW�I�����_PL~7�AL_ �ސJR�A��B�(0C���Df�$Eh��ւ�C_=�U� � � ���~��J3�0����TIA�4��5��6��MOM������ �B�AD��*��*6 PU70NRW���W R����?� A$PI�6�� �	��)�4l��}69��Q���c�SPEED�PGq�7� D�>D����>t�Mt[��SAM��`痰>��MOV���$��p�5��5$�D�1�$2�� �����{�Hip�IN?,{�F(b+=$��H*�(_$�+�+GA�MM�f�1{�$G#ET��ĐH�D����=
^pLIBR�ѝ]I��$HI��_��HȐ*B6E��*8A$>G086LW=e6\<G9@�686��R��ٰV���$PDCK��Q�H�_���� ;"��z�.%�7�4*��9� �$I/M_SRO�D�s"����H�"�LE�O�0\H��6@�@�U� ��ŀ�P�qUR_�SCR�ӚAZ��S_SAVE_D�,�E��NO��CgA�� ���@�$����I��	 �I� %Z[� ��RX " ��m���"�q�' "�8�Hӱt�W �UpS��ћ�L;@���O㵐.'}q��Cg@���@ʣ����S�M�A�Â� � $P9Y��$WH`'�NGp���H`��Fb��0Fb��Fb��PLM����	� 0h�H�{�X��O���z�Z�eT�M����# pS��C��O@__0_B_�a��_%�� |S����@	�v ��v �@���w�v��9EM��% FR�frJ�B�ː��ftP��PM��QU� ��U�Q��Af�Q�TH=�HOL��Q7HYS�ES�,��UE��B��O#��  ��P0�|�gAQ�(��ʠu���O��ŀ��ɂv�-�A;ӝR#OG��a2D�E��Âv�_�ĀZ�INF�O&��+����b�v�AOI킍 ((@SLEQ/�#� �����o���S`c0QO�0�01EZ0sNUe�_�AUT�Ab�COPY��Ѓ�{��@M��N�����1h�P�
� ��RGI������X_�Pl��$�����`�W��P���j@�G���EX_T_CYCtb����p����h�_N�A�!$�\�<�R�O�`]�� � 9m��POR�ㅣ\���SRVt�)��6��DI �T_l����Ѥ{�ۧ��ۧ �ۧ5*٩6٩7٩8���AiS�B쐒��$�)F6���PL�A�A^�TAR��@E `��Z�����<��d� �,(@FLq`h��@Y�NL���M�C���GPWRЍ�쐔e�ODELAѰ�Y�p�AD#qX� �QSwKIP�� ĕ�Zx�O�`NT!� ��P_x���ǚ@�b �p1�1�1Ǹ�?�  �?��>��>�&�>��3�>�9�J2R�;쐖 4��EX� TQ����ށ�Q����[�KFд���RD�CIf� �U`�X}�R�#%M!*�0�)�~�$RGEAR_0sIO�TJBFLG�L�igpERa��TC݃�������2TH2N���� 1� ��Gq T�0 I����M���`Ib�\��qREF�1�� l�h��ENA9B��lcTPE?@�� ��!(ᭀ����Q�#��~�+2 H�W���2�Қ���"�4�F�X�W P��3�қ{�@��������j�4�����
��.�@�R�j�5�ҝu�����������j�6�Ҟ��P(:Lj�7�ҟo@�����j�8�����"4Fj��SMSK�� � �+@��E�A�QR�EMOTE�������@ "1��Q�I�O�5"%I��P��Rrd�Wi@쐣  �@����X�gpi�쐤���Y"$DSB_SICGN4A�Qi�̰C�о�tRS232%��Sb�iDEVICE�US#�R�RPAR�IT�!OPBI�T�Q��OWCONTR��Q�ѓ�R�CU� M�SUXTASK�3NB��0�$oTATU�P�IS@@쐦F�6�_�P�C}�$FREEFROMS]p�ai��GETN@S�UPD2l�ARBA"SP%0��ߧ� !m$USA���az9�L��ERI�0f��pRY$�5~"_�@f�P�1�!N�6WRK��D9��F9ХFRIEND�Q4bUF��&�A@oTOOLHFMY5��$LENGTHw_VT��FIR�p�qC�@�E� IUF�IN�R���RGyI�1�AITI:�bxGX��I�FG2�7�G1a����3�B�GP1RR�DA��O_� o0e�I1RER�đ�3&����TC���AQJV ��G|�.2���F� �1�!d�9Z�8+5K�+5౑E�y�L0�4�XS �0m�LN�T�3�Hz��89��%�4�3G���W�0�W�RdD �Z��Tܳ��K�a3d���$cV 2����1��I1H�02*K2sk3K3Jci �aI�i�a�L��SL���R$Vؠ�BV�EVPk�]V*R��� �,6 Lc���9V2F{/P:Bֵ�PS_�E��$prr�C�ѳ$A0���wPR���v�U�cS�k�� {���2��� 0���VX`�!�tX`A��0P�Ё�
�5�SK!� �-qRH��!0���z�NJ SAX�!h�A�@LlA���A�THIC�1p�������1TFE��|�q>�IF_CH�3�A�I0�����G1@�x������9�Ɇ7_JF҇PR(����RVAT��� �-p��7@����D9O�E��COU(���AXIg��OFF{SE+�TRIG�S K��c���Ѽ�e�[�K��Hk���8�IGMA�o0�A-��ҙ�OR?G_UNEV���� �S�쐮d� �$������GgROU��ݓTO2���!ݓDSP��JO1G'��#	�_P'�2�OR���>P6KE�Pl�IR�0�PML�RQ�AP�Q��E�08q�e���SYSG��"v��PG��BRK*Rd�r�3�-��������ߒ<pAD��ݓJ�B�SOC� N�D?UMMY14�p\@�SV�PDE_OP�3SFSPD_O+VR��ٰCO��&"�OR-��N�0.��Fr�.��OV�S!Fc�2�f��F��!�4�S��RA�"LCH�DL�RECOV(��0�W�@M�յF�RO3��_��0� @�ҹ@VE}RE�$OFS�@3CV� 0BWDG�Ѵ`C��2j�
�TR�!���E_FDO>j�MB_CM��U�B �BL=r0�w�=q�tVfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�<#�8$CA�{�|����8$HBK|1,c��IO��.�:!aPPA"�N�3�^��F���:"�DVC_DB�C��d�w"���D�!��1���ç�3��^��ATIO� �q�0�UC�&CAB�BS�PⳍP��䖁�_0c�SUB'CPUq��S�Pa  aá�}0�Sb��c��r"~ơ$HW_C���� :c��IcA�A-�l_$UNIT��l���ATN�f����CY{CLųNECA���[�FLTR_2_�FI���(��}&��L�P&�����_SCT@SF_��F����G����FS|!�¹�CH�AA/����2��RSD�x"ѡb�r�: ;_T��PRO��OÖ� EM�_��8u�q u�q���DI�0e�RAIL�AC��}RMƐLOԠdC��:anq��wq�����PR��SLQ��pfC�ѷ 	��F�UNCŢ�rRIN�kP+a�0 ��!RA� >R 
Я��ίWAR�BLFQ��A������DA�����L�Dm0�aB9��nqBTIvrbؑ��μPRIAQ1�"AFS�P�!�����`(%b���M�I1UÇDF_j@��y1°L�ME�FA�@HRDiY�4��Pn@RS@Q��0"�MULSE�j@f�b�q �hX��ȑ���$.A[$�1$c1Ó~���� x~��EG�0ݓ�q!AR����09>B�%AXE��ROB���W�A4�_�-֣S�Y���!6��&S�'W�R���-1���ST�R��5�9�E��C 	5B��=QB90`�@6������OT�0�o 	$�ARY�8�w20���	%�F�I��;�$LINQK�H��1�a_63��5�q�2XY�Z"��;�q�3@��1��2�8{0B�{`D��� CFI���6G��
�{�_J���6��3aOP_dO4Y;5�QTBmAd"�BC
�z�DU"�z66CTURN3��vr�E�1�9�ҍGFL�`���~ �@�5<:y7�� 1�?0%K�Mc�68Cb�8vrb�4�ORQ��X �>8�#op������wq�Uf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W�� �Tυ� ;����QH� !`�ҽ��U�Q�WkeK#�kecXER��	BGE	0��S�dAWa Ǣ:D���7!�!AX�rB!{q��1 uy-!y�pz�@ z�@z6Pz\Pz�  z1v�y�y� +y�;y�Ky�[y��ky�{y��y�q�yD7EBU��$�����L�!º2WG`  A!B!�,��SV���� 
w���m���w� ���1���1���A���A ��6Q��\Q���!�m@���2CLAB3B��U�����S � ÐER���� �� $�@� Aؑ!p�PO��Z�q0�w�^�_MRAȑ�/ d  T�Ĵ�ERR��TYz�B�I�V3@�cΑ'TOQ�d:`L� �d�2�]�X�C[! /� p�`T}0i��_V1�r�a'�
4�2-�2<����@Pq�����F�$W���g��V_!�l�$��P����c��q"�	��SFZN_C;FG_!� 4��?� ��|�ų����@�ȲW� ?]���\$� �n���Ѵ��9c�Q���(�FA�He�,�XEDM�(�����!s��Q�g�P{RV HE�LLĥ� 5�6�B_BAS!�R�SR��ԣo �#S���[��1r�%��2�ݺ3ݺ4ݺ5ݺ6�ݺ7ݺ8ݷ��ROaOI䰝0�0NLK!ưCAB� ��AC-K��IN��T:�1��@�@ z�m�_PUf!�CO� ��OU��P� Ҧ) ��޶���TPFWD_KA1Rӑ��RE~��qP��(��QUE������P
��CSTOPI_AL�����0�&���㰑�0SEM�l�b�|�M��d�TYf|�SOK�}�DI������(���_TM>\�MANRQ�ֿ0�E+�|�$KEY?SWITCH&	����HE
�BEAiT����E� LEҒ���U��FO�����O_HOM�On�REF�PPRzP��!&0��C+�OA��ECO��B�r�IOCM�D8׵��]���8�` � DH�1����U��&�MHx�»P�CFORC��f� ���OM�  � @V��|�U,3P� 1-�`� �3-�4�p �SN�PX_ASǢ� �0ȰADD�����$SIZ��$VsARݷ TIP]�)\�2�A򻡐� ��]�_� �"S꣩!yCΐ��FRIF��S�"�c���NFp��V ��` � x�`SI�TES�R6S�SGL(T�2P&���AU�� ) STM�TQZPm 6BW<�P*SHOWb���SV�\$��; ���A00P�a �6�@�J�T�5�	6�	7�	8
�	9�	A�	� �!� �'��0�F�0 u�	f0u�	�0u�	@�@u[Pu%12U1?1L1Y1fU1s2�	2�	2�	U2�	2�	2�	2�	U222%22U2?2L2Y2fU2s3P)3�	3�	U3�	3�	3�	3�	U333%32U3?3L3Y3fU3s4P)4�	4�	U4�	4�	4�	4�	U444%42U4?4L4Y4fU4s5P)5�	5�	U5�	5�	5�	5�	U555%52U5?5L5Y5fU5s6P)6�	6�	U6�	6�	6�	6�	U666%62U6?6L6Y6fU6s7P)7�	7�	U7�	7�	7�	7�	U777%72U7?7,i7Y7Fim7s�'��VP��UPD��  ���|�԰
��YS�LOǢ� �  z��и���o�E��`>�8^t��АALUץ�����CU���wFOqIgD_L�ӿuHI�z�I�$FILE_���t��$`�^�Ms;SA��� h���?E_BLCK�#�|C,�D_CPU<� {�<�o����t��޴�R ��
P�W O� ��LA���S��������RUNF�Ɂ��Ɂ����F��ꁡ�ꁬ��TB�Cu�C� �Xw -$�LENi� �v������I��G�LOW_AXI�SF1��t2X�M��д�D�
 ��I�� ��}�TOR����Dh��� L=��⇒p�s���#�_MA`�p��ޕ��ޑTCV����T���&��ݡ ����J�����J�����Mo���J�Ǜ �������2�Ѓ v�ة���F�JK��VK�i�Ρv�Ρ3��J0l�ңJJڣJJ�AALң�ڣ��e4�5z�&�N1-�P9���␅�L~�_V�j�;������ =` �GROU�pD���B�NFLIC���REQUIREa�EBUA��p����2¯������c�� \��A�PPR��C���
v�EN�CLOe��S_M v�,ɣ�y
���� ����MC�&���g�_M	G�q�C� �{�9����|�BRKz�NO�L��|ĉ R��_L!I|��Ǫ�k�J����P
���ڣ�����&����/���6��6��8�������� ��8�%�W�2�e�PATHa�z�p�z��=�vӥ�ϰ�x�CN�=�CA�����p�I�N�UC��bq��CO�UM��YZ������qE%���2������PAYLOA��J{2L3pR_AN��<�L��F�B�6�R�{��R_F2LSHR��|�LOG��р���|����ACRL_u� ������.���H�p��$H{���FLE�X
�s�J�� :�/����6��2�����;�M�_�F1 6����n���������ȟ��Eҟ����� ,�>�P�b���d�{� �����������5�	T��X��v��� EťmFѯ���� ���&�/�A�S�e��D�Jx�� � `������j�4pAT��l��n�EL  �%jøJ���ʰJE��gCTR�Ѭ�TN���F&��HAND_�VB[
�pK�� $F2{�6� �rSWm�U���O $$Mt�h�R�À08��@<b 35��^6A@�p3�k��q{9t�A���p��A��A�ˆ0��TU���D��D��P��G��IST��$A��$AN��DYˀ�{� g4�5D���v�6�v��@5缧�^�@��P�� ���#�,�5�>�+p�K�� &0�_��ER!V9�SQASYM$��] �����x�������_SHl����� ��sT�(����(�:�JA���S�cir��_VI�#Oh9�``V_UNI��td�~�J���b�E�b��d ��d�f��n�������H��uN���xQ2�H������"Cq3EN� a�DI��>��ObtC�Dpx�� ��2IxQA����q ��-��s �� s������ ��OMMEB��rr/�TVpPT�P ���qe�i�A���P�x ��yT�P�j� $DUM�MY9�$PSm_��RFq�  ��:� s���!~q�� X����K�ST�s�ʰSBR��M�21_Vt�8$S/V_ERt�O��z����CLRx�A  O�r?p? Oր �� D $GLOB���#LO��Յ�$�o��P�!SYS�ADR�!?p�pT�CHM0 � ,x����W_NA��c/�e�$%SR�?�l (:] 8:m�K6�^2m�i7m� w9m��9���ǳ��ǳ� ��ŕߝ�9ŕ��� i�L���m��_�_�_|�TD�XSCRE�jƀ�� ��STF�Ƶ�}�pТ6�7�D�] _v AŁ� 9T����TYP�r�@K��u�!u���-O�@IS�!��tvC�UE{t� �����H�S���!RSM�_�XuUNEXCcEPWv��CpS_�� {ᦵ�ӕ���÷����COU ��� [1�O�UET�փr|���PROGM� {FLn!$CU��cPO*q��c�I_�p}H;� � 8��.N�_HE
p��Q�~�pRY ?����,�J�*��;�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� D�C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!$��VSHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3��H���w�2u�sqV�rzu��%�DJU��~|#�WAIT�������%ONE���YBOư ?�� $@p%�vC�SBn)TPE��NEC��x"�$t$��.�*B_T��R��% �qR� ���sB�%�tM�+��t�.�F�R!�݀��OPm�MAS��_DOG�OaT	�D����C3S�	�O2DELAY���e2JO��n8E��Ss4'#�J�aP6%�����Y_��O2$��2���5���`? sqZA�BCS��  �$�2��J�
���$�$CLAS�����AB�sp'@@�VIRT��O.@A�BS�$�1 <E�� < *AtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v���8��M@[�AXLրK��*B�dC  ���IqN��ā��PRE������LAR�MRECOV �<I䂥�NG�� �\K	 A  � J�\�M@PPLIMC�?<E�E��Handl�ingTool ��� 
V7.5�0P/28[�  o��c��
�w_SW�� UP*A7� ��F0ڑ���AG@�� S20��*A���:�ާ��oFB �7DA5�� ��'@�cy@��None������� ��T�'*A4�b+xl�_��V����:g�UTOB���������HGAPO�N8@��LA��U��D� 1<EfA����������� Q 1שI Ԁ��Ԑ�:�i�n��܍�#BGB �3��\�HE�Z��r�HTTHKY ��$BI�[�m����� 	�c�-�?�Q�o�uχ� �ϫϽ��������_� )�;�M�k�q߃ߕߧ� ���������[�%�7� I�g�m������� ������W�!�3�E�c� i�{������������� ��S/A_ew �������O +=[as�� �����K//'/ 9/W/]/o/�/�/�/�/ �/�/�/G??#?5?S? Y?k?}?�?�?�?�?�? �?COOO1OOOUOgO yO�O�O�O�O�O�O?_�	__-_K_Q_��(�T�O4�s���DO_C�LEAN��e��SN�M  9� ��9oKo]ooo�o�D?SPDRYR�_%�HI��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ|��g�PLUGGҠ��Wߣ��PRC�`B�`9��o�=�OxB��oe�SEGF��K������o%o�����#�5�m���LAP �oݎ����������џ �����+�=�O�a�>��TOTAL�.����USENUʀ�׫ �X���R(�RG�_STRING �1��
��M��Sc�
��_�ITEM1 �  nc��.�@�R�d�v� ��������п������*�<�N�`�r��I/O SIGN�AL��Try�out Mode��Inp��Simulated��Out��O�VERR�` = �100�In �cycl���P�rog Abor������Stat�us�	Hear�tbeat��M?H FaulB�K�AlerUم�s߅� �ߩ߻��������� �S���Q�� f�x���������� ����,�>�P�b�t�p������,�WOR�� ����V��
.@ Rdv����� ��*<N`PO��6ц��o �����//'/ 9/K/]/o/�/�/�/�/��/�/�/�/�DEV �*0�?Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�OPALTB��A�� �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_�oo(o:o�OGRI �p��ra�OLo�o�o�o �o�o�o*<N `r������`o��RB���o�>� P�b�t���������Ώ �����(�:�L�^�xp����PREG�N ��.��������*� <�N�`�r����������̯ޯ���&�����$ARG_��D �?	���i���  w	$��	[}��]}���Ǟ�\�SB�N_CONFIG� i��������CII_SAV/E  ��۱Ҳ�\�TCELLSE�TUP i�%�HOME_IO��͈�%MOV_8�2�8�REP����V�UTOBACK�
�ƽF�RA:\�� X�Ϩ���'` ���x������ �� ��$�6�c�Z�lߙ���������������� �!凞��M�_�q�� ���2��������� %�7���[�m������ ��@�������!3E$���Jo��p�����INI�@���ε��MESSAG����q�>�ODE_D$��ĳ�O,0.��PA�US�!�i� ((Ol���� ���� /�// $/Z/H/~/l/�/�'a~kTSK  qx�����UPDT%��d0;WSM�_CF°i��еU�'1GRP 2�h�93 |�B��A|�/S�XSCRD+1;1
1; ����/�?�?�? OO$O ��߳?lO~O�O�O�O �O1O�OUO_ _2_D_�V_h_�O	_X���GR�OUN0O�SUP�_NAL�h�	ܢĠV_ED� 1�1;
 �%-B?CKEDT-�_`�!oEo$���a�o�����ߨ���e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[8�5GED4�n�#�� ~�j���ED5Z��Ǐ6� ~��8�}���ED6�����k�ڏ ~G���!�3�ED7��Z��~� ~�8V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W�Ư�
}3�����CR o�����3�տ@ϯ�����P�PNO_DE�L�_�RGE_UN�USE�_�TLAL_OUT q��c�QWD_ABO�R� �΢Q��ITR�_RTN����N'ONSe����CAM_PARA�M 1�U3
 �8
SONY �XC-56 234567890�H� � @����?���( Щ�V�|[r؀~�X�HR5k�|U�Q��ο�R57����A�ff��KOWA SC310M|[�r�̀�d @6�|V��_�Xϸ� ��V��� ���$�6���Z�l��CE_RIWA_I857ЍF�1��R|].��_LIO4W=� ���P<~�F<�GwP 1�,����_GYk*C*�  ��C1� 9J� @� G� �CL�C]� d� l� s��R� ��[�m�� v� � �� ��� C�� �"��|W��7�HEӰON�FI� ��<G_P_RI 1�+P� m®/���������'CHKPAU�S�  1E� ,�>/P/:/t/^/�/ �/�/�/�/�/�/?(?@?L?6?\?�?"O������H�1_MO5R�� �0�5 	 �9 O�?$O@OHO6K�2	���=$9"�Q?55��C�P)K�D3P������a�-4�O__|Z
�OG_�7�PO��� ��6_��,xV�AD�B���='�)
m�c:cpmidb�g�_`��S:�(�����Yp�_)o�S`	�BBi�P�_mo8j�(�Koo�o9i+�(��og�o�o
�m�of�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`(ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCo��C|��Cq�D��C����C�{iSZE@D���F.��F���E⚵F?,E�ٙ�E@�F�N�IU���I?O�I<#�I6�I洤SY���vqG��T�Em�(�.��(��(��<�q�G�x�2��Ң �� a�D��j���E�e��EX��EQ�EJ�P F�E�F�� G�ǎ^�F E�� FB�� H,- Ge���H3Y����  >�33 s���xV  n2xQ@��5Y��8B� yA�AST<#�
�� �_'�%��wRS/MOFS���~2��yT1�0DE ��O c
�(�;��"�  <�6�z�Rb���?�j�C4�)�SZm� W��{�Jm�C��B-G�C�`�@$�q��T{�FPROG %i����c�I��� �Ɯ��f�KEY_TBL�  �vM�u� �	�
�� !�"#$%&'()�*+,-./01�c�:;<=>?@�ABC�pGHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������p���͓���������������������������������耇���������������������9�!j�LCK��.�<j���STAT����_AUTO_DO���W/�INDTO_ENB߿2R���9�+�T2w�XSTsOP\߿2TRLl��LETE����_�SCREEN �ikcsc���U��MMENU� 1 i  <g\��L�SU+�U� ��p3g�������� ����2�	��A�z�Q� c��������������� .d;M�q ������ N%7]�m� ��/��/J/!/ 3/�/W/i/�/�/�/�/ �/�/�/4???j?A? S?y?�?�?�?�?�?�? O�?O-OfO=OOO�O sO�O�O�O�O�O_�O�_P_Sy�_MAN�UAL��n�DBC�OU�RIG���DOBNUM�p��<����
�QPXWOR/K 1!R�ү�_�oO.o@oRk�Q_A�WAY�S��GC�P ��=��df_A!L�P�db�RY����t���X_�p 1"�� , 
�^��P�o xvf`MT�I^��rl@�:sONTImM������Zv�i
õ�cMOTN�END���dREC�ORD 1(R�8a��ua�O��q� �sb�.�@�R��xZ� ������ɏۏ폄� ��#���G���k�}��� ��<�ş4��X��� 1�C���g�֟������ ��ӯ�T�	�x�-��� Q�c�u���������� >����)Ϙ�Mϼ� F�࿕ϧϹ���:��� ����%�s`Pn&�]�o� �ϓ�~ߌ���8�J��� ��5� ��k����� ���J�����X��|� ��C�U�����������0�����	��dbTOLERENCqdsBȺb`L�͐P�CS_CFG �)�k)wdMC�:\O L%04dO.CSV
�Pc��)sA �CH� z�P)~���hM�RC_OUT �*�[�`+P SG�N +�e�r���#�10-MAY�-20 10:3�3*V17-FEB�j9:09�k PQ�8��)~��`pa�m�?�PJPѬ�VERSION �SV2.�0.8.|EFLO�GIC 1,�[ 	DX�P7)�P�F."PROG_E�NB�o�rj ULS�ew �T�"_WRSTJNEp�V�r`d�EMO_OPT_�SL ?	�es
� 	R575 )s7)�/??*?<?'>�$TO  �-�l�?&V_@pEX�W�d�u�3PATHw ASA\�?��?O/{ICT�aF�o`-�gds�egM%&AST?BF_TTS�x�Y�^C��SqqF�PM�AU� t/XrMSWR.�i6.|S/�Z!D_N�O0__�T_C_x_g_�_�tSB�L_FAUL"0��[3wTDIAU 1�6M6p�A�12345678#90gFP?Bo Tofoxo�o�o�o�o�o �o�o,>Pb��S�pP�_ �� �_s�� 0`��� ��)�;�M�_�q��� ������ˏݏ��|)gUMP�!� �^��TR�B�#+�=�P�MEfEI�Y_TE{MP9 È�3@8�3A v�UNI�.(�YN_BRK �2Y)EMGDI�_STA�%WЕN�C2_SCR 3��1o"�4�F�X� fv���������#��ޑ14����)��;�����ݤ5�����x�f	u�ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/߭P�b�t��  ��xߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N���r������� ��������&8 J\n����� ���"`�FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/4 ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O?�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�O�O�o�o�o 
.@Rdv� �������� *�<�N�`�r����o�� ��̏ޏ����&�8� J�\�n���������ȟ�ڟ����H�ETM�ODE 16��]� ��ƨ�
R�d�v�נRRO�R_PROG �%A�%�:߽�  ���TABLE  A������#�L��RRSEV_NU�M  ��Q���K�S���_AU�TO_ENB  q��I�Ϥ_NOh�� 7A�{�R��  *������������^�+��Ŀֿ迄�HISO�͡I��}�_ALM 18.A� �;�����+�e�wωϛϭ����_H���  �A���|��4�TC�P_VER !�A�!����$EXTLOG_REQ�s�{�V�SIZ_�~Q�TOL  ͡{Dz��A Q�_BWD����r����n�_DI�� 9��}�z�͡m���STEP����4��_OP_DO����ѠFACTORY�_TUN�dG�E�ATURE :�����l�H�andlingT�ool ��  -� CEngl�ish Dict�ionary��O�RDEAA �Vis�� Mas�ter���96 �H��nalog �I/O���H55�1��uto So�ftware Update  ���J��matic �Backup��P�art&�gr�ound Edi�t��  8\ap�Cameraz��F��t\j6R��ell���LOA�DR�omm��sh�q��TI" ��cyo��
! o����pane�� �
!��tyle select��H59��nD���o�nitor��48�����tr��Rel�iab���adi�nDiagn�os"����2�2 u�al Check� Safety �UIF lg\a���hanced �Rob Serv> q ct\��lUser FrU���DIF��Ext�. DIO ��f�iA d��en]dr Err L@���IF�r��  �П�90��FCT�N MenuZ v�'��74� TP �In��fac � SU (G�=�p��k Exc�n g�3��Hig�h-Sper Sk]i+�  sO�H9 ~� mmunic!��onsg�teurh� ����V����^conn��2��{EN��Incr�stru���5.�fdKARE�L Cmd. L�?uaA� O�R�un-Ti� EnIv����K� ��+%��s#�S/W��74���License|T�  (Au* �ogBook(S�y��m)��"
�MACROs�,V/Offse6��ap��MH� �����pfa5�Mec�hStop Pr3ot��� d�b =i�Shif���/j545�!xr ��#��,�qb o�de Switc]h��m\e�!oz4.�& pro��4��g��Mul�ti-T7G��n�et.Pos Regi��z�}P��t Fun����3 Rz1��Nu!mx �����9m�1>�  Adjuj��O1 J7�7�* ��<���6tatuq1EIKRDMt�ot��scove�� ��@By- }Ouest1�$Go� �� U5\SNPX b"���YA�"Libr����#b�� �$~@h�pd]0��Jts in VCCM�����0�q  �u!��2 R�0��/I�08��T�MILIB�M J�92�@P�Acc�>�F�97�TPT�X�+�BRSQelZ0�M8 Rm��q%��692��Une�xceptr mo�tnT  CVV�P���KC����+�-��~K  II)��VSP CSXC��&.c�� e�"�� =t�@Wew�gAD Q�8bvr �nmen�@�iP�� a0y�0�pfG�ridAplay !� nh�@*�3R�1�M-10iA(B�201 �`2V" y F���scii��load��83 �M��l����Gua=r�d J85�0�maP'�L`���stua�Pat�&]$Cyc8���|0ori_ x%oData'Pqu���ch�1��g`� mj� RLJam�5����IMI De�-B(\A�cP" #�^0C  etk}c^0asswo%q.�)650�ApU��Xnt��Pven��CTqH�5�0�YELLOW BqO?Y��� Arc�0�vis��Ch�W�eldQcial44Izt�Op� ��gs�` 2@�a��p�oG yRjT1� NE�#HT� xyWb��! �p�`!gd`���p\� =P���JPN ARCP�*PR�A�� �OL�pSup̂f�il�p��J�� ��cro�670�1C~E��d��SS�pe�t�ex�$ �P� Soz7 t� ssagN5� <Q�BP:� �9 �"0�QrtQC��P�l0dpn�笔�r�pf�q�e�ppm�ascbin4p�syn�' ptx�]08�HELNC�L VIS PK�GS �Z@MB �&��B J8@I�PE GET_V�AR FI?S (�Uni� LU�OO�L: ADD�@2/9.FD�TCm���E�@DVp���`A��ТNO WTWTOEST �� ��!���c�FOR ��E�CT �a!� AL�SE ALA`�CPMO-130���� b D: HAN?G FROMg���2��R709 D�RAM AVAI�LCHECKS �549��m�VPC�S SU֐LIM�CHK��P�0x�F_F POS� F��� q8-12� CHARS�ER>6�OGRA ��Z@wAVEH�AME��G.SV��Вאn$���9�m "y�TR}Cv� SHADP��UPDAT k�0>��STATI���? MUCH ����TIMQ MOTN-003��@�OBOGUIDE? DAUGH���b8��@$tou� �@�C� �0��PATH|�_�MOVET��� R64��VMX�PACK MAY ASSERTjS޴�CYCL`�TA���BE COR �71�1-�AN��R�C OPTION�S  �`��APSwH-1�`fix��2�SO��B��XO򝡆��_T��	�i��0j���du�byz p cwa��y�٠HI������U�pb XSP�D TB/�F� \�hchΤB0���EmND�CE�06\Q��p{ smay In@�pk��L ���traff#�	� ���~1from �sysvar s�cr�0R� ��d�DJU���H�!A���/��SET ER�R�D�P7����N�DANT SCR�EEN UNRE�A VM �PD�D���PA���R�I�O JNN�0�F�I��B��GROUNנD Y�Т٠��h�SVIP 5�3 QS��DIGI?T VERS��k���NEW�� P0�6�@C�1IMAG��ͱ���8� DIx`���pSSUE�5���EPLAN J=ON� DEL���1�57QאD��CALLI���Q��m����IPND}�IMG� N9 PZ�19޴�MNT/��ES� ���`LocR HCol߀=��2�Pn� �PG:��=�M��c�an����С: �3D mE2vie�w d X��e�a1 �0b�pof �Ǡ"HCɰ�AN�NOT ACCE�SS M cpite$Et.Qs a� {loMdFlex)a�:��w$qmo G
�sA9�-'p~0��h0�pa��eJ AU�TO-�0��!ip�u@Т<ᡠIABL�E+� 7�a FPL�N: L�pl lm� MD<�VI�����WIT HOCv�Jo~1Qui�t�"��N��USB�@��Pt & rem�ov���D�vAxi�s FT_7�PG�ɰCP:�OS-�144 � h s� 268QՐOST��p  CRASH� DU��$P��W�ORD.$�LOgGIN�P��P:	��0�046 iss�ueE�H�: Solow st��c�`6����໰I�F�IMPR��SPOT:Wh4���N1�STY��0VMGqR�b�N�CAT��-4oRRE�� � 58�1��:%�R�TU!Pe -M a�SE:�@pp���AGp�L��m@al�l��*0a�OCB �WA���"3 CN�T0 T9DWro>O0alarm�ˀm0d t�M�"0�2�|� o�Z@OME�<�� ��E%  #1�-�SRE��M�st�}0g     �5KANJI5n�o MNS@�I�NISITALI�Z'� E�f�we���6@� dr�@ f�p "��SCII� L�afails� w��SYSTaE[�i��  � tMq�1QGro8�m n�@vA����&���n�0q��RWR=I OF Lk���� \ref"�
�u�p� de-rel}a�Qd 03.�0�SSchőbet�we4�IND e�x ɰTPa�DOȬ l� �ɰGi�gE�soperawbil`p l,��aHcB��@]�le�Q0cflxz�Ð���OS {����v4pwfigi GLA�$��c2�7H� la�p�0ASB� Ifz��g�2 l\c�0��/�E�� EX'CE 㰁�P���$i�� o0��Gd`]���fq�l lxt��EFal��#0��i�O�Y�n�CLOSn��SRNq1NT^��F�U��FqKP�AN�IO V7/ॠ1p�{����DB �0ء�ᴥ�ED��DE�T|�'� �bF�N�LINEb�BUG�T���C"RLIB���A��ABC J�ARKY@��� r7key�`IL���P�R��N��ITGAR
� D$�R �Er�� *�T��a�U�0��h�[�ZE V� �TASK p.vr�P2" .�XfJ��srn�S谥dIB�P	c���B/��B�US��UNN�  j0-�{��cR'���LOE�DIVS�C�ULs$cb����BW!��R~�W`P���&��IT(঱tʠ�{OF��UNEXڠ�+���p�FtE��S�VEMG3`NML� 505� D*�C?C_SAFE�P*�p �ꐺ� PET��8'P�`�F  !���IR����c i S�>� K��K�H �GUNCHG��S^�MECH��M��T*�%p6u��tP�ORY LEAKr�J���SPEg�D��2V 74\G�RI��Q�g��CTLN��TRe @�_��p ���EN'�IN�������$���r��T�3)�i�STO�A$�s�L��͐X	����q��Y� ��TO2�J m��0F<�K�����DU�S��O��3$ 9�J F�&�����SSVGN-18#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRKC�TR/"� �q\j5���_�Q�S�qINVJ0D ZO�Pݲ�� �s��г�Ui ɰ̒�a��DUAL� J�50e�x�RVO1/17 AW�TH!�Hr%�N�247%�5q2��|�&aol ���R���at�Sd�cU8���P,�LER��i�x�Q0�ؖ  ST����Md�Rǰt� \fosB�A�0Np�cб���{�U��RO�P 2�b�pB��ITP4M��b !�AUt c0< � pl�ete�N@� �z1^qR635 (�AccuCal2zkA���I) "�(ǰ�1a\�Ps��ǐ � bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etaca2��AT���PC�`��슰�_p�.pc�!Ɗ��:�circB���5�tl��Bɵ��:�fm+�Ί�V�b��ɦ�r�upfrma.����ⴊ�xed�8�Ί�~�pedA�D ��}b�ptlib0B�� �_�rt�߄	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̆�D����c�Ӳ�5�j>ʌ����tcȐ��	�r(����mm 1��T�#sl^0��T�mѡ�&#�rm3��ub Y��q�std}��pl�;�&�ckv�=�r�vaf�䊰��9�vi������ul�`�0fp�q� �.f��� d�aq; i Data� Acquisi
��n�
��T`���1�89��22� DMCM RR[S2Z�75��9 ?3 R710�o�59p5\?��T{ "��1 (D�T� nk@���������E Ƒȵ��Ӹ�et3dmm ��ER����gE��1�q\mo?۳�=(G����[(

�2�` ! ��@JMACRO���Skip/Of�fse:�a��V�4�o9� &qR662����s�H�
 6�Bq8����9Z�4_3 J77� 6�J783�o ���n�"v�R5IK�CBq2 PTLC�Zg R�3 (�s, ��������03�	зJԷ\�sfmnmc "MNMC����ҹ�%wmnf�FMC"�Ѻ0ª etmcr�� �8����� ,�qD�q�   874�\prdq>,jxF0���axisH�Process �Axes e�rol^PRA
�Dp� �56 J81j�5-9� 56o6� ��l�0w�690 98� �[!IDV�1��2(8x2��2ont�0�
 ����m2���?C���etis "I�SD��9�� FpraxRAM�P� D��defB�,�G�isbasicH�B�@޲{6�� 70U8�6��(�Acw: ������D
�/,��AMOX�� ��DvE��?�;T��>Pi� RAFM';�]�!PAM�V�W��Ee�U�Q'
bU�7y5�.�ceNe� �nterfaceh^�1' 5&!54�K<��b(Devam±��/�#���/<�Tane`"DNEWE���btpdnui �A�I�_s2�d_rsCono���bAsfj|N��bdv_arFv�f�xhpz�}w��hkH9xstc��gAp�onlGzv{�ff ��r���z�3{�q'Td>pcha�mpr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�!��pcchmp]aM�P&B�� �mpe�v�����pcs���YeS�� MacKro�OD��16Q! )*�:$�2U"_,��Y�(PC ��$_;�������o��J�geg{emQ@GEMSW�|~ZG�gesndy�<�OD�ndda��Sƕ�syT�Kɓ�su^Ҋ���n�m���L��O  ���9:p'�ѳ޲��spotplusp���`-�W�l�J�s��t[�׷p�key�ɰ�$��s��-Ѩ�m���\fea;tu 0FEAWD�oolo�srn '!2 p���a�As3���tT.� (N. A.)��!e!(�J# (j�,��o�BIB�oD -�.�n6��k9�"K��u[�-�_���p� "P�SEqW����wop "sEЅ�&�:� J������y�|��O8� �5��Rɺ���ɰ[� �X�������%�(
 ҭ�q HL�0k� 
�z�a!�B�Q�"(g�Q�����]�'� .�����&���<�!ҝ_�#��tpJ�H�~Z�� j�����y������2 ��e������Z����V� �!%���=�]�͂���^2�@iRV� on��QYq͋JF0� 8�ހ�`�	(^�dQueue���X\1����`�+F1tpvtsen��N&��ftpJ0v �RDV�	f���J1 Q���v�eyn��kvstk���mp��btkcl�rq���get�����r��`k�ack�XZ�st1rŬ�%�stl��~Z�np:!�`�� �q/�ڡ6!l�/Yr$�mc�N+v3�_`� ����.v�/{\jF��� �`�Q�΋ܒ�N50 (�FRA��+��͢f?raparm��Ҁ��} 6�J643�p:V�ELSE
�#�VAR $SG�SYSCFG.$��`_UNITS �2�DG~°@�4Jgfqr��4A�@FRL-� �0ͅ�3ې���L�0 NE�:�=�?@�8�v�9~Qx304��;�B�PRSM~QA�5T�X.$VNUM_�OL��5��DJ50�7��l� Functʂ"qwAP��琉�G3 H�ƞ�kP9jQ��Q5ձ� ��@jLJ zBJ[�6N�kAP�����S��"TPPRp���QA�prna�SV�ZS��AS8Dj5k10U�-�`cr�`8 ��ʇ�DJR`jYȑH  �Qm �PJ6�a21���48AAVM3 5�Q�b0 lB�`�TUP xbJ�545 `b�`61�6���0VCA�M 9�CLI�O b1�5 ����`MSC8�
rP� R`\sSTYL MNIN�`oJ628Q  �`�NREd�;@�`SC�H ��9pDCSU� Mete�`OR�SR Ԃ�a04 �kREIOC ��a5�`542�b9 vpP<�nP�a�`�R�`�7�`�MAS�K Ho�.r7 <�2�`OCO :��r�3��p�b�p���r0�X��a�`13\mn��a39 HRM"��q�q��LCH}K�uOPLG B��a03 �q.�pH�CR Ob�pCpP�osi�`fP6 i=s[rJ554�òp'DSW�bM�D�pqR��a37 }Rjr0 L�1�s4 �R6�7���52�r5 �2�r7� 1� P6���Re�gi�@T�uF�RDM�uSaq%�4�`930�uSNB�A�uSHLB̀\�sf"pM�NPI��SPVC�J5�20��TC�`"M�NрTMIL�I=FV�PAC W�poTPTXp6.%��TELN N M�e�09m3U�ECK�b�`UFR��`��VCOR��V�IPLpq89qSX9C�S�`VVF�J��TP �q��R62]6l�u S�`Gސ~�2IGUI�C���PGSt�\ŀH863�S�q�����q�34sŁ684`���a�@b>�3 :B抂1 T��96 :.�+E�51 y�q353�3�b1 ���b31 n�jr9 ���`�VAT ߲�q75� s�F��`�sAWSyM��`TOP u��ŀR52p���a809 
�ށXY q���s0 ,b�`885�QXрOLp}�"pE�v��tp�`LCMDў�ETSS���6� �V�CPE o�Z1�VRCd3
�NuLH�h��001m2�Ep��3 f��p��4� /165C��6�l���7PR��00�8 tB��9 -2[00�`U0�pF�1&޲1 ��޲2L"����p��޲4��5 �\hmp޲6 RB�CF�`ళ�fs�8� �Ҋ��~�J�7 OrbcfA�L�8\P0C����"�32m0u��n�K�Rٰn�5 5oEW
n�9 zΊ�40 kB��3 ��6ݲ�`00iB%/��6�u��7�u���8 µ������sU0��`�t �1 05\;rb��2 E��K���j���5˰��6A0��a�HУ`:�63�`jAF�_���F�7 ڱ�݀H�8�eHЋ��cUI0��7�p��1u��8u��9 73�������D7� ��5\t�97 ��8U�Q1��2��1�1:����h��1np�"��8�(�U1��\pyl���,࿱v ��B�85E4��1V���D�4��im��1�<���$>br�3pr�4@pGPr�6 B���цp���1����1�`͵15=5ض157 �2�у62�S����1�b��2����1Π"�2L���B6`�1<cf�4 7B�5 DR���8_�B/��18�7 uJ�8 06��90 rBn�1 �(��202 0E�W,ѱ2^��2��9�0�U2�p�2��2 �b��4��2�a"RiB����9\�U2�`xw�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`ڰR,:7 �2��V�2��5���2^��a^9���qr�����n�5����5᥁"�8Ha�Ɂ}�5B���5������`UA���� ��8�6 �6 S�0��5��p�2�#�529 ��2^�b1P�5�~�2`���&P5���8��5��u�!�5\��ٵ544��5��	R�ąP nB^z�c (�4�����SU5J�V�5��1�1@^��%�����5 �b21��gA��5m8W82� rb��95N�E�5890r�: 1�95 �"�� ����c8"a��|�L (���!J"5|6��^!"�6��B�"8�`#���+�8%�6B�AM�E�"1 iC��622�Bu�6V��d� �4��84�`ANR�SP�e/S� �C�5� �6� ��� \@� �6� �V� 3t��?� T20CA�R���8� Hf� 1DH��� AOE� ��w ,�|�� �0X\�� �!64K��ԓ�rA� �1 (M-7�!/50T�[PM��P�Th:1�C�#P�e� �3�0� 5`M�75T"� �D8p�! �0Gc� u�4��i1�-710i�1� S�kd�7j�?6�:-HS,� �RN�@�UB��f�X�=m75sA*A6an���!/CB�B2.6A �0;A�C�IB�A�2�QF1�UB2:�21� /70�S� �4����Aj1�3p����r#0 B2\m*A@C��;bi"i1K��u"A~AAU� imm7c7��ZA@I�@�Df�A�D5*A�E� #0TkdR1�35Q1�" *�@�Q�1�QC)P�1 *A�5*A�EA�5B�4>\77
B7=Q�D�2H�Q$B�E7�C�D/qA	HEE�W7�_|`jz@@� 2�0�Ejc7(�`�E"l7�@7�A
1��E�V~`�W2%Q�R9\ї@0L_�#��� �"A���b��H3s=rA/2�R5nR4�7�4rNUQ1ZU�A�s\m9
1M92L2�!F!t^Y�ps� 2ci��-?�qhimQ�t  w0 43�C�p2�mQ�r�H_ �H20�Evr�QHsXBFSt62�q`s����� ��Pxq350_�*A3I)�2�d�u0X�@� '4TX�0�pa3i1A3sQ25L�c��st�r�VR1%e�q0
��j1��O 2 �A�UEiy�.�‐� �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ�� qA!Pvs� 5	15aU ���?PŅ���ဝQG9A6�zS*�7�q�b5�1����Q��00	P(��V7]u�aitE1 ���ïp?7� !?�z���rbUQRB1P�M=�Qa9��H��QQ�25L�������Q���@L��8ܰ��y0�0\ry�"R2B�L�tN  ��w� �1D�q�2�qeR�5���_bx�3�X]1m1lcqP!1�a�E�Q� 5F����!5���@M-16 Q�� f���r��Q�e�� ��� PN�LT_`�1��i1��9453�p�@�e�|�b1l>�F1u*AY2�
��R8`�Q����RJ�J3�D}T� 85
Qg�/0�� *A!P�*A�Ð𫿽�Y2ǿپ6t�6=Q����Pȓ��� AQ� g�*ASt]1^u�a jrI�B����~�|I��b��yI�\m�Qb�I �uz�A�c3Apa9q� B6S��S��m����}�85`N�N�  �(M���f1����6����161��5�s`�SC��U��A�����5\set036c����10�y�#h8��a6��6��9r�2HS ���Er���W@}�a��I�lB� ��Y�ٖ�m�u�C������5�B��B��h `�F���X0���A:���C�M��AZ��@��4��6i����� e�O�- 	���f1��F ������1F�Y	���T6HL3��U66~`���Ur�dU�9D20Lf0 ��Qv� ��fjq��N� �����0v
� ��i	��	��72lqQ2�������� \chngmove.V���d���@2l_arf	�f~�� 6������9C�Z��0�~���kr41 S���0��V��t����8��U�p7nuqQ%��A]��V�1\�Qn�BJ�2W�E�M!5���)�#:�648��F�e50S�\� �0�=�PV���e�� ����E������m7shqQSH" U��)��9�!A��(����� ,�sq�ॲTR1!�L��,�60e=�4F�d����2��	 R-�� ���������Ж��4���LSR�)"�!lOA��Q�) %!� 16�
U/��2��"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D�� �5V��@2cVE��pȖ�T��pt갖�1L ~E�#�F�Q��9E�#Dce/��RT��59�� �	�A�EiR�������9\m20�20 ��+�-u�19r4�`� E1�=`O9`�1"ae��O�2��_$W}am41�4�3�/d?1c_std��1�)�!�`_T��r�_ 4\jdg�a�q�P J%!~`-�r�+bg8B��#c300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W �"PsA��e��� �t�i�P�W.�� c�FX.�e�kE1�4�44�~6\j4�443sj��r�j4up���\E19�h�PA�T�=:o�A Pf��coWo!\�[2a��2A;_2��QW2�bF�(�V11ă23�`��X5�Ra2�1�J*9�a:88�J9X�l5�m1a`첚��*���(85�& �������P6����R,52&A����,8fA9IfI50\u�z��OV
�v��}E֖J0���Y>� 16r�C �Y��;��1��L���A q�&ŦP1��vB)e��m�����1p� .�1D�q�27�F��KAREL Us�e S��FCTN<��� J97�FA+�� (�Q޵�p%�L)?�Vj9F?(�j�R�tk208 "Km�6Q�y�j��iæP�r�9�s#��v�kr;cfp�RCFt3����Q��kcctme��!ME�g����6�mWain�dV�� ��Cru��kDº�c��0�o����J�dt�F9 �»�.vrT�f�����E%�!��5�FR�j73B�K���UtER�HJ�O  J��# (ڳF���F�q� Y�&T��p�F�z��19�tkvBr���V�h�9p�E�y�<�k������p��;�v���"CT�� f����)�
І��)� V	�6���!��qFF ��1q���=�����O�@?�$"���$��je����TCP Aut��r�<520 H5n�J53E193��9��96�!8��9���	 �B574��5�2�Je�(�� Se%!Y�����u��ma>�Pqtool�ԕ������conr�el�Ftrol �Reliable��RmvCU!��H51������ a55�1e"�CNRE ¹I�c�&��it��l\sfutst "UTա��"X�\u��g@�i�6Q]V�0�B,Eѝ6A�  �Q�)C���X��Yf�hI�1|6s@6i��T6IU��vR�d�
$ae%1��2�C58�E6��8�Pv�iV4OFH�58SOeJ� mvBM6E~O58�I�0�E �#+@�&�F�0���F �P6a���)/++�</>N)0\tr1������P ,�qɶ�rmwaski�msk�a$A���ky'd�h	A	��P�sDispla�yIm�`v����J887 ("A��+Hyeůצprds�ҨIϩǅ�h�0pl�2"�R2��:�Gt�@��PRD�TɈ�r�C�@�Fm��D�Q�AscaҦ� V<Q&��bVvbrl�eې@��^Sp��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@�P�firmQ����P@p�2�=bk�6�r�3��6��tppl��PAL���O�p<b�ac�q 	��g1J�U�d�J��gait_9e��Y��&��Q���	�Sha�p��eratio�n�0��R674�51j9(`sGen@�ms�42-f��r�p`�5����2�rsgl��E��p�G���qF�20�5p�5S���Ձ�re�tsap�BP�O�\}s� "GCR��z�? �qngda�AG��V��st2ax�U��Aa]��bad��_�btputl�/�&�e���tpli1bB_��=�2.����5���cird�v�sqlp��x�hex���v�re?�Ɵx�key�v�pm��x�sus$�6�gcr���F������[�q27j9�2�v�ollis�mqSk�9O�ݝ� �(pl.���t��p!o��29$Fo8��cg�7no@�tptcls` CLS�o�b�F\�km�ai_
�s>�v�o	�t�b���ӿ�E�H��6�1e_nu501�[m���utia|$cal�maUR��CalMwateT;R51%�i=1]@-��/V� ���Z�� �fq1�9 "�K9E�L����2m�CLMTq�S#��3et �LM3!}t �F�c�nspQ�<c���c_moq��� ��c_e�����su��ޏ �_ �@�5�G�join�i�j��oX���&cWv	 �̆�N�ve��C�cl�m�&Ao# �|$fi�nde�0S�TD ter FiLANG���R��
��n3���z0Cen���r, ������J����� � ��K��Ú�=���_�����r� "FNCDR�� 3��f��tguid�䙃N�."��J�tq�� ��� ����������J����_������c��	m��Z��\fndrA.��n#>
B2p��>Z�CP Ma������38A��� c��6� (���N�B���@���� 2�$�81�B�m_���"ex� z5�.Ӛ��c��0bSа�efQ���	��RBT;�OPTN �+#Q� *$�r*$��*$r*$%/ s#C�d/.,P�/0*ʲDPN��$����$*�Gr�$k E�xc�'IF�$MA�SK�%93 H5��%H558�$548 H�$4-1�$�d�#1(�$�0 E�$���$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9j0�"M�49�4  ���4�4tpsh���4�P�4- DQ�� �3�Q�4�R�4�pR@%0�2�r�4.b
E\���5�A�4��3adq}\�5K979":E��ajO l "DQ ^E^�3i�Dq ��4�ҲO ?R�? ��q@�5��T��3rAq�OF�Lst�5~��7p�5`��REJ#�2�@av^E�ͱ�F���4��.�5y� N� �2il(iqn�4��31 JH1��2Q4�251ݠ�4r'mal� �3)�RE o�Z_�æOx����4��8^F�?onorTf��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱ�4$�REM���4yݱ"u<@�RER5932fO��47Z��5lity�,�U��e"Dil�\�5��o ��79�87�?�25 �3hk910�3��FE�0�=0P_�Hl\mhm �5��qe�=$�^��
E��u�IAympt�m�U��BU��vst e�y\�3��me�b�Dv I�[�Qu�:F�Ub�*_0�
E,�su��_	 Er��ox���4huse�E-�?�sn�������FE��,�Gbox�����c݌ ,"�������z���M��g��pdspw )�	��9���b���(��1���c�� Y�R�� �>�P���W�@�������'�0ɵ��[��͂��� � � ,�@�� �A�bu�mpšf��B*�BCox%��7Aǰ60�pBBw���MC� (6��,f�t I�s� ST��*��}B������w��"BBF�
�>�`���)��\�bbk968 "��4�ω�bb�9�va69����etb�Š��X�����ed�	�F��u�f� �s�ea"������'�\���,���b�ѽ�oH6�H�
�x�$�f����!y���Q[�! toperr�fd� �TPl0o� Rec�ov,��3D��R/642 � 0��C@�}s� N@��(U�rro���yu2r���  �
 � ����$$CL~e� ������������$z�_�DIGIT��������.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�o$j��+c:PR�ODUCTM�0\�PGSTKD��V�&ohozf99��D����$FEAT_INDEX���xd�� � 
�`ILEC�OMP ;����#��`�cSET�UP2 <�e��b�  N ��a�c_AP2BC�K 1=�i G �)wh0?{%&c����Q�xe% �I�m���8� �\�n����!���ȏ W��{��"���F�Տ j���w���/�ğS�� �������B�T��x� �����=�үa����� �,���P�߯t���� ��9�ο�o�ϓ�(� :�ɿ^���Ϗϸ� G���k� �ߡ�6��� Z�l��ϐ�ߴ���U� ��y����D���h� �ߌ��-���Q����� �����@�R���v�� ��)�����_����� *��N��r�� 7��m�&��3\�i
pP }2#p*.VRc�*��� /��PC/1/�FR6:/].��/+T�`�/�/F%��/�,�`r/?�*#.F�8?	H#&?�e<�/�?;STM� �2�?�.K �?�=�iPenda�nt Panel�?;H�?@O�7.O�?8y?�O:GIF�O�O��5�OoO�O_:JPG _J_�56_�O_�_��	PANEL1'.DT�_�0�_�_�?O�_2�_So�W Ao�_o�o�Z3qo�o@�W�o�o�o)�Z4�o�[�WI��
�TPEINS.XSML��0\����qCustom� Toolbar�	��PASSW�ORDyFR�S:\L�� %�Password Config�� �֏e�Ϗ�B0��� T�f����������O� �s������>�͟b� �[���'���K��� �����:�L�ۯp��� ��#�5�ʿY��}�� $ϳ�H�׿l�~�Ϣ� 1�����g��ϋ� ߯� ��V���z�	�s߰�?� ��c���
��.��R� d��߈���;�M��� q������<���`��� ����%���I������ ��8����n��� !��W�{" �F�j|�/ �Se��/�/ T/�x//�/�/=/�/ a/�/?�/,?�/P?�/ �/�??�?9?�?�?o? O�?(O:O�?^O�?�O �O#O�OGO�OkO}O_ �O6_�O/_l_�O�__ �_�_U_�_y_o o�_ Do�_ho�_	o�o-o�o Qo�o�o�o�o@R �ov��;�_ ���*��N��G� �����7�̏ޏm�� ��&�8�Ǐ\�돀�� !���E�ڟi�ӟ��� 4�ßX�j�������� įS��w������B��#��$FILE_�DGBCK 1=���/���� ( �)�
SUMMARY�.DGL���MD�:�����Di�ag Summa�ry��Ϊ
CONSLOG��������D�ӱConso?le logE�ͫ���MEMCHECCK:�!ϯ���X��Memory D�ata��ѧ�{�)��HADOW�ϣϵ�J���Sh�adow Cha�ngesM�'�-��)	FTP7�Ф�3ߨ���Z�mment TBD���ѧ0=4)ET?HERNET��������T�ӱEth�ernet \�f�iguratio�nU�ؠ��DCSV�RF�߽߫������%�� veri?fy all��'��1PY���DIF�F�����[���%=��diff]�������1R�9�K���c ���X��CHGD������cB��r����2Z8AS� ��GD���k��qz��FY3b8I[� �/"GD���s/�����/*&UPDATES.� �/��?FRS:\�/�-�ԱUpdate?s List�/���PSRBWLD.CM(?���"<?�/�Y�PS_ROBOWEL��̯�?�?� �?&�O-O�?QO�?uO OnO�O:O�O^O�O_ �O)_�OM___�O�__ �_�_H_�_l_o�_�_ 7o�_[o�_lo�o o�o Do�o�ozo�o3E �oi�o���R �v���A��e� w����*���я`��� ������O�ޏs�� ����8�͟\����� '���K�]�쟁���� 4���ۯj������5� įY��}������B� ׿�x�Ϝ�1���*� g�����Ϝ���P��� t�	�ߪ�?���c�u� ߙ�(߽�L߶��߂� ��(�M���q� �� ��6���Z������%� ��I���B�����2�����h����$FoILE_� PR� ���������MDO?NLY 1=.��? 
 ���q ����������~ %�I�m �2��h��!/ �./W/�{/
/�/�/ @/�/d/�/?�//?�/ S?e?�/�??�?<?�? �?r?O�?+O=O�?aO �?�O�O&O�OJO�O�O �O_�O9_�OF_o_
?VISBCKL6>[*.VDv_�_>.PFR:\�_�^�.PVisio�n VD file�_�O4oFo\_joT_ �oo�o�oSo�owo �oB�of�o� +������� +�P��t������9� Ώ]�򏁏��(���L� ^�������5���ܟ k� ���$�6�şZ���~�����
MR_�GRP 1>.�L��C4  B���	 W������*u����RHB ���2 ��� ��� ���B����� Z�l���C���D��������Ŀ��K�G��J���I��6�T���F�5U�P�����ֿ �E�M.G��E$��;n���:G��@O����@�5P@����fZ�@���W@���*λ?� F@ ��������J��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<,6\b�π+�&�(�a�L߅�p�A��A��߲�v���r� �����
�C�.�@�y� d���������������?�Z�lϖ�BH�� �Ζ��������
0�PS@�P��TW��ܿ� �B���/ ��@�33�:��.�gN�UU�U�U��q	>u.�?!rX���	�-=[z��=�̽=V�6<�=�=�ߎ=$q������@8�i7G���8�D�8@9!�7�:�����D�@ D��� Cϥ��C������'/0-�� P/����/N��/r��/ ���/�??;?&?_? J?\?�?�?�?�?�?�? O�?O7O"O[OFOO jO�O�O�O�O�гߵ� �O$_�OH_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooVohoSo�owo�o �i��o�o�o��) ;�o_J�j�� �����%��5� [�F��j�����Ǐ�� �֏�!��E�0�i� {�B/��f/�/�/�/�� �/��/A�\�e�P��� t��������ί�� +��O�:�s�^�p��� ��Ϳ���ܿ� ��O H��o�
ϓ�~ϷϢ� ���������5� �Y� D�}�hߍ߳ߞ����� ���o�1�C�U�y� �߉���������� ��-��Q�<�u�`��� ������������ ;&_J\��� �������ڟ�F �j4������ ���!//1/W/B/ {/f/�/�/�/�/�/�/ �/??A?,?e?,φ? P�q?�?�?�?�?O�? +OOOO:OLO�OpO�O �O�O�O�O�O_'__ K_�o_�_�_�_l��_ 0_�_�_�_#o
oGo.o koVoho�o�o�o�o�o �o�oC.gR �v�����	� ��<�`�*<�� `�����ޏ��)� �M�8�q�\������� ˟���ڟ���7�"� [�F�X���|���|?֯ �?�����3��W�B� {�f�����ÿ������ ���A�,�e�P�u� ��b_�����Ϫ_��� ��=�(�a�s�Zߗ�~� �ߦ�������� �9� $�]�H��l���� ��������#��G�Y�  �B�������z����� ��
ԏ:�C.gR d������	 �?*cN�r �����/̯&/ �M/�q/\/�/�/�/ �/�/�/�/?�/7?"? 4?m?X?�?|?�?�?�? �?��O!O3O��WOiO �?�OxO�O�O�O�O�O _�O/__S_>_P_�_ t_�_�_�_�_�_�_o +ooOo:oso^o�o�o p��o�� ��$�� o�o�~�� �����5� �Y� D�}�h�������׏ ����
�C�.�/v� <���8������П�� ��?�*�c�N���r� �������̯��)� �?9�_�q���JO��� ��ݿȿ��%�7�� [�F��jϣώ��ϲ� ������!��E�0�i� T�yߟߊ��߮��߮o �o��o>�t�> ��b����������� +��O�:�L���p��� ����������' K6oZ�Z�|�~� ����5 Y Di�z���� ��/
//U/@/y/ @��/�/�/�/���/^/ ???Q?8?u?\?�? �?�?�?�?�?�?OO ;O&O8OqO\O�O�O�O �O�O�O�O_�O7_���$FNO ����VQ��
F0fQ �kP FLAG8�(�LRRM_CHK�TYP  WP�\�^P�WP�{Q{OM�P_MIN�P�����P�  �XNPSSB_C�FG ?VU ��_����S ooIUTP_D�EF_OW  ���R&hIRCO�M�P8o�$GENOVRD_DO�Vs�6�flTHR�V� d�edkd_EN�BWo k`RAV�C_GRP 1@�WCa X"_�o_ 1U<y�r �����	��-� �=�c�J���n����� ���ȏ����;�"��_�F�X���ibROUr�`FVX�P��&�<b&�8�?��埘�������  D?�јs�6��@@g�B�7�p�p)�ԙ���`SMT�cG�mM���� �LQ�HOSTC�R1H����P��at�kSM��f�\����	127.0z��1��  e�� ٿ�����ǿ@�R��d�vϙ�0�*�	anonymous��`���������[�� � �����r� ���ߨߺ�����-�� �&�8�[�I�π�� �����1�C�� W�y���`�r������� ��������%�c�u� J\n������� ��M�"4FX ��i������ 7//0/B/T/�� �m/��/�/�/? ?,?�/P?b?t?�?�/ �?��?�?�?OOe/ w/�/�/�?�O�/�O�O �O�O�O=?_$_6_H_ kOY_�?�_�_�_�_�_ 'O9OKO]O__Do�Oho zo�o�o�o�O�o�o�o 
?o}_Rdv� ��_�_oo!�Uo *�<�N�`�r��o���� ��̏ޏ�?Q&�8��J�\���>�ENT {1I�� P!�.��  ����՟ ğ�������A��M� (�v���^�����㯦� �ʯ+�� �a�$��� H���l�Ϳ�����ƿ '��K��o�2�hϥ� ���ό��ϰ����� ��F�k�.ߏ�R߳�v� �ߚ��߾���1���U���y�<�QUIC�C0��b�t����1 �����%���2&����u�!ROUT�ERv�R�d���!�PCJOG�����!192.16?8.0.10��w�NAME !��!ROBOT�p�S_CFG 1�H�� ��Auto-st�arted�tFTP����� �� 2D��h z����U�� 
//./�v���/ ���/�/�/�/�/� !?3?E?W?i?�/?�? �?�?�?�?�?��� AO�?eO�/�O�O�O�O �?�O�O__+_NO�O J_s_�_�_�_�_
OO .OoB_'ovOKo]ooo �oP_>o�o�o�o�oo �o5GYk}�_ �_�_��8o�� 1�C�U�$y������� �ӏf���	��-�?� ����Ə���ϟ �����;�M�_� q���.�(���˯ݯ� �P�b�t�����m��� ������ǿٿ����� !�3�E�h��{ύϟ� �����$�6�H�J�/� ~�S�e�w߉ߛ�jϿ� �������*߬�=�O��a�s��YT_ER�R J5
���P�DUSIZ  j��^J����>��?WRD ?t���  guest}��%�7��I�[�m�$SCDMNGRP 2Ktw�������V$�K�� 	�P01.14 8~��   y�����B   � ;����� ����������
 �������?�����~����C.gR|����  i  ��  
��������� +�������
���l �.r���"�l��� m
d����|��_GROU��]L�� �	�����07EQUPD'  	պ�J��TYa ����T�TP_AUTH �1M�� <!iPendany���6�Y!K?AREL:*��
-KC///A/ �VISION �SETT�/v/� "�/�/�/#�/�/
? ?Q?(?:?�?^?p>�CTRL N�����5�
�F�FF9E3�?��FRS:DEFA�ULT�<FA�NUC Web �Server�:
 �����<kO}O�O�O��O�O��WR_CONFIG O��� �?��IDL_CPU_PC@��B��7P�BHUMIN(\��<T?GNR_IO�������PNPT_S_IM_DOmVw[�TPMODNTO�LmV �]_PRT�Y�X7RTOLNK 1P����_o�!o3oEoWoio�RMA�STElP��R�O�_CFG�o�iUO���o�bCYCLE��o�d@_ASG s1Q����
 ko ,>Pbt��� ������sk�bNUM����K@�`�IPCH�o��`R?TRY_CN@oR<��bSCRN����Q��� �b�`�b�R���Տ��$J�23_DSP_E�N	����OB�PROC�U�iJ[OGP1SY@��?8�?�!�T��!�?*�POSRE��zVKANJI_@�`��o_�� ��T�L��6͕����CL_�LGP<�_���EYL_OGGIN�`�����LANGU�AGE YF7ReD w���LG��YU�?⧈�x� ������=P��'�0��$ NM�C:\RSCH\�00\��LN_D?ISP V��
�0�������OC�R.R�DzVTA{�OGB?OOK W
{��`i��ii��X������ǿٿ�����"��6	h������e�?�G_BUF/F 1X�]��2	աϸ������� ����!�N�E�W߄� {ߍߺ߱�����������J���DCS� Zr� =����^�+�ZE������|��a�IO 1[
{G ُ!� �!� 1�C�U�i�y������� ��������	-A Qcu�����z��EfPTM  �d�2/ASew �������/ /+/=/O/a/s/�/�/���SEV���.�TYP�/0??y͒�RS@"�|�×�FL 1\
������?�?�?�?0�?�?�?/?TP6���">�NGNA�M�ե�U`�UPSF��GI}�𑪅mA�_LOAD�G �%�%DF_�MOTN���O�@MAXUALRM<���J��@sA�Q����(WS ��@C �]m�-_����MP2�7�^
{k ر�	�!P��+ʠ�;_/��Rr�W�_�WU�W�_�� �R	o�_o?o"ocoNo so�o�o�o�o�o�o�o �o;&Kq\� x������� #�I�4�m�P���|��� Ǐ���֏��!��E� (�i�T�f�����ß�� ӟ���� �A�,�>� w�Z�������ѯ���� د���O�2�s�^� ������Ϳ���ܿ��'��BD_LDXD�ISAX@	��ME�MO_APR@E {?�+
 �  *�~ϐϢϴ�����������@ISC 1_�+ ��IߨT�� Q�c�Ϝ߇��ߧ��� ��w����>�)�b�t� [����{������� ���:���I�[�/��� ���������o����� 6!ZlS�� s����2� AS'�w��� �g��.//R/d/��_MSTR �`�-w%SCD 1am͠L/�/H/�/�/ ?�/2??/?h?S?�? w?�?�?�?�?�?
O�? .OORO=OvOaO�O�O �O�O�O�O�O__<_ '_L_r_]_�_�_�_�_ �_�_o�_�_8o#o\o Go�oko�o�o�o�o�o �o�o"F1jU g������� ��B�-�f�Q���u�𮏙�ҏh/MKCF/G b�-㏕"�LTARM_��c�L�� �σQ�N�<�METP�UI�ǂ���)N�DSP_CMNT�h���|�  d�.��ς�ҟܔ|�_POSCF�����PSTOL 1e�'�4@�<#�
 5�́5�E�S�1�S�U� g�������߯��ӯ� ��	�K�-�?���c�u������|�SING_?CHK  ��;�/ODAQ,�f��Ç���DEV 	�L�	MC:!�HOSIZEh��-��TASK %6��%$123456�789 �Ϡ��T�RIG 1g�+ l6�%���ǃ��0���8�p�YP[� ���EM_INF �1h3� �`)AT&F�V0E0"ߙ�)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ�����ԁH�����A���A�I�q�,��|����  ���ߵ�����J��� n������W������� ����"����X�� /����e���� ��0�T;x�= �as��/�,/ c=/b/�/A/�/�/ �/�/��?��� ^?p?#/�?�/�?s?}/ �?�?O�?6OHO�/lO ?1?C?U?�Oy?�O�O 3O _�?D_�OU_z_a_��_�ONITORG ?5�   �	EXEC1TɃ�R2�X3�X4�XQ5�X���V7�X8�X9Ƀ�RhBLd�RLd �RLd�RLd
bLdbLd "bLd.bLd:bLdFbLcU2Sh2_h2kh2whU2�h2�h2�h2�hU2�h2�h3Sh3_h�3�R�R_GRP?_SV 1in����(����C?B�PP�A4�>%���gY�>r3��x�_D=R^���PL_NAME� !6��p�!�Default� Persona�lity (from FD) ��RR2eq 1j)TUX)TX��q��X dϏ8�J�\� n���������ȏڏ� ���"�4�F�X�j�|������2'�П��� ��*�<�N�`�r��<��������ү������,�>�P�b� �R�dr 1o�y �\��, �3��~�� @D�  ��?�����?䰺�㱏A'�6����;��	lʲ	 �xJ����� ��< �"�� ��(pK�K� ��K=*�J����J���J�V���Z�����rτ́p@j��@T;f���f���ұ]�l��I�o��������������b��3���o�  ��`�>�����bϸ�z��{Ꜧ���Jm��
� B�H�˱]����q�	� p��  P�pQ�p�>�p|  Ъ�g����c�	'� �� ��I� ��  ����:��È
�È=����"�nÿ�	�ВI�  �n @@B�cΤ�\��ۤ���q�y�o�N���  �'�����@2��@�����/��C��C�C�@� C������
��A�W�@<�*P�R�
h�B�b�A��j�����:����Dz۩��߹������j��( ?�� -��C�`��'�7�����q��Y����� �?�ff ��gy ����o��:a��
>+�  PƱj�(����7	����|�?���xZ�p<
6b�<߈;܍��<�ê<� �<�&Jσ�A�I�ɳ+���?ff�f?I�?&�k�@��.��J<?�`�q�.�˴ fɺ�/��5/���� j/U/�/y/�/�/�/�/��/?�/0?q��F �?l??�?/�?+)��?�?�E�� E��I�G+� F� �?)O�?9O_OJO�OXnO�Of�BL޳B� ?_h�.��O�O��%_�O L_�?m_�?�__�_�_x�_�_�
�h�Îg>��_Co�_`goRodo�o�GA�ds�q�C�o�o�o|����$]Hq�m��D��pC����pCHmZZ7t����6q�q��ܶN'�3�A�A�AR1�AO�^?�$��?�K/�±
�=ç>�����3�W
=�#�\W��e��9������{����<���(�B��u��=B�0�������	L��H�F�G����G��H��U`E���C��+���I#��I��HD��F��E��R�C�j=��
�I��@H�!�H�( E<YD0q�$��H� 3�l�W���{������� �՟���2��V�A� z���w�����ԯ���� ����R�=�v�a� �����������߿� �<�'�`�Kτ�oρ� �ϥ��������&�� J�\�G߀�kߤߏ��� ��������"��F�1� j�U��y������� �����0��T�?�Q�t���(���3/�E����u�������q3�8�x����q4Mgs�&IB+2D�a���{�^ ^	������u%P2P7Q4_A���M0bt��R�������/   �/�b/P/�/ t/�/ *a)_3/�/�/�%1a?�/?;?8M?_?q?  �?�/��?�?�?�?O 2 �F�$�vGb��/�A��@�a�`�qC��C@�o�Ot���K�F� DzH@��� F�P D�!��O�O�ys<O!_�3_E_W_i_s?��W�@@pZ�42�2!2~
 p_�_�_�_	oo -o?oQocouo�o�o�o��o��Q ��+���1��$MSK�CFMAP  ��5� ��6�Q�Q"~�cONR�EL  
�q3�bEXCFE�NB?w
s1uXqF�NC_QtJOGO/VLIM?wdIpMr]d�bKEY?w�u]�bRUN�|�u��bSFSPDT�Y�avJu3sSIG�N?QtT1MOT��Nq�b_CE_�GRP 1p�5s\r���j����� T��⏙������<� �`��U���M���̟ ��🧟�&�ݟJ�� C���7�������گ��������4�V�`TC�OM_CFG 1�q}�Vp�����
�P�_ARC_\r�
jyUAP_CP�L��ntNOCHE�CK ?{ 	r��1�C� U�g�yϋϝϯ����������	��({NO_?WAIT_L�	u6M�NTX�r{�[�m�_ERRY�29sy3� &�������r�c� �촯T_MO��t��,�  �<$�k�3�P�ARAM��u{�	�[���u?��� =9@345678901��&��� E�W�3�c�����{�������������=�UM_RSP�ACE �Vv��$ODRDSP����jxOFFSET�_CARTܿ�D�IS��PEN_FILE� �q��c����OPTION_�IO��PWOR�K v_�ms �P(�R�Q
�j.j	 ��Hj&�6$� RG_DS�BL  �5Js��\��RIENTkTO>p9!C��P�qfA� UT_SIM_D
r�b� �V� LCT w�w�bc��U)+$_P�EXE�d&RAT�p �vju�p��2X�j�)TUX)TX�>##X d-�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?O�H2�/oO �O�O�O�O�O�O�O�O_]�<^O;_M___q_ �_�_�_�_�_�_�_o����X�OU[�o(��(���$}o�, ���IpB` @D�  &Ua?�[cAa?p]a�]�DWcUa쪋l;��	lmb�`��xJ�`��p���a�<; ��`� ��b���H(��H3k7�HSM5G�22�G���Gp
��
���'|��KCR�>�>q�Gs�uaT�3���  �4spBpyr  ]�o�*SB_�����j]��t�q� ��rna ��,���6  U��PQ��|N�M�,k���	�'� � ���I� �  {��%�=��ͭ�迋ba	���I  �n @� �~���p�����r��N	 W�  '!�o�:q�pC	 C�@�@sBq�|��� m�
S�!�h@ߐ�n�����*�B	 �A8���p� �-�qbz��P��t�_�������( �� -��恊�n�ڥ[A]Ѻ�b4�'!�5�(p �?�fAf� ��
����O�Z�R*�85�z���>N΁  Pia��(5� ��@���ک�a�c�dF#/?��5�x��*��<
6b<߈�;܍�<�ê�<� <�&�o&�)�A�lcΐIƾ*�?fff?�?y&c���@�.u��J<?�`�� Yђ^�nd��]e��[g ��Gǡd<����1�� U�@�y�dߝ߯ߚ��� �߼�	���-�������&��"�E�� E���G+� F� ������������&���J�5��bB��A T�8�ђ��0�6���>� ��J�n�7��[mx�0��h��1��>�M�I`
�@��A�[��C-�)��?���� /�
YĒ��Jp��vav`#CH/�������}!@I�Y�'��3A�A�AR�1AO�^?�$��?����±�
=ç>�����3�W
=�#�����+e��ܒ������{�����<��.(��B�u��=�B0�������	�*H�F��G���G���H�U`E����C�+�-I#��I��HD��F��E���RC�j=U>
�I��@H��!H�( E<YD0/�?�?�? �?�?O�?3OOWOBO TO�OxO�O�O�O�O�O �O_/__S_>_w_b_ �_�_�_�_�_�_�_o o=o(oaoLo�o�o�o �o�o�o�o�o' $]H�l��� ����#��G�2� k�V���z���ŏ��� ԏ���1��U�g�R� ��v�����ӟ��������-��(���������a�����Q�c�,!3�8��}���,!4Mgs8����ɢIB+կ���a���{� ��A�/�e�S���w�J�P!�P��������7��ӯ�ϑ�R9�Kτ�oχϓϥ�  ���χ���� )��M������z���{߉ߛ���ߒߤ�p������  )�G�q�_���2� F�$�&Gb	���n�[ZjM!C�s�@j/�A�S�~=�F� Dz����� F�P DC��W����)������������x?̯��@@
9�R=�=��=��
 v��� ����*<pN`�*P �������1��$PA�RAM_MENU� ?-���  DEFPULSEl�	WAITTM�OUT�RCV�� SHEL�L_WRK.$CUR_STYL�;,OPT�/�PTB./("C�R?_DECSN��� ,y/�/�/�/�/�/�/ ?	??-?V?Q?c?u?��?�USE_PR_OG %�%�?\�?�3CCR������7_HOST !�!�44O�:AT̰�?PCO)ARC|�O�;_TIME��XB�  �GD�EBUGV@��3G�INP_FLMS�K�O�IT`��O�EP+GAP �L��#[�CH�O�HTYPE
����?�?�_�_ �_�_�_oo'o9obo ]ooo�o�o�o�o�o�o �o�o:5GY� }����������1�Z��EWOR�D ?	7]	�RS`�	PNS2�$��JOE!>��TEs@WVTRA�CECTL 1xv-�� ������ɆDT� Qy-����D � �� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� T�(�v����������� ����*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_j��_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�_����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv��������//"#�$P�GTRACELE�N  #!  ���" ��8&_UP z����g!o S!�h 8!_CFG {g%Q#"!x!��$J �#|"DEF�SPD |�,l!!J �8 IN �TRL }�-�" 8�%�!PE_C�ONFI� ~g%O�g!�$�%��$LID�#�-~74GRP 1�7�Q!�#!A ����&ff"!A+�33D�� D]�� CÀ A@+6�!�" d�$�9�9�*1*0� 	 �+9�(�&�"�? ´	C�?�;B@3AO�?�OIO3OmO"!>�T?�
5�O�O�N��O =��=#�
�O_�O_J_5_ n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_Roxoco�o �o�o�o�o�o�o�>)bM��;
�V7.10bet�a1�$  �A�E�rӻ��A " �p?!G�^�q>���r��0��q�ͻqBQ��qA\�p�q�4�q*�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏� ��4��1�j�U���y� ����֟������0� �T�?�x�c������� ү����!o�,�ۯP� ;�M���q�����ο�� �ݿ�(��L�7�p�x+9��sF@ �� �ͷϥ�g%������ +�!6I�[߆������� �ߠ���������!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ���=(aL ^������ �'9$]�Ϛ��� ��������/<� 5/`�r߄ߖߏ/>�/ �/�/�/�/?�/1?? U?@?R?�?v?�?�?�? �?�?�?O-OOQO<O uO`O�O�O�O�O���O _�O)__M_8_q_\_ n_�_�_�_�_�_�_o �_7oIot���o�o ���o�o�o(/!L/ ^/p/�/{*o��� ������A�,� e�P�b���������� Ώ��+�=�(�a�L� ��p������Oߟ񟠟 � �9�$�]�H���l� ~�����ۯƯ���#� No`oro�on��o�o�o �oԿ���8J\ ng����vϯϚ��� ����	���-��Q�<� u�`�r߫ߖ��ߺ��� ����;�M�8�q�\� ��������z������ %��I�4�m�X���|� ����������:�L� ^���Z�������� ���$�6�H�S wb����� ��//=/(/a/L/ �/p/�/�/�/�/�/? �/'??K?]?H?�?�� �?�?f?�?�?�?O�? 5O OYODO}OhO�O�O �O�O�O�O&8J4_ F_����_�_��_ �_"4-o�O*oco No�oro�o�o�o�o�o �o)M8q\ �������� �7�"�[�m��?���� R�Ǐ���֏�!�� E�0�i�T���x����� ���_$_V_ �2�l_�~_�_�����R�$P�LID_KNOW�_M  �T������SV� ��U͠�U��
��.� ǟR�=�O�����mӣ�M_GRP 1�T�!`0u��T@ٰ)o�ҵ�
���P зj��`���!�J� _�W�i�{ύϟϱ���`������߱�MR��Ņ��T��s�w�  s��ߠ޴߯߅��ߩ� ������A���'�� ����������� ��=���#����������}������S��ST^��1 1��U# ����0�_ A  .��,>Pb�� ������3 (iL^p���(��2*��'�<-/3/)/;/M/4f/x/�/�/�5�/�/�/�/6 ??(?:?7S?e?w?�?8�?�?�?�?~MAD  d�#`PARN_UM  w�\%OSCH?J ME�
�G`A�Iͣ�EUP�D`OrE
a�OT_CMP_��B@�P@�'˥TER_C;HK'U��˪?R�$_6[RSl�¯��_#MOA@�_�U_�_RE�_RES_G � �>�oo8o+o\o Oo�oso�o�o�o�o�o@�o�o�W �\�_ %�Ue Baf�S�  ����S0��� �SR0��#��S�0>� ]�b��S�0}������R�V 1�����rB@�c]��t�(@�c\����D@�c[�$���RTHR_INRl�DA��z˥d,�MASS9�� ZM�MN8�k�M�ON_QUEUE� ���˦��x� URDNPUbQN{�P[��END���_ڙ�EXE�ڕ�@BE��ʟ��OPTIO�Ǘ�[��PROGR�AM %��%�ۏ�O��TASK�_IAD0�OCFG� ���tO��ŠD�ATA���Ϋ@��27�>�P�b�t� ��,�����ɿۿ������#�5�G���INFOUӌ�������� �Ͽ���������+� =�O�a�s߅ߗߩ߻�@�������^�jč�� yġ?PDIT� �ίc���WE�RFL
��
RG�ADJ �n�A	����?����@���?IORITY{�QV}���MPDSPH������Uz����O�TOEy�1�R�� (!AF4�E��P]���!tc�ph���!ud|��!icm���ݏ6�XY_ȡ��R��ۡ)� *0+/ ۠�W :F�j���� ��%7[B��*��PORTT#�BC۠�����_CARTREP�
�R� SKSTA�z��ZSSAV����n�	2500H863���r�$!�U�R����q��n�}/�/�'� URGeE�B��rYWF� #DO{�rUVWV��$��A�WRUP_DELAY �R�>�$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?3A_QSKIP!�n�;l#x 	1/+O + OROdOvO9Hn��O �G�O�O�O�O�O_�O _D_V_h_._�_z_�_ �_�_�_�_
o�_.o@o Roovodo�o�o�o�o �o�o�o*<L�r`���n��$�RCVTM���]��pDCR!�L�ЈqB��C�*J�C$�>��$ >5?-;���04M¹�O���ǃ�������~��9On�Y��<
6b<߈�;܍�>u.��?!<�& {�b�ˏݏ��8���� �,�>�P�b�t����� ����Ο���ݟ�� :�%�7�p�S������ ʯܯ� ��$�6�H� Z�l�~�������ƿ�� �տ���2�D�'�h� zϽ��ϰ��������� 
��.�@�R�d�Oψ� �߅߾ߩ������� ��<�N��r���� ����������&�8� #�\�G�����}����� ������S�4FX j|������ ���0T?x �u����'/ /,/>/P/b/t/�/�/ �/�/�/�/�?�/(? ?L?7?p?�?e?�?�? ��?�? OO$O6OHO ZOlO~O�O�O�?�?�O �O�O�O __D_V_9_ z_�_�?�_�_�_�_�_ 
oo.o@oRodovo�X��qGN_ATC �1�� AT&FV0E/�� ATDP/6/9/2/9�h�ATA�n,�AT%G1%B�960/�++U+�o,�aH,�q�IO_TYPE � �u�sn_�oR�EFPOS1 1}�P{ x�o�Xh_�d_��� ��K�6�o�
���.�ාR����{{2 1�P{���؏V�ԏxz����q3 1���$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����<�>��S6 1�ѯ����/�����ѿO�S7 1�f�x���ĿB��-�f��S8 1� ����Y�������y��SMASK 1��P  
9�G��XNOM���a~߈�~�qMOTE  h��~t��_CFG ᢥ����рrPL_�RANG�ћQ��POWER ��e���SM_DRYPRG %i��%��J��TART� �
�X�UME_PRO'�9��~t�_EXEC_EN�B  �e��GS�PD������c��T3DB���RM���MT_!�T����`OBOT_NA_ME i�����iOB_ORD_�NUM ?
��\qH863�  �T���������bPC_TIMoEOUT�� x�`oS232��1��k� LTEA�CH PENDA1N �ǅ�}����`Mainte�nance Co#ns�R}�m
"{�d?KCL/Cg��Z� ��n� ?No Use}�8	��*NPO��Ѯ����(C7H_L��������	�mMAVA#IL��{��ՙ��SPACE1 2��| d��(>��&���p��M,?8�?�ep/ eT/�/�/�/�/�W/ /,/>/�/b/�/v?�? Z?�/�?�9�e�a�=? ?,?>?�?b?�?vO�O�ZO�?�O�O�Os�2�/O*O<O�O`O �O�_�_u_�_�_�_�_[3_#_5_G_Y_o }_�_�o�o�o�o�o[4.o@oRodovo $�o�o����"�	�7�[5K]o� �A����	�̏�?�&�T�[6h�z��� ����^�ԏ���&�� ;�\�C�q�[7���� ����͟{���"�C�@�X�y�`���[8�� ��Ưدꯘ��0�?π`�#�uϖ�}ϫ�[Gw �i� ��:�
G� ���� $�6�H�Z�l�~ߐ��8  ǳ�����߈��d(���M�_�q�� ����������?� ��2�%�7�e�w����� ��������������� !�RE�W����� �����?�Q `�� @ 0��ߖrz	�V_�����
/ L/^/|/2/d/�/�/�/ �/�/�/?�/�/�/*? l?~?�?R?�?�?�?�?@�?�?�?2O�?
���O[_MODE � �˝IS �"��vO,*ϲ��O-_��	M_v_#dCWORK_AD�M�-��%aR  ���ϰ�P{_�P_?INTVAL�@�����JR_OPTI[ON�V �EBp�VAT_GRP �2����#(y_Ho �e_vo �o�oYo�o�o�o�o�o *<�bOoNDp w������	� ��?�Q�c�u����� /���ϏᏣ����)� ;���_�q��������� O�ɟ���՟7�I� [�m�/�������ǯٯ 믁��!�3���C�i� {���O���ÿտ��� ϡ�/�A�S�e�'ω� �ϭ�oρ������� +�=���a�s߅�Gߕ� �����ߡ���'�9� K�]��߁����y� ���������5�G�Y���E�$SCAN_GTIM�AYuew��R �(�#(�(�<0.a+aPaP
TqA>��Q��oX�����OO�2/��:	d/JaR��WY��^��p�^R^	r  P���� � � 8�P�	�D��GYk} ��������Qp/@/R/x/)P;�o\T���Qpg-�t�_DiKT��[  � lv%��� ���/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OWW �#�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o lO~Od+No`oro�o�o �o�o�o�o�o& 8J\n����8��u�  0�"0g �/�-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q�����$o ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E��� ��Do��������ҿ� ����,�>�P�b�t� �ϘϪϼ���������w
�  58�J�\� n߀ߒߜկ������� ��	��-�?�Q�c�u�p����� �� -����� �2�D�V�@h�z�������������������& ���%	123�45678�" +	��/� ` r������� �(:L^p ������� / /$/6/H/Z/l/~/� �/�/�/�/�/�/? ? 2?D?V?h?�/�?�?�? �?�?�?�?
OO.O@O o?dOvO�O�O�O�O�O �O�O__*_YON_`_ r_�_�_�_�_�_�_�_ ooC_8oJo\ono�o �o�o�o�o�o�oo "4FXj|���������	���s3�E�W�{�C�z  Bp��  � ��2���z��$SCR_GRP� 1�(�U8(�\x^ �@  �	!�	 ׃�� �"�$� ��-��+���R�w����D!~�����#����O����M-10i�A 890990�5 Ŗ5 M61CA >4��Jׁ
� ���0�����#�1�	"�z���О���¯Ҭ � ��c���O�8�J� ������!�����\ֿ��B�y����������A��$�  !@��<� �R�?��d����Hy�u�O���F@ F�`�§�ʿ �϶�������%��I� 4�m��<�l߃ߕ��߹�B���\���� 1��U�@�R��v�� ����������;���*<=�
F���?�<d�<�>7�����s@�:��� B����ЗЙ���EL�_DEFAULT�  �����B�MIP�OWERFL  ��$1 WFD�O $��ER�VENT 1������"�pL!�DUM_EIP���8��j!AF�_INE �=�!'FT���9!��4 ��[�!RPC_MAIN\>�J�n'VISw=���o!TP�PU��	d�?/!
PM�ON_PROXY@/�e./�/"Y/��fz/�/!RDMO_SRV�/�	g�/�#?!R C?�h,?o?!
pM�/��i^?�?!RLSgYNC�?8�8�?>O!ROS�.L�4�?SO"wO�#DO VO�O�O�O�O�O_�O 1_�OU__._@_�_d_ v_�_�_�_�_o�_?o�ocoiICE_K�L ?%y (�%SVCPRG�1ho8��e���o�m3��o�o�`4 �`5�(-�`6PU�`7@x}�`���l9��{�d:?��a�o� �a�oE��a�om��a ���aB���aj叟a ���a�5��a�]� �a����a3����a[� ՟�a�����a��%��a ӏM��a��u��a#��� �aK�ů�as���a�� mob�`�o�`8�}�w� ������ɿ���ؿ� ��5�G�2�k�VϏ�z� �Ϟ����������1� �U�@�y�dߝ߯ߚ� �߾�������?�*� Q�u�`������� �����;�&�_�J� ��n������������sj_DEV ~y	�MC:���_OUT�",REC� 1�Z� d �   	�    ��@�� ����A�����
 �PS?D#6 r��UO� �� �� `��� �Z�{� �r� *�  +X�- � I- �- !
- � �X�YZ��PSJ;4 ��?  (� E � ��R ���� E- �� �/e/�l!4�/��� X� (,/>/P/�/�/*�""4� =�!� � ؀  ?"S1h��'!�/���("- ��\?�?$=�= �?�?�?"OOFO4OjO |O^O�O�O�O�O�O�O �O_ __T_B_x_f_ �_�_�_�_�_�_�_o ooPo>oto�oho�o �o�o�o�o�o(
 L:\�p���w,����4� "�X�F�|���p����� ֏ď����0��@� f�T���x�����ҟ� Ɵ���,��<�b�P� ��h�z������ί� �(�:��^�L�n�p� ������ܿ�п� � 6�$�Z�H�jϐ�rϴ� �����������2�D� &�h�Vߌ�z߰ߞ��� ��������
�@�.�d��R��ZjV 1��w P����j� 
�� ��<��
TYPEV�FZN_CFG ;��5d��4�GRP 1��A�c ,B� A�� D;� B����  B4�RB21HE�LL:�(
��?x���<%RS'! ��H3lW� {������`2Vh������%w�����#!�1�����7�2�0d�����HK 1��� �k/f/x/�/�/�/ �/�/�/�/??C?>?�P?b?�?�?�?�?��OMM ����?���FTOV_ENB� ���+�HOW_R�EG_UIO��I_MWAITB�.JKOUT;F��LIwTIM;E���O�VAL[OMC_UN�ITC�F+�MON�_ALIAS ?�e�9 ( he ��_&_8_J_\_B_ �_�_�_�_j_�_�_o o+o�_Ooaoso�o�o Bo�o�o�o�o�o' 9K]n��� �t���#�5�� Y�k�}�����L�ŏ׏ ������1�C�U�g� ���������ӟ~��� 	��-�?��c�u��� ����V�ϯ����� �;�M�_�q������ ��˿ݿ����%�7� I���m�ϑϣϵ�`� ������ߺ�3�E�W� i�{�&ߟ߱������� ����/�A�S���w� ����X������� ���=�O�a�s���0� ������������' 9K]���� b���#�G Yk}�:��� ���/1/C/U/ / f/�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_O
O�O�O�O �O�OvO�O__%_7_��C�$SMON_�DEFPRO ����`Q� *SY�STEM*  d�=OURECAL�L ?}`Y (� �}6copy� frs:ord�erfil.da�t virt:\�temp\=>1�92.168.4��P46:8188� 12>_�_�_l}.�V*.d�_�^�_�`oro�oe
xyz�rate 61 �+o=oOo�o�oe �g�o�a�o�ocu��b9�_�Xmpback�oRr���l]0�rmdb(`*��� �b�t���c4x�t:\)���;�SqpU����
� }5��a�����W׏h�z�� ��:�Տ���
�� ��A�ӟd�v�����.� ;�я��������� O�`�r�������2�͟ ޿���'�¿K�\� nπϓ���8�ɯ���� ���#���G��j�|� �o�g+�=�O������|)2244 �� ��c�u���5�6� �������"Ͻ�5��� b�t����Ϭ߾�:�U� ����
߮������� hz��1CU�0�
�E�52Tp� �cu����5�6 ����"��5��b/t/�/c�_�_B�1660 W/�/�/�/ o�/�)�/`?r?�?� �o;?M?�?�?O' �4�?�?cOuO�O�� 5/�'�O�O�O/"/�O �(�Ob_t_�_���� KTV_�_�_o�_�_ >@�_hozoo�O�O:_ �_�o�o
_�oA_�o dv��_.o;�_� ��o��Oo`�r� ���o�o2�oޏ��� 'K\�n�������$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1����?���%֟ ��&�	��\�?�f� ��u��������ϯ�� "��F�)�;�|�_��� ����ֿ��˿��� B�%�f�I�[Ϝ�Ϧ� �ϵ�������,��6� b�E߆�i�{߼ߟ��� ��������L�/�V� ��e��������� ���6��+�l�O�v� �������������� 2V9K�o� ������& R5vYk��� ��/��<//F/ r/U/�/y/�/�/�/�/ ?�/&?	??\???f? �?u?�?�?�?�?�?�? "OOFO)O;O|O_O�O �O�O�O�O�O_�O_ B_%_f_I_[_�__�_ �_�_�_�_�_,oo6o boEo�oio{o�o�o�o �o�o�oL/V �e������ ��6��+�l�O�v��������PARAM� ����� ��	��P�����OFT_K�B_CFG  �⃱���PIN_S_IM  ����C�U�g�����RVQSTP_DSB,��򂣟����SR ��/�� & � AR�����T�OP_ON_ER�ސ���PT�N /�@��A	�RINGo_PRM� ���VDT_GRP �1�ˉ�  	 ������������Я� ����*�Q�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߣߠ߲� ����������0�B� i�f�x�������� �����/�,�>�P�b� t��������������� (:L^p� ������  $6HZ�~�� �����/ /G/ D/V/h/z/�/�/�/�/ �/�/?
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8___\_��VP�RG_COUNT���@���REN�BU��UM�S��__�UPD 1�/�8  
s_�oo *oSoNo`oro�o�o�o �o�o�o�o+&8 Jsn����� ����"�K�F�X� j���������ۏ֏� ��#��0�B�k�f�x� ��������ҟ����� �C�>�P�b������� ��ӯί�����UYSDEBUG�P��P�)�d�YH�SP�_PASS�UB�?Z�LOG �V�U�S)�#��0�  ��Q)�
�MC:\��6���_MPC���U���Q�ñ8� �Q�SA/V �����ǲ�%�ηSV;�T�EM_TIME �1��[ (�P"��T!y�ؿT1SV�GUNS�P�U'��U���ASK_OPTION�P�U�Q��Q��BCCFGg ��[u� n�X�G�`a�gZo��� �ߕ��߹������� :�%�^�p�[���� ������ �����6�!� Z�E�~�i���������%�������&8�� nY�}�?�� ԫ ��(L :p^����� ��/ /6/$/F/l/ Z/�/~/�/�/�/�/�/ �/�/2?8 F?X?v? �?�??�?�?�?�?�? O*O<O
O`ONO�OrO �O�O�O�O�O_�O&_ _J_8_n_\_~_�_�_ �_�_�_�_o�_ o"o 4ojoXo�oD?�o�o�o �o�oxo.TB x��j���� ����,�b�P��� t�����Ώ��ޏ�� (��L�:�p�^����� ��ʟ��o��6� H�Z�؟~�l������� د���ʯ ��D�2� h�V�x�z���¿��� Կ
���.��>�d�R� ��vϬϚ��Ͼ����� ��*��N��f�xߖ� �ߺ�8��������� 8�J�\�*��n��� ���������"��F� 4�j�X���|������� ������0@B T�x�d���� �>,Ntb ������/� (//8/:/L/�/p/�/ �/�/�/�/�/�/$?? H?6?l?Z?�?~?�?�? �?�?�?O�&O8OVO hOzO�?�O�O�O�O�O �O
__�O@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<o^o�oro �o�o�o�o�o�o  J8n$O��� ��X���4�"��X�B�v��$TBC�SG_GRP 2��B�� � �v� 
 ?�  ������׏ �������1��U�g��z���ƈ�d,� ���?v�	 H�C��d�>�����e�CL  B�p��Пܘ������\)��Y  A��ܟ$�B�g�B�Bl�i�X�ɼ���X��  D	J���r�����C����үܬ	���D�@v�=�W�j� }�H�Z���ſ���������v�	�V3.00��	�m61c�	*`X�P�u�g�p�>���2v�(:�� ��p���  O�����p�����z�JCFG� �B��� ,���������=��=�c�q�K� qߗ߂߻ߦ������ ��'��$�]�H��l� ������������#� �G�2�k�V���z��� �����������p *<N���l�� �����#5G Y}h���� v�b��>�// /V/ D/z/h/�/�/�/�/�/ �/�/?
?@?.?d?R? t?v?�?�?�?�?�?O �?*OO:O`ONO�OrO �O�O��O�O�O_&_ _J_8_n_\_�_�_�_ �_�_�_�_�_�_oFo 4ojo|o�o�oZo�o�o �o�o�o�oB0f T�x����� ��,��P�>�`�b� t�����Ώ������ �&�L��Od�v���2� ����ȟʟܟ� �6� $�Z�l�~���N����� دƯ�� �2��B� h�V���z�����Կ¿ ����.��R�@�v� dϚψϪ��Ͼ����� ��<�*�L�N�`ߖ� �ߺߨ����ߚ��� ����\�J��n��� ��������"���2� X�F�|�j��������� ������.TB xf������ �>,bP� t�����/� (//8/:/L/�/�ߚ/ �/�/h/�/�/�/$?? H?6?l?Z?�?�?�?�? �?�?�?O�?ODOVO hO"O4O�O�O�O�O�O �O
_�O_@_._d_R_ �_v_�_�_�_�_�_o �_*ooNo<oro`o�o �o�o�o�o�o�o& �/>P�/��� ������4�F� X��(���|�����֏ ����Ə0��@�B� T���x�����ҟ���� ��,��P�>�t�b� ������������� �:�(�^�L�n����� ��2d�����̿� $�Z�H�~�lϢϐ��� �����Ϻ� ��0�2� D�zߌߞ߰�j����� �����
�,�.�@�v� d����������� ��<�*�`�N���r� ������������& J\�t��B ������F 4j|��^��p��/�  2 �6# 6&J/6"��$TBJOP_G�RP 2����  ?i�X,i#�p,� ��x�J� �6$�  �_< �� �6$� @2 �"	 ߐC�� �&b � Cق'�!�!>�c��
559>�0�+1�33=�{CL� fff?+0?�ffB� J1�%�Y?d7�.��/>��2\)?0�5����;��hC=Y� �  @� �!?B�  A�P?�?��3EC�  Dp�!�,�0*BOߦ?��3JB��
:���Bl�0��0�$�1��?O6!Aə�A�ДC�1D�G6��=q�E6O0�p���B�Q�;��A�� ٙ�@L3D	�@�@__�O�O>B�\JU�OHH��1ts�A@333@?1� C�� �@�_�_&_8_>��D��UV_0�LP�Q30<'{�zR� @�0�V �P!o3o�_<oRifoPo ^o�o�o�oRo�o�o�o �oM(�ol�pP~��p4�6&�q�5	V3.00��#m61c�$�*(��$1!6�A� �Eo�E���E��E��F��F!��F8��FT��Fqe\F�N�aF���F�^�lF���F�:�
F�)F���3G�G���G��G,I�R�CH`�C��dTDU�?D���D��DE(�!/E\�E���E�h�E��ME��sF�`F+'\FD���F`=F}�'�F��F��[
F���F���M;S@;Q�*�|8�`rz@/&�
8�6&<��1�w��^$ESTPARS�  *({ _#HR���ABLE 1̒p+Z�6#|�Q� (� 1�|�|�|�5'T=!|�	|�
|�|�T˕6!|�|�|����RDI��z!�ʟܟ� ��$���O ������¯ԯ�����	S��x# V���˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �U-����ĜP�9�K� ]�o��-�?�Q�c�u����6�NUM  V�z!� > � Ȑ����_CFGG �����!@b �IMEBF_TT�����x#��a�VER腣b�w�a�R 1=�p+
 (3�6"	1 ��  6!���� ������ �9�$�:�H� Z�l�~����������� ����^$��_���@x�
b MI_CWHANm� x� k�DBGLV;0o��x�a!n ETHER_AD ?�� �y�$"�\&n oROUT��!p*�!*�SNM�ASK�x#�255.h�fx^$�OOLOFS_D�I��[ՠ	ORQCTRL �p+ ;/���/+/=/O/ a/s/�/�/�/�/�/���/�/�/!?��PE_�DETAI��P�ON_SVOFF��33P_MON ��H�v�2-9ST�RTCHK ����42VTCOMPATa8�24:0�FPROG %�%CA)&O�3?ISPLAY��L:_INST_MPe GL7YDUS���?�2LCK�LPKQ?UICKMEt �O��2SCRE�@>�
tps��2 �A�@�I��@_Y����9�	SR_GRP� 1�� ���\�l_zZg_�_ �_�_�_�_�^�^�o j�Q'ODo/ohoSe� �oo�o�o�o�o�o�o !WE{i�������	1?234567���!���X�E1�V[
� �}ipnl�/a�gen.htmno��������ȏ~��Panel _setup̌}�?���0�B�T�f�  ��񏞟��ԟ��� o����@�R�d�v��� ���#�Я����� *���ϯůr������� ��̿C��g��&�8� J�\�n�����϶��� ������uϣϙ�F�X� j�|ߎߠ����;��߀����0�B��*NU�ALRMb@G ?�� [���� �������� ��%�C��I�z�m�������v�S�EV  �����t�ECFG �Ձ=]/BaA$ �  B�/D
  ��/C�Wi{�� ����� PRց; �To\�o�I�6?K0(% ����0����� //;/&/L/q/\/�/0�/�/l�D �Q��/I_�@HIST� 1ׁ9  �(  ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1?pv?�?�?�?�� >?P=962c?�?
OO0.O�?�?�136�?|O �O�O�OAOSOeO�O_ _0_�HM___q_�_�_ �_�_H_�_�_oo%o 7o�_[omoo�o�o�o Do�o�o�o!3E ��a81�ou�� ����o���)� ;�M��q��������� ˏZ�l���%�7�I� [���������ǟٟ h����!�3�E�W�� ��������ïկ�v� ��/�A�S�e�Pb ������ѿ������ +�=�O�a�s�ϗϩ� ��������ߒ�'�9� K�]�o߁�ߥ߷��� �����ߎ�#�5�G�Y� k�}���������� �����1�C�U�g�y� ��v�����������	 �?Qcu�� (����) �M_q���6 ���//%/�I/ [/m//�/�/�/D/�/ �/�/?!?3?�/W?i? {?�?�?�?�����?�? OO/OAOD?eOwO�O �O�O�ONO`O�O__ +_=_O_�Os_�_�_�_ �_�_\_�_oo'o9o Ko�_�_�o�o�o�o�o �ojo�o#5GY �o}������?���$UI_PA�NEDATA 1�������  	�}��0�B�T�f�x��� )����mt�ۏ��� �#�5���Y�@�}��� v�����ן��������1��U�g�N������ �1��Ïȯگ ����"�u�F���X� |�������Ŀֿ=��� ���0�T�;�x�_� �Ϯϕ��Ϲ������,ߟ�M��j�o߁� �ߥ߷������`�� #�5�G�Y�k��ߏ�� ������������� C�*�g�y�`������� ��F�X�	-?Q c����߫��� �~;"_F ��|����� /�7/I/0/m/���� �/�/�/�/�/�/P/!? 3?�W?i?{?�?�?�? ?�?�?�?O�?/OO SOeOLO�OpO�O�O�O �O�O_z/�/J?O_a_ s_�_�_�_�O�_@?�_ oo'o9oKo�_oo�o ho�o�o�o�o�o�o�o #
GY@}d� �&_8_����1� C��g��_�������� ӏ���^���?�&� c�u�\�������ϟ�� �ڟ�)��M��� ��������˯ݯ0�� ���7�I�[�m���� ������ٿ�ҿ��� 3�E�,�i�Pύϟφ�`�Ϫ���Z�l�}���@1�C�U�g�yߋ�)� ��#������� ��$� 6��Z�A�~�e�w�� ����������2���V�h�O�����v�p���$UI_PANELINK 1�v��  ��  ��}1�234567890����	-?G  ���o����� a��#5G�	�����p&���  R�����Z ��$/6/H/Z/l/~/ /�/�/�/�/�/�/�/ 
?2?D?V?h?z??$? �?�?�?�?�?
O�?.O @OROdOvO�O O�O�O �O�O�O_�O�O<_N_``_r_�_�_�0,�� �_�X�_�_�_ o2oo VohoKo�ooo�o�o�o �o�o�o��,> r}�������� ����/�A�S�e� w��������я��� tv�z����=�O� a�s�������0S��ӟ ���	��-���Q�c� u�������:�ϯ�� ��)���M�_�q��� ������H�ݿ��� %�7�ƿ[�m�ϑϣ� ��D��������!�3� Eߴ_i�{�
�߂��� �߸������/��S� e�H���~��R~'� '�a��:�L�^�p� ��������������  ��6HZl~� ��#�5���  2D��hz��� ��c�
//./@/ R/�v/�/�/�/�/�/ _/�/??*?<?N?`? �/�?�?�?�?�?�?m? OO&O8OJO\O�?�O �O�O�O�O�O�O[�_ ��4_F_)_j_|___�_ �_�_�_�_�_o�_0o oTofo��o��o� �o�o�o,>1 bt����K� ���(�:���� {O������ʏ܏�uO �$�6�H�Z�l����� ����Ɵ؟����� � 2�D�V�h�z�	����� ¯ԯ������.�@� R�d�v��������п ���ϕ�*�<�N�`� rτ��O�Ϻ�Io���� �����8�J�-�n߀� cߤ߇����߽���� o1�oX��o|��� �����������0� B�T�f���������� ����S�e�w�,>P bt��'��� ��:L^p ��#���� / /$/�H/Z/l/~/�/ �/1/�/�/�/�/? ? �/D?V?h?z?�?�?�? ??�?�?�?
OO.O�� ROdO�߈OkO�O�O�O �O�O�O_�O<_N_1_ r_�_g_�_7OM��m�$UI_QU�ICKMEN  }��_�AobRESTOR�E 1�  �|��Rto�o�im�o�o�o �o�o:L^p �%������o ����Z�l�~��� ��E�Ə؏���� � ÏD�V�h�z���7��� ����/���
��.�@� �d�v�������O�Я �����ßͯ7�I� ��m�������̿޿�� ��&�8�J��nπ� �Ϥ϶�a�������Y� "�4�F�X�j�ߎߠ� �������ߋ���0�xB�T�gSCRE`�?#mu1�sco`u2��3���4��5��6��7��8��bUSER�q�v��Tp���ksT����4��5��6���7��8��`NDO_CFG �#k�  n` `PD�ATE ����NonebS�EUFRAME � �TA�n�RTOL_ABRTy��l��ENB����G�RP 1�ci/a?Cz  A�����Q�� $6HRd��`U�����?MSK  ������Nv�%�U�%����bVISCA�ND_MAX��I��FAILO_IMG� �PݗP�#��IMREG�NUM�
,[S�IZ�n`�A��,VONTMOU4��@���2���a��a�����FR:\� � M�C:\�\LOGn�B@F� !��'/!+/O/�Uz �MCV�8#7UD1r&EX{+�S��PPO64_t��0'fn6PO��LIb�*r�#V���,f@�'޻/� =	�(SZ�V�.����'WA�I�/STAT ����P@/�?�?��:$�?�?��2D�WP  ��P� G@+b=���� H�O_JMP�ERR 1�#k
�  �2345678901dF�ψO {O�O�O�O�O�O_�O *__N_A_S_�_
� MLOWc>
 �g_TI�=�'�MPHASE  ���F��PSH�IFT�1 9�]@<�\�Do�U#o Io�oYoko�o�o�o�o �o�o�o6lC U�y������ ��	�V�-�e2�����	VSFT1��2	VM�� S�5�1G� ���%�A�  B8̀�̀�@ pكӁ˂�у��z�ME@�?�q{��!c>&%�a�M1��k�0�{ ��$`0TDINEND��\�O� �z�����S��w��P�{��ϜRELE�Q��Y���\�_AC�TIV��:�R�A ��e���e�:��RD� ���YBO�X �9�د�6���02����190.0.�8�3��254t��QF�	 ��X�j��1�r�obot���   p�૿�5pc��̿������7�����-�f�ZA+BC�����,]@U� �2ʿ�eϢωϛϭ� ������ ���V�=� z�a�s߰�E�Z��1�Ѧ