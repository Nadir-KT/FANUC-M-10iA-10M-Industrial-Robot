��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 � �1�K(�|UREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8GW�+0�$Y $DB\� 6COMW!2�MO� H.	 �\rVE�1$F8�RA{$O�UD�cB]CTMP1_FtE2}G1_�3�B�2�GXD�#
� d $CARD_EXIST4�$FSSB_T�YP!AHKBD�_SNB�1AGN G�n $SLO�T_NUM�AP�REV4DEBU�� g1� ;1_EDI}T1 � 1�G=� S�0%�$EP�$O�P�U0LEToE_OK�BUS�oP_CR�A$;4xAV� 0LACIw�1�R�@k �1$@M{EN�@$D�V��Q`PvVA{G B�L� OU&R ,�A�0�!� B� L�M_O�
eR�"C�AM_;1 x�r$ATTR84�@� ANNN@5�IMG_HEIG�H�AXcWIDTH�4VT� �UU0F�_ASPEC�A;$M�0EXP�.@�AX�f�CF�D X $GR� �� S�!.@B�PNF�LI�`�d� UIR�E 3T!GITCH�+C�`N� S�d_LdZ`AC�"�`EDp*�dL� J�4S�0� �<za�!p;G0� � 
$WARNM�0f�!�@� -s�pNST� CORyN�"a1FLTR{u�TRAT� T}p  $ACCa1�p��|{�rORIضP�C�kRT0_S�~B\qHG,I1� [ T�`�"3I��pTYD�@*2 �3`#@� �!�B*HEDDcJ* Cd�2_�U3_�4_�5_�6_��7_�8_�94�ACO�$ <� �o�op�hK3 1#`O_Mc@�AC t � E�#6NGPvABA � �c1�Q8��`,��@Bnr1�� d�P�0Xe���axnpUP@&Pb26���p�"J�pS_R�rPBC��J�rĘߜJV�@U� B��`s}�g1�"YtP_*0wOFS&R @� �RO_K8T��aIT<�3T�NOM_�0�1�p�3� >��D !�� Ќ@��hPV��mCEX�p� �0g0ۤ<�p�r
$TF�2Co$MD3i�TO�3��0U� F� R��Hw2tC1(�Ez�g0#E{"F�"F�F40CP@�a2 �@$�PPU�3N�)ύRևAXd�!DU��AI�3�BUF�F=�@1c |pp���pPIT�� PP�M�M��y��F�SIMQSI�"ܢVAڤT�:��Px T�`(z�M��P�B�qFAC5Tb�@EW�P1��BTv?�MC�k �$*1JB`p�*1DEC��F���y=�� �H0�CHNS_EMP�1�$G��8��@_�4�3�p|@P��3�TCc�(r/�0-sx���ܐ� MBi��!����J�R� i�SEGFRR��Iv �aR�Tp9N�C��PVF4>�>bx &��f {uJc!�Ja��� !28�pץ�AJ���SIZ�3S�c�B�TM���g��>JaRSINFȑb� ��q�۽�н�����L�3�B���CRC�e�3CCp���� c��mcҞb�1J�cѿ��.����D$ICb�C q�5r�ե��@v�'���SEV���zF��_�եF,pN��ܫ�p?�4�0A�! �r ���h�Ϩ��p�2��@�a�� �د� �	�>�Cx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�IM�]pUR��QUA1w  $@TITO1�/S@S�!����"0�?DBPXWO��B0=!5�$SK���2M@DBq�!"�"v�PR�� 
� 8=����!# S q1�$2�$z���LB�)$�/���� %�/��$C�!&?�$ENE�q.'*?�Ú �RE�p2(H ���O�0#$L|3$$�#�B[�;�К�FO_D��ROSr�#������3�RIGGER�6P�ApS����ETUR�N�2�cMR_8�T�Uw��0EWM��M�GN�P���B#LAH�<E���P��O&$P� �'P@D�Q3�CkD{��DQฑ�4�11��FGO_oAWAY�BMO��t�Q#!� CS_�o)  �PIS�  I gb {s�C��A��[ �B$�S��AbP�@�EW-�TNTVճ�BV�Q[C�(c`�UWr�P�J��P�$0���SAFE���V_S}V�bEXCLU�:�nONL2��S1Y�*a&�OT�a'�HI_V�4��B���_ *P0� 9�9_z��p ��A;SG�� +nrr� @6Acc*b��G�#@E��V.iHb?fANNU�N$0.$fdID�U�2�SC@�`�i�a��j�f/�!�pOGI:$2,O�$FibW$�}�OT9@�1 ?$DUMMYT��d�a��dn�� � �E-o ` ͑HE4�(sg�*b�SAB��SU�FFIW��@CUA=�c5�g6r�!MSW�E. 8�Q�KEYI5���T�M�10s�qA�vIN����ї!��/ Dބ�HOST_P! �rT��ta��tn��tsp��pEMӰV��� S�BLc ULI�0 � 8	=ȳ�r��DTk0�!1 � �$S��ESAMPL��j�۰f璱f����I�0��[ $SUB�k�#0�C��T�r#a�SAVʅ��c��`�C��P�fP$n0yE�w YN_B#72 0Q�DI{dlp�O(��9#$�R�_I�� �EN�C2_S� 3 ! 5�C߰�f�-  �SpU����!4�"g��޲�1T���5@X�j`ȷg��0�0K�4x�AaŔAVER�q8ĕ9g�DSP�v��PC��r"��(����ƓVALUߗHE4�ԕM+�IPճ���OPP ��TH��֤��P�S� �۰	F��df�J� ����C1+6 H>�bLL_DUs�~a�3@{��3:���OT�X"���so��0NO�AUTO�!7�p!$)�$�*��c4�(��C� 8�C, ���&�L�� 8H *8�LH <6� ���c"�`, `Ĭ�k� ��q��q��sq��~q���7��8��9��0T����1��1̺1ٺU1�1�1 �1ʕ1�2(�2����2�̺2ٺ2�2�2� �2�2�3(�3R��3��̺3ٺ3�U3�3 �3�3�=4(�C(���?��!9 <�9�&�z���I��1���M��QFqE@'@� : ,6���Q? �@P?Q9��5�9�E�@�A��a�A� ;p�$TP�$VA�RI:�Z���UP2f�P< ���TDe� ��K`Q�����wBAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�H  ���P���@`�!>�t ;E��sC�ST�D� D���c�<� 	C��{� �_���l���R  �����FORCEUP�?b��FLUS�`H��N>�F ���RD_CM�@E������ p��@vMP��REMr F�Q��1k@���7�Q
K4	NJ�5EF1Fۓ:�@IN2Q��sOVO�OVA�	�TROV���DT<Հ�DTMX�  ��@�
ے_PH",p��CL��_TpEȓ@�pK	_(�Y_T���v(��@A;QD� ������!0tLܑ0RQ���_�ad����M�7�CL�d�ρRIV'�{��E�ARۑIOHPCȸ@����B�B��CM�9@���R �GC3LF�e!DYk(Ml�ap#5TuDG��p�� �%��FSSD �s? P�a�!�1��E�P_�!�(�!1���E�3�!3�+5�&��GRA��7�@��4;�PW��ONn��EBUG_SD2H�P�{�_E A �L����T�ERM`5Bi5�p��ORI#e0Ci5w?��SM_�P��Ze0D�9TA�9E�6� �UP\�Fg� -�A{�AdP|w3S@B$SEG�:v� EL{UUSE�@NFIJ�B$�;1x젎4�4C$UFlP=�$,�|QR@��_G90Tk�D�~SwNST�PAT��<��APTHJ��E�p%B`�'EC����AR$P�I�aS�HFTy�A�A�H_�SHORР꣦6 ��0$�7PE��E�O#VR=��aPI�@��U�b �QAYLOW���IE"�r�A��?���ERV��XQ� Y��mG>@�BN��U�\��R2!P.uAScYMH�.uAWJ0G�ѡEq�A�Y�R�Ud>@��EC���EaP;�uP;�6WOR>@�M`�0SMT6�G3�GR��13�a�PAL@���`�q�uH� � ���T�OCA�`P	P�`$OP����p�ѡ��`0O��RE�`R4C�AO�p낎Be�`R�Eu�h�A���e$PWR�IMu�RR_�cN��q.=B I&2H���p�_ADDR��H_LENG�B�q�q�q�$�R��S�JڢSS��SKN��u\��u̳�uٳSE�A�jrmS��MN�!K������b����OL�X��p����`ACRO3pJ�@��X�+�p�Q��6�OUP3��b_�IX��a�a1 ��}򚃳���(��H ��D��ٰ��氋�+IO2S�D���x��	�7�L $d�<�`Y!_OFFr��PRM_��ɡH�TTP_+�H:�M; (|pOBJ]"�p���$��LE~C|d���N � ��.֑AB_�Tqᶔ�S�`H�LVh�K�R"uHITCOmU��BG�LO�q���h�����`���`SS� ���HW��#A:�Oڠ<`I�NCPU2VISIOW�͑��n��to���to�ٲ �IOL]N��P 8��R��^p$SLob oPUT_n�$p¾�P& ¢��Y F_�AS�"Q��$L ������Q  U�0	P�4A��50��ZPHY`��-��x��UOI �#R `�K��� �$�u�"pPp�k���$������UeJ5�S-���NE6W�JOGKG̲DISĖ��Kp���#T �(�uAVF�+`�CTyR�C
�FLAG2v�LG�dU ����؜�13LG_SIZ����b�4�a��a�FDl�I`�w� m� _�{0a�^��cg���4� ����Ǝ���{0��� �SCH_���a�SLN�d�VW���AE�"����4��UM��Aљ`LJ�@�DAUf�EAU�p��d|�r��GH�b6�OGB�OO��WL ?�6 IT��y0�wREC��SCR �ܓ�D
�\���MARGm�!��զ ��dH%�����S����W���U� �JGM[�M�NCHJ���FNK�EY\�K��PRGƂ�UF��7P��FW�D��HL��STP���V��=@��А�RES��HO`����C9T@��b ��7�[�UL����6�(RD� ����Gt��@PO��������MD�FOCU��RwGEX��TUI��	I��4�@�L� ����P����`���P��NE��CANAx��Bj�VAILI��CL !�UDCS_CHII4��s�O�D(!�S���S���/��_BUFF��!X�?PTHA$m���v`����a�!Y�?P��j�\3��`OS1Z2Z�3Z��_�� Z � ��[aEȤ��.ȤIDX�dPSRraO���zA�STL��R}�Y&�� Y$E�C���K��&&��п![ L Q��+00�	P���`#q�dt
�U�dw<���_ \ ?�4Г�\���Ѩ#\0C4�] ���CLDPL��UTRQLI��dڰ�)�$FLG&�� 1�#b�D���'B�LD�%�$�%ORGڰ5�2 �PVŇVY8�s�T�r�$}d^ ���$6��$
�%S�`T� �B0�4}�6RCLMC�4`]?o?�9세�MI�p�}d_ d=њRQz��DSTB�pƽ ;F�HHAX��R JHdLEXC#ESr��BM!p�a`��/B�T8B�j�`a�p=F_A7J�i��KbOtH� K�db� \Q���v$MB�C�LI|�)SREQUIR�R�a.\o�AXODEBUZ�ALt M��c�b�{P����2ANDRѧ`�`ad;�2�ȺSDC��N�INl�K�x`��XB� N&��aZ���UwPST� ezr7LOC�RIrp�EX<fA�p�9AA�ODAQ��f XfY�OND�rMF,� �Łf�s"��}%�e/�� �8FX3@IGG>�� g ��t"���ܓs#N�s$R�a%��iL��hL�v�@��DATA#?pE��%�tR��Y�Nh t $MD`qI}�)nv� ytq�yt�HP`�Pxu��(�zsANSW)�yt@��yu�D+�)\b���0o�i[ �@CUw�V�p� 0XeRR2��j �Du�{Q��7Bd$C'ALIA@��G���2��RIN��"�<NE�NTE��Ck�r`^�آXb]���_N�q�lk���9�D���Bmn��DIVFDH�@t���qnI$V,���S�$��$Z �X�o�*�����oH �$BE�LT�u!ACCE�L�.�~�=�IR!C�� ���D�T�8�O$PS�@�"LD��r��#^�S�Eы T�PATH3���I�"��3x�p�A_W���ڐ���2nC��4�_{MG�$DD��<T���$FW�Rp`9��I�4��DE7��PPABN��ROTSPEE�[g�� J��[�C@4�D�?$USE_+�VPi��SYY���1- qYN!@A�Ǧ�OFF�qǡMOUf��NG���OL����INC�tMa6���HB��0HBENCS�+�8q9Bp�4�FDm�IN�IԒ]��B���VE��#�y�23_�UP񕋳LOWL����p� B���D�u�9B#P`�x ���BC<v�r�MOSI��B�MOU��@�7PERoCH  ȳOV�� â
ǝ����D��ScF�@MP����� Vݡ�@y�j�LUk��Gj�p�UP=ó���Ķ�TRK��AYLOA�Qe��A��Ԓ��p��N`�F�RTI�A$��MOUІ�HB�B S0�p7D5���ë��Z�DUM2ԓS�_BCKLSH_CԒk����ϣ����=���ޡ �	ACLAL"q��1м@�էCHK� �S�RTY��^�%E1Qq9_�޴_UM�@�9C#��SCL0�r��LMT_J1_LD��9@H�qU�EO��p�b�_�e�k�e�SP�C��u���N�PC��N�Hz \P��C��0~"XT��CN�_:�N9��I�SF!�?�V���U�/����ԒT���CB!�SH �:��E�E1T�T��`��y���T��PA �&�_P��_� =�@�����!����J6 1L�@��OG�G��TORQU��ON ֹ��E�R��H�E�g_W2���_郅����I�I�I��Ff`xJ�1�~1�VC3�0BD:B��1�@SBJR�KF9�0DBL�_SM��2M�P_sDL2GRV�`���fH_��8d���COS���LNH��� �����!*,�a1Z���fMY�_(��TH��)THE{T0��NK23��ت"��CB�&CB�CAA�B�"��!�!�&SB� 2�%GTS�Ar�CIMa������,4#97#$DU���H\1� �:B�k62�:AQ(rSf$N	E�D�`I��B+5��$̀�!A�%�5�78���LPH�E�2���2SC%C%@�2-&FC0JM&̀V�8QV�8߀LVJV!KUV/KV=KVKKVYKVgIH�8FRM��T#X!KH/KH=KHKKUHYKHgIO�<O�8�O�YNOJO!KO�/KO=KOKKOYKOM&F�2�!+i%0d�7�SPBALANC�E_o![cLE0H_�%SPc� &�b&|�b&PFULC�h`�b�g�b%p�1k%��UTO_��T13T2�i/�2N��"� {�t#�Ѱ`�0�*��.�T��OÀ<�v I�NSEG"�ͱREqV4vͰl�DIF��f��1lzw��1m���OBpq�я?�MI�{���nLCHWA�RY�_�AB��!�$MECH�!o �,�q�AX��P���8�7Ђ�`n 
�d�(�U�ROB��CR�ԒH���8(�M�SK_f`�p P+ �`_��R/�k�z�����1S�~�|�z��{���z��qINUq��MTCOM_C|� �q  ����pO�$NORE�n����pЂr �8p GRe�uSD��0AB�$XY�Z_DA�1a���D�EBUUq������su z`$��COD��G L���p��$BUFIND�X|�  <�MO�Rm�t $فU A��֐���Ԑ<���rG��u � ?$SIMUL  S��*�Y�̑a�OBJE|�`̖ADJUSꘞݐAY_IS�Dp�3����_FI�=��Tu 7�~�6� '��p} =�C�}p�@bŝD��FRIr��T&��RO@ \�E}'�=y�OPWOYq��v0Y�SYSByU/@v�$SOPġ�d���ϪUΫ}pPR�UN����PA��Dp���rɡL�_OUo�顢q�$)�I�MAG��w��0Pf_qIM��L�INv��K�RGOVRDt��X�(�P*�J�|��0L_�`]��0�SRB1�0��M�񦷺ED}��p ��N��PMֲ�୐�w�S�L�`q�w x �$OVSL4vSDI��DEX��Đ�#���-�V} *�N 4�\#�B�2�G�B�_�M�x� �q�E� x Hw��p�ЯATUSW���Cp�0o�s���BTM��*��I�k�4��x�\԰q�y Dw�E&���@E�r��7����З�EXE��ἱ������f q�z @�w���UP'��$�pQ�XN������ļ��� �PG΅{� h $SUB�����0_���!�M/PWAIv�P7ãՓLOR���F\p˕�$RCVFAILs_C���BWD΁|�v�DEFSP!p | Lw����p��\���UNI+������H�R�+�}_�L\pP��y�P��p�}H�> �*�j��(�s`~�N�`KET�B�%�J�PE Ѓ~z��J0SIZE	 ���X�'���S�OR~��FORMAT�``��c ��WrEM�t���%�UX��G�%�c�PLI��p� � $ˀP_S�WI�p{��J_P�L��AL_ ������A��B��� C���D�$E���.�C_�U�� ?� � ����*�J3K0����TI�A4��5��6��MOM��������ˀB��AD������l����PU� NR������)H��m���� A$PI �6q��	����� K4�)6�U��w`��_SPEEDgPG� �������Ի�4T��� � @��SAMr`��\�]��MOV_�_$�npt5���5���1���2���������'�S�Hp�IN�'�@� +����4($4+T+�GAMMWf�1'��$GET`�p���D�a���

pLIBRt>�II2�$HI=�!_g�t��2�&E;��(1A�.� �&LW�-6 <�)56�&]��v�p���V��$PD#CK���q��_?�����q�&���7����4���9+� ��$IM_SR�pD`�s�rF��r�rLE��¹Om0H]��0��-�pq��PJqUR_SCRN�FA����S_SAVE_�D��dE@�NOa�C AA�b�d@�$q�Z�I ǡs	�I� �J�K� �� ��H�L��>�"hq ������ɢ��� bW^US�A�,M4���a��)q`��3��WW�I@v�_�q�.M�UAo�� � $sPY+�$W�P�vNG�{��P:��R`A��RH��RO�PL��@���q� ��s'�X;�	OI�&�Zxe ���m�G� p��ˀ�3s��O�O�O�O�O�aa�_т� |��q�d@�� .v��.v��d@��[wFvr��E���% -�r;B�w�|�tPn���PMA�QUa ��Q8��1�wQTH�HOLG�oQHYS��ES�F�qUE�pZB��Oτ�  ـPܐ(�AP����v�!�t�O`�q��u�"���FA��IGROG�����Q2����o�"��p��INFOҁ�׃V����R��G3�I��� (�0SLEQ�������Y���O���Á�D�P0Ow0���!�E0NU��AUyT�A�COPY�P=�/�'��@Mg�N���=�}1������ ��RiG��Á���X_�P��$;ख�`��W��P��@�������EXT_CYC b!HᝡRpÁ�r��7_NAe!А����ROv`	�� � ���PORp_�1�E2�SRV ��)_�I�DI��T_ �k�}�'���dЇ������5��6��7��8�i�H�SdB���2��$��F�p��GPL8eAdA
�TAR�Б@ ���P����n�d� ,�0FL`L�o@YN��K�M��=Ck��PWR+�9�z����DELA}��dY�pAD�a� ��QSKIP4�� �A�$�OB`NT2�} ��P_$�M� ƷF@\bIpݷ�ݷ� ݷd����빸��Š��Ҡ�ߠ�9���J2R� ��� 46V�EX� TQQ�� ��TQ������ ��`����RDC�V� �`��X)�R�p������r��m$RGEA�R_� IOBT�2FcLG��fipER��DTC���Ԍ���2T�H2NS}� 1����G T\0 ����u�M\Ѫ`I��d��REF�1�Á� l�h��ENsAB��cTPE�0 4�]����Y�]��ъQ n#��*��"�������2�Қ�߼���������3�қ'�9�K�]�o�� ����4�Ҝ�����������
�5�ҝ!�3�E�W�(i�{��6�Ҟ��������������7�ҟ�-?Qcu�8�Ҡ������^�SMSKÁ�l���a��EkA��MO[TE6�����@0�݂TQ�IO}5�QISTP�QR�W@��� �pJ�����p����E�"$DSB_SIGN�1�UQ�x�C\�TP��S�232���R�iDEVICEUS�|XRSRPARIT���4!OPBIT�Q�I�OWCONTR`+�TQ��?SRCU� �MpSUXTASK�3N�p�0p$TATU�P�PH �0������p_XPC)��$FREEFRO�MS	pna�GET\�0��UPD�A�2ΙqRSP� :���� !$US�AN�na&����ER1I�0�RpRYq5*"�_j@�Pm1�!�6WRK9KD���6��~QFRIEND�Q��RUFg�҃�0TO�OL�6MY�t$�LENGTH_VT\�FIR�pC�@�ˀE> +IUFINt-RM��RGI�1�ÐAITI�$GX�ñ3IvFG2v7G1`���p3�B�GPR�p�1F�O_n 0��!�RE��p�53҅U�T�C��3A�A�F �G((��":���e1n!���J�8�%���%]�� �%�� 74�XS O0�L��T�3�H&��8���%b453G�E�W�0�WsR�TD ����T��M����Q�T�]�$V 2�����1�а91�8�02*�;2k3�;3�:i fa�9-i�aQ��NS���ZR$V��2BVwEVP�	V�B;�����& �S�`��F�"�k�@�2�a�PS�E��$pr1C��_$Aܠ�6wPR��7vMU�cS��t '�/89�� 0�G�aV`��p�d`����50�@��-�
25S^�� ��aRW�����B�&�N�A)X�!�A:@LAh�^�rTHIC�1I�8��X�d1TFEj��q>�uIF_CH�3�qaI܇7�Q�pG1Rx�V���]��:�u�_�JF~�PRԀƱ��RVAT��� ���`���0RҦ�DO�fE��COUԱ��A�XI���OFFS=E׆TRIGNS����c����h�����Hx�Y��IGMA0�PA�pJ�E�ORG�_UNEV�J� ��S�����d ӎ$CА�J�GR3OU����TOށ�!DSP��JOG�Ӑ�#��_Pӱ�"O��q����@�&KEPF�IR��ܔ�@M}R&��AP�Q^�Eh0��K�SYS�q"K�;PG2�BRK�B��߄�pY�=�d�����`AD������BS�OC���N��DU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR-���C��ˢΓ�OR٧3N]0ڦF��ڦ��OV��SF��p���F+�r!���CC��1q"LCHD}L��RECOVʤc0��Wq@M������#RO�#��Ȑ_+���� @0�e@VER��$OFSe@CV/ �2WD�}���Z2���TR�!|���E_FDO��MB_CM���B��BL�bܒ#��adt�VQR�$0p���G$�7�AM5��� e����_M;��"'����8$CA��'�E�>8�8$HBK(1���IO<�����QPPA������
���������DVC_DBhC;��#"<Ѝ�r!"S�1[ڤ�S�3[֪�/ATIOq 1q� �ʡU�3���CAB Ő�2�CvP��9P^�B��_� �SUBCPU�ƐS�P � M�)0NS�cM�"r�?$HW_C��U���S@��SA�A�pl$�UNITm�l_�A�T���e�ƐCYC=Lq�NECA����FLTR_2_F�IO�7(��)&B�LPxқ/�.�_SCT�CF_`�Fb�l���|��FS(!E�e�CHA��1��4�D°"3�RS�D��$"}����_Tb�PRO����� KEMi_��a�8!�a !�a��D�IR0�RAILAiCI�)RMr�LO��C���Qq��#q��V��PR=�S�A�p�C/�� 	��FUsNCq�0rRINP`�Q�0��2�!RAC �B ��[���[gWARn���BL�A�q�A����D�Ak�\���LD@0���Q��qeq�TI"r��K�hPgRIA�!r"AF��Pz!=�;��?,`�R�K���MǀI�!�D�F_@B�%1n�LM��FAq@HRDY4�4_�P@RS�A�0|� �MULSE@x���a ���ưt��m�$�1-$�1$1o������ x*�EaGE ����!AR���Ӧ�09�2,%� 7�wAXE��ROB���WpA��_l-��SY�[�W!‎&S�'WR�U�/-1��@�STRП�����Eb� !	�%��J��AB� ����&9�����OTo0v 	$��ARY�s�#2��Ԓ�	ёFI�@��$LINK(|�qC1�a_�#����%kqj2XYZ@��t;rq�3�C1j2J^8'0B��'�40����+ �3FI���7`�q����'��_Jˑp���O3�QOP_�$2;5���ATBA�2QBC��&�DUβ�&=6��TURN߁"r��E11:�p��9GFL��`_���* �@�5�*7���Ʊ 1�� KŐM��&8���"r��ORQ��a �(@#p=�j�g�#qXUp�����mTOVEtQ:�M��i���U��U��VW�Z�A�Wb��T {�, ��@;�uQ���P \�i��UuQ�We�eL�SERʑe	��!E� O���UdAas���4S�/7����AX��B�'q��E1�e ��i��irp�jJ@�j �@�j�@�jP�j@ �j �!�f��i��i��i ��i��i�y�y��'y�7yTqHyDEBU8�$32����qͲf2G + AB�����رnSVS�7� 
#�d��L�#�L� �1W��1W�JAW��AW� �AW�QW�@!E@?\D2�3LAB�29U�4�Aӏ��C  �o�ERf�5� �� $�@_ A��!�PO��à�0#��
�_MRAt�� �d � T��ٔEcRR����;TY&����I��V�0�cz�TOQ�d�PL[ �d�"��� ?�w�! �� pp`T)0���_�V1Vr�aӔ����2Bٛ2�E����@�H�E���$W�����5V!��$�P��o�cI��aΣ	 HELL_CFG!ߵ 5��B_7BASq�SR3��.� a#Sb����1�%��2��3���4��5��6��72��8���RO�����I0�0NL�\CAB8+�����ACK4������,�\@2@�&�?�_�PU�CO. U�OUG�P~ ����m�������TPհ_KA1R�[@_�RE*��qP���|�QUE����uP����CSTOPI_AL7�l�k0���h��]�l0SEM��4�(�M4�6�TYfN�SO���DIZ��~�A�����m_TM>�MANRQ��k0�E����$KEY?SWITCH����m���HE��BEAiT��|�E- LE~�����U��F!Ĳ���B�O_HOM=OnGREFUPPR&P��y!� [�C��O��-ECOC��Ԯ0_�IOCMWD
�a��	�m��� � DHh1���UX���M�xβgPgCFORC��n� ��OM.  � @�5(�U�#P, 1��, �3��45��NPXw_ASt�� 0���ADD���$S�IZ��$VAR\���TIP/�.�
�A�ҹM�ǐ��/�H1�+ U"S�U!Cz����FRIF��J�S0���5Ԓ�NF�� ܍� � xp`SIƗ�TE�C���CSG%L��TQ2�@&���x�� ��STMT��2,�P �&BWuP���SHOW4���S�V�$�� �Q�A00�@Ma}����� �����&���5���6��7��8��9��A��O ���Ѕ�Ӂ���0��F��� G�� 0G���0G���@GP��PG��1	1	U1	1+	18	1E	U2��2��2��2��U2��2��2��2��U2��2��2	2	U2	2+	28	2E	U3��3��3��3��U3��3��3��3��U3��3��3	3	U3	3+	38	3E	U4�4��4��4��U4��4��4��4��U4��4��4	4	U4	4+	48	4E	U5�5��5��5��U5��5��5��5��U5��5��5	5	U5	5+	58	5E	U6�6��6��6��U6��6��6��6��U6��6��6	6	U6	6+	68	6E	U7�7��7��7��U7��7��7��7��U7��7��7	7	U7	7+	78	7E�	�VP��UPD>s�  �`Nм��5�YSLOt�� � L��d���A�aTA�0d��|��ALU:ed�~�CU�ѰjgF!aID_L��ÑeHI�jI��$FILE_���d���$2�fSA>��� hO��`E_BL�CK��b$��hD_CPUyM�yA��c�o�db����R ��Đ
PW��!� -oqLA��S=�ts�q~tRUN�qst �q~t���qst�q~tw �T��ACCs��X -$�qLEN;��tH��ph��_�I��ǀLOW_7AXI�F1�q�d2*�MZ���ă��W��Im�ւ�aR�TOR���pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v��������TCV��؁��T ��ي�����t�V��$��V�Jj�R�MA����J��m�u�b����q2j�#�U�{�t�K�JK��VK;���H����3��J0����J�J��JJ��AAL���ڐ��ڐԖ4Օ5���N1���ʋƀJW�LP�_(�g��м�pr�� `�`GGROUw`��B�ПNFLIC��f�R�EQUIRE3�E�BU��qB���w�2�����p���q5�p��� \��APPRҒ�C}�Y�
ްEN�٨CLO7��S_!M��H���u�
�qu�o� �`�MC��8���9�_MG��C��Co��`M�в�N�B;RKL�NOL|�N�:[�R��_LINђ�$|�=�J����Pܔ�� ���������������Q6ɵ�̲8k�D�>���� ��
���q)��7�PATH3�L�B�L��H�w�ڡ��J�CN�CA��Ғ�ڢB�IN�rU�CV�4a��C!�UMB��Y,���aE�p�����ʴ���PAYwLOA��J2L`OR_AN�q�Lpp����$�M�R_F�2LSHR��N�L�Oԡ�Rׯ�`ׯ�ACRL_G�ŒЛ�� ��Hj`߂$H�M���FLEXܣ��qJ�u� : �������������1�F1�V�j�@�R�d�v�������E ����ȏڏ����"� 4�q���6�M���~�� U�g�y�ယT��o�X��H������藕? �����ǟِݕ�ԕ@����%�7��JJ�� � V�h�z����`AT�採@�EML�� S��J|��Ŝ�JEy�CTR,��~�TN��FQ��HAND_VB-�q��v`�� $���F2M����ebSW���q'��� $$MF�:�Rg�(x� ,4�%��0&A�`�=��aM)F�AW�Z`i�Aw�A��X X�'pi�UDw�D��Pf�G�p��)STk��!x��!N��DY�pנM�9$`% Ц�H��H�c�׎���0� ��Pѵڵ㵀����������� ���1��R�6���QASYMvř����v��J���cі�_SH>��ǺĤ�ED� ���������J�İ�%��C�IDِ�_VI�!X�2PV_UCNIX�FThP�J�� _R�5_Rc�cTz�pT�V ��@���İ�߷��U �����
(�T2��Hqpˢ��a3EN�3�DI�����O4d�`J�� x g"IJAAȱz�aa bp�coc�`a�pdq�a�� ��OMMEB��� �b�RqAT(`PT�@� S��a7�;�AȠ�@�h�a�iT�@�<� $DUM�MY9Q�$PS�_��RFC��$v �p���Pa�� XƠ���ST�E���SBRY�M�21_VF�8$S/V_ERF�O��Ls�dsCLRJtA��O�db`O�p �� D $GLOBj�_LO���u�q��cAp�r�@aSYS��qADR``�`T�CH  � ,x��ɩb�W_NA��c�7��SR��?�l ��� 
*?�&Q�0"?�;'?� I)?�Y)��X���h��� x������)��Ռ�Ӷ� ;��Ív�?��O�O�O|�D�XSCRE�j�p����ST�F�s}y`�����/_HA�q� TơgpTYP�b����G�aG���Od0IS_䓀e�;UEMd� ����p�pS�qaRSM_��q*eUNEXCE1P)fW�`S_}pMрx���g�z�����ӑC�OU��S�Ԕ 1-�!�UE&��Ubwr���PROGM�F�L@$CUgpP�O�Q��5�I_�`H>� � 8�� �_HE�PS�#��`?RY ?�qp�b���dp�OUS>�� � @6p�v�$BUTTp�R|pR�COLUMq�<e��SERV5��PANEH�q� w� �@GEU��Fy��)$HE�LPõ)BETERv�)ෆ���A  � ��0��0��0�ҰIN簪c�@N(��IH�1��_�o ֪�LN�r'� �qpձ_ò=��$H��TEX8l����FLA@��/RELV��D`���������M��?,@�ű�m����"�USRVIEW�q�� <6p�`U�`��NFI@;�FOsCU��;�PRI� �m�`�QY�TRI}P�qm�UN<`�Md� #@p�*eW�ARN)e6�SRT+OL%��g��ᴰ�ONCORN��RA�U����T���w�V�IN�Le� =$גPATH9�ג�CACH��LOG�!�LIMKR���x�v���HOST��!�b�R��OgBOT�d�IM>�	 �� ���Zq��Zq;�VCPU_�AVAIL�!�EX	�!AN���q�`�1r��1r��1 ��\��p�  #`C�����@$TOOLz�$��_JMP�� ���e$S�S����SHIF��Nc�P�`ג��E�ȐR����OSU�R��Wk`RADILѮ��_�a��:�9a���`a�r��LULQ�$OUTPUT_3BM����IM�ABp �@�rTIL'SCO��C7� ������&��3 ��A���q���m�I�2G��1V�pLe��}��yDJU��N_�WAIT֖�}Ҵ�{�%! NE�u��YBO�� ��� $`�t�S�B@TPE��NE�Cp�J^FY�nB_T��R�І�a$�H[YĭcB��dM� ��F� �p�$�pb��OP?�MAS�_�DO�!QT�pD���ˑ#%��p!"DE�LAY�:`7"JO Y�@(�nCE$��3@` �xm��d�pY_[�!"g�"��[���P?� �1ZABC~%��  $�"�R��
ϐ�$$C�LAS����i��!ϐϐ � �VIRT]��/ 0A�BS����1 5�� < �!F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ8i{0-�AXL�pl��!�63  �{tIqN��qztPRE�����v�p�uLAR�MRECOV �9�rwtNG�� �.;	 A  � �.�0PPLIMC��?5�p��Handl�ingTool �o� 
V7.5�0P/23-�  o�PB��
��w_SWt� UP�!7� x�F0��t��A� v� �864�� �it��y� N�" 7DA5��� j� QB�@ϐo�None�isͅ˰ ���T�]�!LAAWx>�_l�V�utT��s9�UTO�"�Њt�y��HGAPCON
0g�1��Uh�oD 1581����̟ޟry����/Q 1���p �,�蘦���;�@���q_��"�" g�c�.�H����D�HTTHKYX��"�-�?�Q��� ɯۯ5����#�A�G� Y�k�}�������ſ׿ 1�����=�C�U�g� yϋϝϯ�����-��� 	��9�?�Q�c�u߇� �߽߫���)����� 5�;�M�_�q���� ����%�����1�7� I�[�m���������� !����-3EW i{����� �)/ASew ����/��/ %/+/=/O/a/s/�/�/ �/�/?�/�/?!?'? 9?K?]?o?�?�?�?�? O�?�?�?O#O]����TO�E�W�DO_CLEAN�����C�NM  � �__/_A_S_�DSPDRYR�O&��HIc��M@�O�_ �_�_�_oo+o=oOo aoso�o�o���pB��v# �u���aX�t�������9�PLUGGp���G��U�PRCvPB�@��_�or�Or_��SEGF}�K[mwxq�O�O������?rqLAP�_�~q�[�m���� ����Ǐُ����!�|3�x�TOTAL�f| yx�USENU�p��� �H���B��R�G_STRING� 1u�
�kMn�S5�
ȑ�_ITEM1Җ  n5�� ��$�6� H�Z�l�~�������Ư�د���� �2�D��I/O SIG�NAL̕Tr�yout Mod�eӕInp��S�imulated�בOut���OVERR�P =� 100֒In� cycl��ב�Prog Abo�r��ב��Sta�tusՓ	Hea�rtbeatїMH Faul��Aler'�W�E� W�i�{ύϟϱ������� �CΛ�A�� ��8�J�\�n߀ߒߤ� �����������"�4��F�X�j�|���WOR {pΛ��(ߎ����� � �$�6�H�Z�l�~��� ������������ 2PƠ�X �� A{������ �/ASew������SDEV[�o�#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g?>y?PALTݠ1 ��z?�?�?�?�?O"O 4OFOXOjO|O�O�O�O��O�O�O�O_�?GRI�`ΛDQ�?_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o�o2_l�R��a\_�o "4FXj|� ���������0�B�T��oPREG �>�� f���Ə؏� ��� �2�D�V�h�z� ������ԟ���Z���$ARG_��D ?	���;���  �	$Z�	[�O�]O��Z�p�.�S�BN_CONFIOG ;��������CII_SA_VE  Z������.�TCELLSETUP ;��%HOME_I�OZ�Z�%MOVq_��
�REP�l�U�(�UTOBAC�Kܠ���FRA:\z� �\�z�Ǡ'`�pz���ǡi�INI�0�z���n�MESSAG���ǡC�>��ODE_D����ą�%�O�4�n�PA�USX!�;� ((O>��Ϟˈ� �Ϭ���������� *�`�N߄�rߨ߶�g�~l TSK  w�x��_�q�UPDT+���d!�A�WSM�_CF��;����'�-�GRP 2�:�?� N�BŰA|��%�XSCRD1�;1
7� �ĥĢ����������*� ������r��������� ��7���[�&8J�\n��*�t�GR�OUN�UϩUP�_NA�:�	�t��_ED�1�7�
 �%-B?CKEDT-�2��'K�`���-(t�z�q�q�z���2t1�����q�k�(/��ED3/��/�.pa/�/;/M/ED4�/ t/)?�/.?p?�/�/ED5`??�?<?.p�?O�?�?ED6O �?qO�?.MO�O'O9OED7�O`O_�O.p�O\_�O�OED8L_,�_�^-�_ oo_�_ED9�_�_]o��_	-9o�oo%oCR_ 9]�oF�o�k� � NO_D�EL��GE_U�NUSE��LA�L_OUT �����WD_AB�ORﰨ~��pIT_R_RTN��|ONONSk����˥CAM_PAR�AM 1;�!�
� 8
SONY� XC-56 2�34567890� ਡ@����?��( С�\�
���{����^�HR5q�̹��ŏ�R57ڏ�Af�f��KOWA �SC310M
��x�̆�d @ <�
���e�^��П \����*�<��`��r�g�CE_RIA�_I�!�=�Ff��}�z� ���_LIU�]������<��FB�GP� 1��Ǯ��M�_�q�0�C* Y ����C1��9���@��G���CR�CU]��d��l��s��QR�����[Դm���v���������W C����(���숁=�HE�`ONF�Iǰ�B�G_PR/I 1�{V�� �ߖϨϺ�����������CHKPAUS��� 1K� , !uD�V�@�z�dߞ߈� ���߾������.��R�<�b���O���������_MOR��� �6��� 	 �����*�� N�<�������?Ғ�q?;�;����K���9�P���ça�-:���	�

��M���pU�ðț�<��,~��DB��튒)
mc�:cpmidbgX�f�:����u��	p�/���H�
� �s>�܌�Q�?��g�/��f�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����o=L���*MC��1����?43���1��t�īCz�  BHH�>'��B�$�9G��<5@@�C���1Y
K�@��D��;A�e�8��.D�� ��1�=B��IE��Ce=�D�<�?X�F���1Y	X���'w�1����s���.�p���b���BDw�M@x8��K�CҨ����g@D��p@�0E��8EX��EQ�EJ�P F�E�F�� G��=F�^F E�� F�B� H,- Ge��H3Y��:��  >�33 ����~  n48�~@��5Y�E>��ðA��Y<#�
�"Q ���+_�'R_SMOFS�p�.�8��)T1��DE ���
Q��;�(P  B_<_���R����	op6C4RP�Y
s@ ]AQ��2s@C�0B3�MaCR�@*cw��UT�p�FPROG %�z�o�oigI�q���v���ldKEY_TB�L  �&S�#� ��	
�� �!"#$%&'(�)*+,-./0�1i�:;<=>?�@ABC� GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇�������������������s���p`LCK�lx4�p`�`STAT ���S_AUTO_D�O���5�IND�T_ENB!���R��Q?�1�T2}�^�S�TOPb���TRL^r`LETE��Ċ�_SCREEN ��Zkcs�c��U��MMEN�U 1 �Y  <�l�oR�Y1� [���v�m���̟���� �ٟ�8��!�G��� W�i��������ïկ ��4���j�A�S��� w�����迿�ѿ��� �T�+�=�cϜ�sυ� �ϩϻ�������P� '�9߆�]�o߼ߓߥ� �������:��#�p� G�Y��������� ��$����3�l�C�U� ��y����������� ���	VY)�_MA�NUAL��t�DB;CO[�RIGڇ
��DBNUM� ���B1 e
�PXWO_RK 1!�[�_�U/4FX�_�AWAY�i�G�CP  b=�Pj_CAL� #�j�Y���܅ `�_�  1">�[ , 
�m�g�&/~&lMZ�I�dPx@P@#ONT�IMه� d��`&�
�e�MOT�NEND�o�RECORD 1(�[qg2�/{�O��! �/ky"?4?F?X?�( `?�?�/�??�?�?�? �?�?)O�?MO�?qO�O �O�OBO�O:O�O^O_ %_7_I_�Om_�O�_ _ �_�_�_�_Z_o~_3o �_Woio{o�o�_�o o �oDo�o/�oS �oL�o����@ ���+�yV,�c� u��������Ϗ>�P� ����;�&���q��� 򏧟��P�ȟ�^�� ����I�[����� � ��$�6�������j�TOLERENC�wB���L���� CS_CFG �)�/'dM�C:\U�L%04�d.CSV�� cl��/#A ��CH��z� //.ɿ��(�S�RC_OUT �*��1/V�S�GN +��"���#�27-JA�N-20 21:�540j�48+? P;��ɞ��/.��f�pa�m��PJPѲ���VERSION� Y�V2�.0.�ƲEFLOGIC 1,�/ 	:ޠ=��ޠL��PROG_�ENB��"p�UL�Sk' ����_WRSTJNK ��"�fEMO_OPT?_SL ?	�#�
 	R575/#=�����0�B�|���TO  ��صϗ��V_F EX�d�%��PAT�H AY�A\p�����5+ICT�-Fu-�j�#�egS�,�STBF_TTS�(@�	d���l#!w�� �MAU��z�^"MS%WX�.�<�4,#�
Y�/�
!J�6�%ZI~m��$SBL_FAUL(�y0�9'TDIA[��1<�<� ����1234567G890
��P�� HZl~���� ���/ /2/D/V/hh/�� P� ѩ�yƽ/��6�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?�,�/�UMP���� �ATR���1OC@�PMEl�OOY_T�EMP?�È�3pF���G�|DUNI���.�YN_BRK �2_�/�EMGDI_STA��]��E�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�a�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��aDzr�A W�_BWD�p��xf�́t�_DI�� 9�5�d�T�asRֆSTEP��:P��OP_DOv��f�PFACTOR_Y_TUNwdM��EATURE �:�5̀rQ�Handling�Tool �� \�sfmEng�lish Dictionary���roduAA� Vis�� Ma�ster����
�EN̐nalog� I/O����g.�fd̐uto S�oftware �Update  �F OR�mat�ic Backu�p��H596�,�ground �Editޒ  1� H5Cam�era�F��OP;LGX�ell𜩐�II) X�omm�Րshw���com揭co���\tp����pane�� � opl��tyl�e select^��al C��nJ�~Ցonitor��gRDE��tr��?Reliab𠧒�6U�Diagno�s(�푥�552�8�u��heck �Safety U�IF��Enhan�ced Rob �Serv%�q )� "S�r�UserG Fr[�����a���xt. DIO 6�fiG� sŢ��wendx�Err�MLF� pȐĳr�r�� ����  !���FCTN Men�u`�v-�ݡ���T�P Inېfac��  ER J�GC�pבk E�xct�g��H55�8��igh-Sp�ex�Ski1�  �2
P��?���m�munic'�on1s��&�l�ur�ې���ST Ǡ��c�onn��2��TX�PL��ncr�s�tru����"FA�TKAREL Cmd. LE�{uaG�545\�ſRun-Ti��E{nv��d
!����ؠ++�s)�S/�W��[�Lic�enseZ��� 4�T�0�ogBook�(Syڐm)��H�54O�MACRO�s,\�/Offs�e��Loa�MH�������r, k�M�echStop �Prot���� l�ic/�MiвSh�if����ɒMixpx��)���xSPS��Mode Swiwtch�� R5W��Mo�:�.�� 7#4 ���g��K��2h�ulti-T�=�M���LN (�Pos�Reg�iڑ������d�ݐtO Fun�ǩ�.�����Num~����Ï lne��ᝰ Adjup������  - W��ta�tuw᧒T��RDMz�ot��s�cove U�9����3Ѓ�uesOt 492�*�o������62;�SNP�X b ���8 Jy7`���Libr��FJ�48���ӗ� ����
�6O�� Pa�rts in VCCMt�32���x	�{Ѥ�J990��{/I� 2 P���TMILIB��Ht���P�AccD��L�
TE$TX܍ۨ�ap1S�Te<����pkey���wգ�d��Un�exceptx�motnZ��������3є�� O��΄� 90J�єSP CSXC<�f�l�Ҟ� Py�We}�Β�PRI�>vr\�t�men�� ��/iPɰa������vGrid�play��v��0�)��H1�M-10iA(B201 ��2\� 0\k/�A/scii�l�Т��ɐ/�Col��ԑG7uar� 
�� /�P-�ޠ"K��stN{Pat ��!S��Cyc�҂�or�ie��IF8�ata- quҐ�� ƶ���mH574��RML��am���Pb�HMI De3�(�b����PCϺ�P�asswo+!��"PE? Sp$�[���stp��� ven���Tw�N�p�YEL?LOW BOE	k$wArc��vis���3*�n0WeldW�cial�7�V#Mt�Op����1y�֠ 2F�a�pocrtN�(�p�T1�`T� �� ��xy]ֹ&TX��tw�ig�j�1� b� ct\��JPN ARC?PSU PR��ovݲOL� Sup�2fil� &PAɰא�cro�� "PM�(����O$SS� enвtex�� r����=�t�ssag$T��P��P@�Ȱ�锱�rtW��H'�>r�dpn��n1#
t�!� z ���ascbin4p�syn��+Aj�M� HEL�NCL� VIS PKG�S PLOA`�McB �,�4VW��RIPE GET_VAR FIEo 3\t��FL[��OOL: ADD� R729.FD/ \j8'�CsQ�Q�E��DVvQ�sQNO WTWTE��>}PD  �^��b�iRFOR ��EC�Tn�`��ALSE� ALAfPCPM�O-130  M�" #h�D: H�ANG FROM�mP�AQfr��R7�09 DRAM �AVAILCHE�CKSO!��sQVP�CS SU�@LIMCHK Q +P~d�FF POS��F��Q R593�8-12 CHA�RY�0�PROGR�A W�SAVE�N`AME�P.SV2��7��$En*��p�?FU�{�TRC|� �SHADV0UPD�AT KCJўRS�TATI�`�P M�UCH y�1��I�MQ MOTN-�003��}�ROB�OGUIDE DAUGH�a���*�Gtou����I� Š�hd�ATH�PepM�OVET�ǔVM�XPACK MA�Y ASSERT��D��YCLfqTA��rBE COR �vr*Q3rAN�pR�C OPTION�SJ1vr̐PSH�-171Z@x�tcǠSU1�1Hp^9R!�Q�`_T�P��'��j�d{tby app wa 5IҌ~d�PHI���p�aT�EL�MXSPD' TB5bLu 1��U�B6@�qENJ`CEV2�61��p��s	�may n�0� �R6{�R� �Rtr�aff)�� 40�*�p��fr��sy�svar scr� J7��cj`DJ�U��bH V��Q/��PSET ERR�`J` 68��PN�DANT SCR�EEN UNRE�A��'�J`D�pPA��pR`IO 1����PFI�pB�pG/ROUN�PD��G���R�P�QnRSVIP� !p�a�PDIGI?T VERS�r}B�Lo�UEWϕ P�06  �!��MA�Gp�abZV�DIx�`� SSUE��ܰ�EPLAN {JOT` DEL�p�ݡ#Z�@D͐CAsLLOb�Q ph���R�QIPND��I{MG�R719���MNT/�PES ��pVL�c��Holp�0Cq���tPG:�`:C�M�canΠ���pg.v�S: 3�D mK�view� d�` �p��eat7У�b� of �P�y���ANNOT �ACCESS M���Ɓ*�t4s a��lok��Fle�x/:�Rw!mo?�PA?�-�����`~n�pa SNBPJ AUTO-�0�6f����TB��PIA�BLE1q 636>��PLN: RG$��pl;pNWFMD�B�VI���tWIT� 9x�0@o��Qu�i#0�ҺPN RR�S?pUSB�� t� & removb�@ )�_��&AxEP7FT_=� 7<`�p�P:�OS-14;4 ��h s�g���@OST� � C�RASH DU �9��$P�pW�� .$��LOGI�N��8&�J��6b0�46 issue� 6 Jg��: �Slow �st~��c (Hos`��c���`IL`IMP�RWtSPOT:Wqh:0�T�STYW =./�VMGR�h��T0CAT��hosB��E�q��� �uO�S:+pRTU' �k�-S� ����E:���pv@�2�� t\�hߐ��m ��al�l��0�  $�H� �WA͐��3 CN�T0 T�� Wr}oU�alarm���0s�d � �0SE1����r R{�OMEpBp���K� 55��REàSEst��g�     �KoANJI�no����INISITA�LIZ-p�dn1we�ρ<��dr�� l�x`�SCII L��fails w��� ��`�YSTE�a���o��Pv� IItH���1W�Gro>P�m ol\wpSh�@�P��Ϡn cfslxL@АWRI ЏOF Lq��p?�F��up��de-r�ela�d "A�Po SY�ch�Ab�etwe:0INDc t0$gbDO����r� `�Gig�E�#operab[ilf  PAbHi�xH`��c�lead�\etf�Ps�r��OS 030�&: f{ig��GLA )P� ��i��7Np t�pswx�B��If��g������5aE>�a EXCE#dU��_�tPCLOS��"�rob�NTdpF�aU�c�!���PNIO V750�Q�1��Qa��DB Ė�P M�+P�QED��DET��-� \�rk��ONLINEhSBUGIQ ߔXĠi`Z�IB�S a�pABC JAR�KYFq� ���0MSIL�`� R�pNД� �p0GAR��D�*pR��P�"! jK�0cT�P�Hl#n��a�ZE V�� TwASK�$VP2(��4`
�!�$�P�`WI[BPK05�!FȐ�B/��BUSY oRUNN�� "��ȁ����R-p�LO��N�DIVY�CU9L��fsfoaBW�p���30	�V��ˠIT`�a5�05.�@OF�UGNEX�P1b�af�@��E��SVEMGN� NMLq� D0pCC_SAFEX �0c�08"qD �PE�T�`N@�#J87�����RsP�A'�M��K�`K�H G�UNCHG۔MEKCH�pMc� T� � y, g@�$ ORY LEAKA8�;�ޢSPEm�Ja:��V�tGRIܱ��@�CTLN�T�Rk�FpepR�j506�EN-`IN������p �`�Ǒk!��Tq3/dqo�STO�0)A�#�L�p �0�@�Q�АY�&�;pb1CTO8pP�s���FB�0@Yp`�`DU��a!O�supk�t4 � PЙF� Bnf�Q�PSVGN-1��V�S'RSR)J�UP��a2�Q�#D�q l �O��QBRKCTR5Ұ�|"-�r�<p�c�j!INVP�D ZO� ��T`h#�Q�cHset,|D��"DUAL� w�2*B�RVO117 A�]�TNѫt�+bTa2�473��q.?��sA�Uz�i�B�comp�lete��604�.� -�`haknc�U� F�Нe8��  ��npJ�tPd!q��`��� 5Nh596p�!5d��� "p�P�P�Q�0�P2@�p�A� xP��R(}\*xPe� aʰI����E��1��p� j � � xSP�^P ��A�AxP�q 5 siug��a��"AC;a���
�bCexPb_p��.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o`�dxP�b]o2�� �c�b�c�ixP�jupf�rm�dxP�o�`ex�e�a�oFdxPtpe�d}o��u`�cptlcibxzxP�lcr�xrxP\�blsazEdxP_fm�}gcxP�x@���o|sp�o�mc(�N�ob_jzop�uD6�wf��t��wms�1q��sld�)��jCmc�o\�n��nuhЌ���|st�e��>�p1l�qp�iwck����uvf0uߒ��lv�isn�Cgacu�lwQ
E F  ;! Fc.fd�Qv��� qw���Dat�a Acquis�i��nF�|1�RR6�31`��TR�QDM�CM �2�P75�H�1�P583xP1���71��59`�5�P57<PxP�Q����¨�(���Q��o p�xP!daq\�o�A��@�� ge/�e�tdms�"DMEsR"؟,�pgdD����.�m���-��qacq.<᡾xPmo��Dh���f{�u�`13���MACROs, Sksaff�@z�����03�SR�Q(��Q6���1�Q9ӡ�R�ZSxh��PxPJ643�@�7ؠ6�P�@�PRS��@���e �Q�UС �PIK�Q52 P�TLC�W��xP3 (��p/O��!�P�n �xP5��03�\sfmnmc "MNMCq�<��Qj��\$AcX�FM�� �ci,Ҥ�X����cd�pq+�
�sk�SKx�xP�SH560�,P��,�y�refp "REFp�d�A��jxP	�of�OF�c�<gy�to�TO�_����ٺ����+je�u��caxi�s2�xPE�\�e�q"�ISDTc��]�porax ��MN�x�u�b�isde܃�h�\�w�xP! is_basic��B�� P]��QAxes��R6������.�(sBa�Q�ess� �xP���2�D�@�z�atis���(�{������~��m��F�Mc�u�{�
ѩ�MNIS��ݝ����x�����ٺ��x� j7}5��Devic��� Interfa�c�RȔQJ7540��� xP�Ne`� �xP�ϐ2�б�����dn� "DNE����
tpdnu�i5UI��ݝ	b�d�bP�q_rs�ofOb
dv_aro��u����>�stchkc���z	 �(}onl��G!ffL+H�@J(��"l"/�n�bx��z�hamp���T�C�!i�a"�59`��S�q��0 (�+�P�o�u�!2��xpc�_2pcchm��C�HMP_�|8бpe�vws��2쳌pc�sF��#C SenxPacro�U·�-�R6�Pd�xPk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GE�M,\i(��Dgesnd�5���H{�}Ha��@sy���c�Isu�xD��Fmd��I��7��4���u���AccuCal�P�4� ��Rɢ7ޠB0��6+56f�6��99\aFF q�S(�U��2�
X�ap�!Bd��cb_��SaUL��  ��� ?�ܖto��ot�plus\tsr�nغ�qb�Wp��t����1��Tool (N. A.)�[K�7�Z�(P�m�����bfcls� k94�"K4p��qt�pap� "PS�9H�stpswo`��p�L7��t\�q ����D�yt5�4�q��@w�q��� �M�uk��rkey����s���}t�sfeatu�6�EA��� cf)t\�Xq�����d�h5���LRC0�md�!�C587���aR�(�����2V��8c?u3l\�pa3}H�&r-��Xu���t,�� �q "�q�Ot��~,���{@�/��1c�}����y�p �r��5���S�XAg��-�y���Wj874��- iRVis<���Queu�� �Ƒ�-�6�1���(����u���tӑ�����
�tpvtsn? "VTSN�3C�t+�� v\pRDV����*�prdq\�Q<�&�vstk=P�������nm&_�դ��clrqν���get�TX��Bd����aoQϿ�0qstr�D[� ��t�p'Z��Ɵ�npv��@�enlIP0��D!x�'�|����sc ߸��tv�o/��2�q���v b����q���!���h�]��(� Con�trol�PRAuX�P5��556�A�@59�P56.@5�6@5A�J69�$@982 J55?2 IDVR7�hq A���16�H���La��� ��Xe�f�rlparm.fn�FRL�am��C9�@(F������w6{���A��QJ6�43�� 50�0L�SE
_pVAR� $SGSYSC���RS_UNIT�S �P�2�4tA�T�X.$VNUM_OLD 5�1�xP�{�50+�"�` Funct���5tA�� }��`#@�`3�a0��cڂ��9���@HA5נ� �P���(�A ����۶}����ֻ}��bPRb�߶~p{pr4�TPSPI0�3�}�r�10�#;A � t�
`���1���96�����%C�� A�ف��J�bIncr �	����\���1o�5qni4�MNINp	xP�`���!���Hour  �� 2�21� �AAVM����0 ��T�UP ��J5�45 ��616�2�VCAM � (�CLI{O ��R6�<N2�MSC "�P �STY�L�C�28~ 13�\�NRE "FwHRM SCH^��DCSU%O�RSR {b�04� �EIOC��1 j 542 �� os| � eg�ist�����7��1�MASmK�934"7 ���OCO ��"3�8��2���� C0 HB��� 4�";39N� Re�� ��LCHK
%OP�LG%��3"%MH�CR.%MC  ; 4l? ��6 dPI�s54�s� DSW%�MD� pQ�K!63!7�0�0p"�1�Р"�4 �6<27 CgTN K � 5 ��%�"7��<25�%/�=T�%FRDM� ��Sg!��930 FB( NBA�P� ( �HLB  Men��SM$@jB( PV3C ��20v��2�HTC�CT�MIL��\@PAC� 16U�hAJ`SA�I \@ELN��<29�s�UECK <�b�@FRM �b�sOR���IPL��}Rk0CSXC ���VVFnaTg@H�TTP �!26� ��G�@ob�IGUI"%IPG�S�r� H863 �qb�!�07r�!34 |�r�84 \so`0! Qx`CC3 Fb�291�!96 rb!g51 ���!53R%� 1!s3!��~�.rp"9js VATFU�J775"��pLR6�^RP�WSMjUCTO�@xT58 F!s80���1XY ta�3!770 ��8�85�UOL  GTS�o
�{` LCM ��r| TSS�EfP6� W�\@CPE �`��0VR� l�QN�L"��@001 i7mrb�c3 =�b0�0���0�`6 w�b^-P- R-�b8n@75EW�b9 �Ґa�� ���b�`ׁ�b2 O2000��`3��`4*5�`5!�c��#$�`7.%�`8 h�605? U0�@B�6E"aRp7� !Pr8 t�a@�tr�2 iB/�1vp3L�vp5 Ȃtr9Σʐa4@-p�r3 	F��r5&�re`u�&�r7 ��r8�U�p9 \h738�a��R2D7"�1�f��2&�7� �3� 7iC��4>w58Ip�Or60 C�L��1bEN�4 I�py�L�uP��@N�-PJ8d�N�8NeN�9 H�(r`�E�b7]�|�⠂8�Вࠂ9 2H��a`0�qЂ5�%?U097 0��@q1�0���1 (�q�3 5R���0 ���mpU��0�0��7*�H@(q�\P"wRB6�q124�b`;��@���@06� 6x�3 pB/x�u ���x�6 H606�a1� ��7 6� ���p�b15�5 ����7jUU1g62 �3 g���4*�65 2ec "_��P�4U1`����B1���`0'�1�74 �q��P�E1�86 R ��P�7� ��P�8&�3 (��90 B/�s1q91����@202��6 3���A�R�U2� d��2 bI2h`��4�᪂2�L4���19v Q�2�*�u2d�Tpt2� ��EH�a2hP�$�5��F�!U2�p�p
�2�p���@5�0-@��84 @�9��TX@�� :�e5�`rb26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0`@�gqGA���a52ѐ��Ḳ6�60ہ5�� ׁ2��8�E��9��EU5@ٰ\�q5�hQ`S�2ޖ5�p\�w�۲�pJ �-P��5��p1\t�H�4��PeCH�7j��phiw��@��P�x��559 ldu� P�D���Q �@������� �`.���P>��8�581l�"�q58�!AM۲�T�A iC�a58�9��@�x����5 �a��12׀0.�1����,�2����,�!P\�h8��Lp ��,�7z��6�0840\��ANRS 0C}A`��p��{��ran���FRA��Д�� ����A%���ѹ�� ������(����Ќ� ��З���������������$�G��1���⨂��������� xS�`q� � �����`64��M���iC/50T-�H������*��)p46��� C��N�����m75s֐� Sp��b46��v��༌ГM-71?�70�З����42�������C��-�а�70H�r�E��/h����O$��rD���c7c7C�q���ą���L��/��2\?imm7c7�g� ������`���(� ��e�����"��������a r��c�T,�Ѿ�"��,�� ��xx�Ex�m77t����k���5�����v)�iC��-HS -� B
_�>���+�Т�7U�]���M*h7�s��7������-9?�/260L_������QB�������]�9p�A/@���q�S��х���h6k21��c��92�������.�)92c 0�g$�@�����)$p��5$���pylH"O"
�21���t?�350����p���$�
�� �350!���0��9�U/�0\m9��M9AA3��4%� s��3M$��X%u���"him98J3����� �i d�"m4~�103�p�� ����h794̂�&R���H�0���� \���g�5AU��՜� �0���*2��00��#06�АՃ���!07{r ����� ���kЙ@����EP�#������?�p�#!�;&07\;!�B1P�߀A��/��CBׂ2�!�:/��?8�ҽCD25L�����0�"l�2BAL
#��B��\20�2 _�r�re���X��1@��N����A@��z��`C�pU��`��#04��DyA�\�`fQ��sU���\��5  ���� p�^P��<$8�5���+P=�ab1l��1LT��lA�8�!uDnE(�20�T��J�1 e�bH8�5���b�Ռ�5[�16Bs��������d�2��x��m6t !`Q����bˀ���b#�(�6iB;S�p�! ��3� ��b�s��-`�_�W8�_���&�6I	$�X5�1�Uc85��R�p6S� ���/�/+q�!�q��`񈓃6o��5m[o)�m�6sW��Q�?��set06p ��3%H�5��10p$����g�/�JrH�� � ��A�856�����F�� ���p/2��h�܅�✐)�5��̑v��(��m6��Y�H�ѝ̑�m�6�Ҝ��a6�DM�����-S�+��H 2�����Ҽ�� �r ̑��✐��l����p1���F���2�\wt6h T6H�� ��Ҝ�'Vl���� ���V7ᜐ/����;3A7��p~S��������4�`圐�V�T��!3��2�PM[�p�%ܖO�chn��vel5����Vq���_arp#��̑�.�~��2l_hemq$8�.�'�6415��� 5���?����F������5g�L�ј[���1���𙋹1����M7NU�М��eʾ����uq$D;��-�!4��3&H�f�c�Ĝ� h������u�� �㜐��ZS�!ܑ4�&��M-����S�$̑�ք �� 0��<������07shJ�H �v�À�sF��S*� ����̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(UL� &�(�,���0�\�?����̑�a�� xS�P���a�e�w�2ȫ�(�	�2�C��A/����\�+p�����2�1 (ܱ�CL S ����B̺��7F��h�?�<�lơ1L� ���c� ���u9�0����e/q��O���98�K��r9 (��,��Rs�ז�5�G�m20c��i��w�A2��:�0`�$��2�2 l�0�k�X�S� ,�ι�2��O���1!4�1w���2T@� _std��G�y� �ң�<H� jdgm���� w0\� �1L���	�P��~�W*�b��t 5P������3�,����E{������LL��5\L��3��L�|#~���~!���4��#��O����h�L6 A�������2璥���44�����[6\j4s��·��@�#��ol�E"w�8P k�����?0xj�H1�1`Rr�>��]�2a�#2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l��0`�&�"��|�`Am1�2@��ػ��3�HqB ��K�R��ˑb�W� ��Fs���)�ѐ�!����a�1����5��16�16C��C<����0\imBQ���d����b��\B5�-���DiL���O�_�<ѠPEtL�E�RH��ZǠPgω�am1l ��u���̑�b�<����<�$�T�̑�F�����Ȋ�Dpb��X"x��hr��p� ����^P��9�0\� �j971\kckrcfJ�F�s������c��e "CTM�E�r���ɛ��a�`main.[��g�`Grun}�_vc�# 0�w�1Oܕ_u����bctme��Ӧ�`�ܑ�j735�-� KAREL U�se {�U���J���1���p� U ̑�9�B@��L�9����7j[�atk208 "K��Kя��\��9��a��̹�����cKRC�a�o ��kc�qJ�&s��� ��Grſ�fsD��:y�0�s�ˑ1X\j|хr�dtB�, ��`.	v�q�� �sǑIf��Wfj52�TKQu�to Set��J�� H5K536�(�932���91�5�8(�9�BA�1(�7�4O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v���! conre;a�#�Controlw Re�ble��CNRE(�T�<�4��2���D�)���S�55i2��q(g�� (����4X�cOux�\s�futs�UTS `�i�栜���t�棈���? 6�T�!�S#A OO+D6����������,!��6�c+� igt�t6iB��I0�TW8 �0��la��vo58�o�b@Få򬡯i�Xh���!Xk�0Y!8\m6e�!6EC���v��6���������<1!6�A���A�6s��ƀ�U�g�T|ώ���rE1�qR��˔Z4�T������,#�eZp)g ����<ONO0���uJ���tCR;��F�a� �xSP�f��prdsuchk �1���2&&?���t��*D %$�r(�✑�娟:r���'�s�qO��<s�crc�C�\At�trldJ"o�\�V�|���Paylo�nfirm�l�!�87��7��A�3ad�! �?ވI�?hplQ��3��3"�q��x pl�`���d87��l�calC�u�Du���;��movx�����initX�:s8O��a�r4 ���r67A4|�e GeneratiڲĐ��7g2q$��g =R� (Sh��c ,|�bE��$ԒA\�:�"��4���4�4�. sg��5��F$d6"e;Qp? "SHAP�T�Q ngcr pGC��a(�&"� ��"G3DA¶��r6�"�aW�/�$dataxX:s�"tpad��<[q�%tput;a__�O7;a�o8�1�yl+s��r�?�:�#�?�5x$�?�:c O�:y O�:H�IO�s`O%g�q�ǒ�?�@0\��"o�j�92;!�Ppl.C�ollis�QSkip#��@5��@J��D ��@\ވ�C@X��7��7�|s2��potcls�LS��DU�k?�\_ et1s�`�< \�Q䜐�@���`dcKqQ�F�C;��J,�n��` (��4eN����T�{���'j(�c������/IӸaȁ��̠GH�����зa��e\mcclmt "CLM�/��� �mate\��lmpALM�?>p7qCmc?����2vm�qp��%�3s��_sv90<�_x_msu�2L�^v_� K�o�{in��8(3r<�c_lo�gr��rtrcW� �v_3�~yac��d�<�ten��der$cCe�' Fiρ�R��Q��?�l�enteAr߄|��(Sd��V1�TX�+fK�r�a�99sQ9+�5�r�\tq\� "FN�DR���S�TDn$LAN]G�Pgui��D�`���S������sp�!ğ֙uf�ҝ�s����$�����e+�=�� �������������w�H�r\fn_�ϣ��|$`x�tcpma��- TCP�����?R638 R�Ҭ���38��M7p, ���Ӡ�$Ӡ�8p0Р��VS,�>�tk��99 �a��B3���PզԠ��0D�2�����UI��t� ��hqB���8��������p���re�ȿ��exe@4φ�B���pe38�ԡG�rmpWXφ�var@�φ�@3N�����vx�!ҡ���q�RBT �$cOPTN ask E0��1��R MAS0�H5�93/�96 H5�0�i�480�5�H0��m�Q�K��7�0�g�Pl�h0ԧ�2�ORDP��@"��_t\mas��0�a@��"�ԧ�����k�� �R����ӹ`m��bL��7�.f��u�d���r��splay�D�E���1w�UPD�T Ub��887 M(��Di{���v�� ��Ԛ⧔��#�B���|����o  ��� �a�䣣��60q��B�����qscan0��B���ad@�������q`�䗣��#��К�`2�� vl v��Ù�$�>�b����! S��Easyy/К�Util��|룙�511 J������R7 ��Nor|֠��inc),<6Q�� �`c��"4�[���986FVRx� So����q�nd 6����P��4�a\ (�@�
  �������d���K�bdZ���men�7���- Me`t!yFњ�Fb�0�T�Ua�577?i 3R��\�5�u?��!� n���f���<���l\mh�Ц�pűE|hmn�	���<\O���eD�1�� l!��y��Ù�\|p����B���Ћmh�@��:. aG!���/�t��55�6�!X�l�.u�s��Y/k)ensu)bL���eK�h��  �B\1;5g?y?�?�?D��?*rm�p�?Ktbox O2K|?0�G��C?A%ds���?1ӛ#� �TR��/� �P�4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?�Ă�Q3t.�P׀al���P+OP51�7��IN0a��Q(8}g��PESTf3u�a�PB�l�ig�h�6��aq��P � sxS��`  n��0mbumpP�Q969g�69�Qq��P�0�baAp�@Q� �BOX��,>vchqe�s�>vetu㒼�=wffse�3� ��]�;u`aW��:z#ol�sm<ub�a-��]D�K�ibQ�c���p�Q<twaǂ tp�Q�҄Taror ROecov�b�O�P�642����a�0q��a⁠QErǃ�QCry�з`�P'�T�`��aar������	{'�p�ak971��71���m���>�pjo@t��PXc��C�1�adb� -�ail��na�g���b�QR629��a�Q��b�P  ?�
  �P���$$CL[q O����������$�PS_DI�GIT���"�!�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����*�璬1:PROD�UCT�Q0\PGSTK�bV,n��99�\����$FEAT_I�NDEX��~��� 搠I�LECOMP ;��)��"���SETUP2 �<��� � N !�_AP2BCK 1=�?  �)}6/"E+%,/i/��W/ �/~+/�/O/�/s/�/ ?�/>?�/b?t??�? '?�?�?]?�?�?O(O �?LO�?pO�?}O�O5O �OYO�O _�O$_�OH_ Z_�O~__�_�_C_�_ g_�_�_	o2o�_Vo�_ zo�oo�o?o�o�ouo 
�o.@�od�o� ��M�q�� �<��`�r����%� ��̏[�������!� J�ُn�������3�ȟ W������"���F�X� �|����/���֯e� �����0���T��x� �����=�ҿ�s�π��,ϻ�9�b�� P�/ 2) *.cVRiϳ�!�*�����������PC��7�!�FR6:D"�c��χ��T� �߽�Lը��ܮx���*.F��>� �	N�,�k��ߏ��STM �����Q������!�iPe�ndant Pa'nel���H��F����4������GIF�������u����JPG&P��<�����	PAN?EL1.DT�́������2 �Y�G��
3w�����//�
4�a/�O///��/�
TPEIN�S.XML�/����\�/�/�!Cus�tom Tool�bar?�PA?SSWORD/�?FRS:\R??� %Passw�ord Config�?��?k?�?O H�6O�?ZOlO�?�OO �O�OUO�OyO_�O�O D_�Oh_�Oa_�_-_�_ Q_�_�_�_o�_@oRo �_voo�o)o;o�o_o �o�o�o*�oN�or ��7��m� �&���\����� y���E�ڏi������ 4�ÏX�j�������� A�S��w�����B� џf�������+���O� ��������>�ͯ߯ t����'���ο]�� ���(Ϸ�L�ۿpς� Ϧ�5���Y�k� ߏ� $߳��Z���~�ߢ� ��C���g�����2� ��V����ߌ���?� ����u�
���.�@��� d������)���M��� q�����<��5r �%��[� &�J�n� �3�W���"/ �F/X/�|//�/�/ A/�/e/�/�/�/0?�/ T?�/M?�??�?=?�? �?s?O�?,O>O�?bO �?�OO'O�OKO�OoO �O_�O:_�O^_p_�O �_#_�_�_Y_�_}_o�_�_Ho)f�$FI�LE_DGBCK� 1=��5`��� (� �)
SUMM?ARY.DGRo�\OMD:�o�o
`�Diag Su�mmary�o�Z
CONSLOG�o��o�a
J�aCo�nsole lo�gK�[�`MEMCHECK@'�o��^qMemor?y Data��W߁)�qHADOW���P��s�Shadow ChangesS��-c-��)	F�TP=��9����w�`qmment T�BD׏�W0<�)�ETHERNE�T̏�^�q�Z��a�Ethernet� bpfigura�tion[��P��DCSVRFˏ��Ï�ܟ�q%�� v�erify alylߟ-c1PY���DIFFԟ��̟a���p%��dif!fc���q��1X�?�Q�� ����{X��CHGD��¯ԯi��px��� �¤�2`�G�Y�� 1��� �GD��ʿ�ܿq��p���Ϥ�F�Y3h�O�a��� 1��(�GD���ψ��y��p�ϡ�0��UPDATES.��Ц��[FRS:�\�����aUpd�ates Lis�t���kPSRBW�LD.CM.��\���B��_pPS_R?OBOWEL���_ ����o��,o!�3��� W���{�
�t���@��� d�����/��Se �����N�r � =�a�r �&�J���/ �9/K/�o/��/"/ �/�/X/�/|/�/#?�/ G?�/k?}??�?0?�? �?f?�?�?O�?OUO �?yOO�O�O>O�ObO �O	_�O-_�OQ_c_�O �__�_:_�_�_p_o �_o;o�__o�_�o�o $o�oHo�o�o~o�o 7�o0m�o� � �V�z�!��E� �i�{�
���.�ÏR� ���������.�S�� w������<�џ`��� ���+���O�ޟH��� ���8���߯n����$FILE_��{PR��������� ��MDONLY 1�=4�� 
 ���w�į��诨�ѿ �������+Ϻ�O�޿ sυ�ϩ�8�����n� ߒ�'߶�4�]��ρ� ߥ߷�F���j���� ��5���Y�k��ߏ�� ��B�����x����1� C���g������,��� P���������?���Lu�VISBC�KR�<�a�*.V�D|�4 FR:�\��4 Vi�sion VD file� :L bpZ�#��Y �}/$/�H/�l/ �/�/1/�/�/�/�/ �/ ?�/1?V?�/z?	? �?�???�?c?�?�?�? .O�?ROdOO�OO�O ;O�O�OqO_�O*_<_ �O`_�O�__%_�_��MR_GRP 1�>4�L�UC4�  B�P	 �]�ol`�*u����RHB� ��2 ���� ��� ��� He�Y�Q`orkbIh�o�Jd�o�Sc�o�oE��� LZo�J�9�F�5U�a�R�J]�o�o �8�e�B����A�b(�Q6���;o}=���=��lq��Q=�ȱxq�o� F@ �r�d�a�}J��NJk��H9�Hu���F!��IP��s}?�`�.9��<9�8�96C'6<,6\b~+A��,�e�P���t�A�PA�����|�ݏx��� %��I�4�F��j��� ��ǟ���֟��!���E�`r�UBH�P@�c������ů�R
6��P;�uP;��˯��e�Q cB�x�P5���@�33@����4�m�,�@UU�U��U�~w�>u.�?!x�^���ֿ���3�R�[z��=�̽=V6�<�=�=��=$q��~��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�Ϡ Cώ���C�
�P��P'�6��_V�  m�o��To��xo�ߜo ������A�,�e�P� b���������� ���=�(�a�L���p� ���������������� *��N9r]�� ������8 #\nY�}�� �����/ԭ//A/ �e/P/�/p/�/�/�/ �/�/?�/+??;?a? L?�?p?�?�?�?�?�? �?�?'OOKO6OoO�O HߢOl��ߐߢ��O��  _��G_bOk_V_�_z_ �_�_�_�_�_o�_1o oUo@oyodovo�o�o �o�o�o�oN u����� ����;�&�_�J� ��n�������ݏȏ� �%�7�I�[�"/�� ������ٟ������� 3��W�B�{�f����� ��կ�������A� ,�e�P�b��������O �O�O��O�OL�_ p�:_�����Ϧ����� ���'��7�]�H߁� lߥߐ��ߴ������� #��G�2�k�2��V w�����������1� �U�@�R���v����� ��������-Q �u���r��6 ��)M4q \n������ /�#/I/4/m/X/�/ |/�/�/�/�/�/?ֿ �B?�f?0�BϜ?f� �?���/�?�?�?/OO SO>OwObO�O�O�O�O �O�O�O__=_(_a_ L_^_�_�_�_���_�� o�_o9o$o]oHo�o lo�o�o�o�o�o�o�o #G2kV{� h������� C�.�g�y�`������� ���Џ���?�*� c�N���r�������� ̟��)��M�_�&? H?���?���?�?�?�� ��?@�I�4�m�X�j� ����ǿ���ֿ��� �E�0�i�Tύ�xϱ� ����������_,��_ S���w�b߇߭ߘ��� ��������=�(�:� s�^��������� ��'�9� �]�o��� ��~����������� ��5 YDV�z ������1 U@yd��v� ����/Я*/��
/ �u/��/�/�/�/�/ �/�/??;?&?_?J? �?n?�?�?�?�?�?O �?%OOIO4O"�|OBO �O>O�O�O�O�O�O!_ _E_0_i_T_�_x_�_ �_�_�_�_o�_/o�� ?oeowo�oP��oo�o �o�o�o+=$a L�p����� ��'��K�6�o�Z� �����ɏ��폴�  ��D�/ /z�D/�� h/ş���ԟ���1� �U�@�R���v����� ӯ������-��Q� <�u�`���`O�O�O�� �޿��;�&�_�J� oϕπϹϤ������ ��%��"�[�F��Fo �ߵ����ߠo��d�!� ��W�>�{�b��� ������������A� ,�>�w�b����������������=���$FNO ����\_�
F0l q � FLAG>�(�RRM_CHKT_YP  ] ���d �] ��O=M� _MIN� 	����� �  �XT SSB_CF�G ?\ �����OTP_DEF_OW  	���,IRCOM�� >�$GENO�VRD_DO���<�lTHR� �d�dq_ENB�] qRAVC_GRP 1@�I X(/ %/ 7//[/B//�/x/�/ �/�/�/�/?�/3?? C?i?P?�?t?�?�?�? �?�?OOOAO(OeOpLO^O�OoROU��F\� ��,�B,�8�?����O�O�O	__���  DE_�Hy_�\@@m_B�=�vR/���I�O�SMT�G��SUoo&oRHoOSTC�1H�I�� ��zMS5M�l[bo�	127.0�`=1�o  e�o�o �o#z�oFXj�|�l60s	ano?nymous��0�����Cao�
&�&��o�x��o ������ҏ�3�� ,�>�a�O�������� ��Ο�U%�7�I��]� ���f�x�������� ү����+�i�{�P� b�t���������� ��S�(�:�L�^ϭ� oϔϦϸ������=� �$�6�H�Zߩ���Ϳ s����������� � 2���V�h�z��߰� ��������
��k�}� �ߡߣ���߬����� ����C�*<Nq� _������-� ?�Q�c�eJ��n� ������/ "/E�X/j/|/�/�/ �%'/?[0? B?T?f?x?��?�?�? �?�??E/W/,O>OPO�bO�KDaENT 1=I�K P!�?�O  �P�O�O�O �O�O#_�OG_
_S_._ |_�_d_�_�_�_�_o �_1o�_ogo*o�oNo �oro�o�o�o	�o- �oQu8n�� ������#�� L�q�4���X���|�ݏ ���ď֏7���[����B�QUICCA0��h�z�۟��1ܟ��ʟ+���2,����{�!ROUTE�R|�X�j�˯!P�CJOG̯��!�192.168�.0.10��}GN�AME !�J!?ROBOT�vN�S_CFG 1H��I ��Auto-sta�rted�$FTP�/���/�?޿#? ��&�8�JϏ?nπ� �Ϥ�ǿ��[������"�4�G�#������� �������������� ��&�8�J�\�n��� �����������/�/ �/F���j��ߎ����� ��������0S� T��x����� !�3��G,{�Pb t��C���� /�:/L/^/p/�/ ���	/�/=? $?6?H?Z?)/~?�?�? �?�/�?k?�?O O2O DO�/�/�/�/�?�O�/ �O�O�O
__�?@_R_ d_v_�_�O-_�_�_�_ �_oUOgOyO�O�_ro �O�o�o�o�o�o�_ &8Jmo�o�� ���o)o;oMoO !��oX�j�|�����o ď֏����/���B��T�f�x���^�ST_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
�FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@�G %j%D�F��GI6���MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�a��3Ŀ�
��؇Mr��?�9�4�"}~q�_DCd~�1PL_NAME !<u�� �!Def�ault Per�sonality� (from FwD) �4RR2k!� 1j)TEX)�TH��!�AX d �?>?P?b?t?�?�?�? �?�?�?�?OO(O:O�LO^OpO�O�O�Ox2 -?�O�O�O__0_B_T_f_x_�b<�O�_�_ �_�_�_�_o o2oDo�Voho&xRj" 1o��)&0\�b, ��9��b�a @D7�  �a?��c�a�?�`�a�aA'�6x�ew;�	l�b�	 �x7Jp��`�`�	p �< ��(p� �.r� K��K ��K�=*�J���J?���JV��kq`q�P�x�|� �@j�@T;f�r�f�q�acrs��I�� ��p����p�r�ph}�3���´  � ��>��ph�`z���꜖"�Jm�q� H�N��ac����dw��  _�  P� Q� }�� |  а��m�Əi}	'� �� �I� ��  ����:��È�È=̣��(�ts�a	����I  �n �@H�i~�ab�Ӌ�b��w��urN0�� � 'Ж�q�p@2?��@����r�q�5�C�pC0C�G@ C����`O
�A1]w@B�UV~X�
nwB0"h�A��p�ӊ�p@����aDz���֏����Я	�pv�( �� -���I��-�=��A�a��we_q�`�p �?�ff ��m��>� ����Ƽ�uq@ݿ�>1�  	P�apv(�`ţ� ��=�qst��?�嚭`x`�� <
6�b<߈;܍��<�ê<� <�&P�ό��AO��c1��ƍ�?f7ff?O�?&��qt�@�.�J<?�`��wi4��� �dly�e߾g;ߪ�t ��p�[ߔ�߸ߣ��߀�� ����6�wh�F0%�r�!��߷��1ى����E�� �E�O�G+� F�!���/���?�e�P����t���lyBL�cB ��Enw4�������+ ��R��s����������h��<��>��I��mXj���A��y�weC�������� #/*/c/N/wi�6����v/C�`� CCHs/`
=$�p�<!��!��ܼ�'�3A��A�AR1A�O�^?�$�?���5p±
=�ç>����3�W
=�#�]��;e��?������{����<��>(�B��u��=B0�������	�R��zH�F�G����G��H��U`E���C��+��}I#�I���HD�F���E��RC��j=�>
I���@H�!H��( E<YD0w/O*OONO9O rO]O�O�O�O�O�O�O �O_�O8_#_\_G_�_ �_}_�_�_�_�_�_�_ "oooXoCo|ogo�o �o�o�o�o�o�o	 B-fQ�u�� �����,��P� b�M���q�����Ώ�� �ݏ�(��L�7�p� [������ʟ���ٟ ���6�!�Z�E�W���:#1($1��9�K����ĥ%��x��Ư!3�8��<�!4Mgs���,�IB+8�J��a?���{�d�d������ȿ���ڼ%P8�P�=:GϚ�`S�6�h�z���R��������������  %�� ��h�Vߌ�z� ��&�g�/9�$�������7����A�S�e�w�  ��������������2 wF�$�&Gb���������!C����@���8�����F�� DzN��� F�P D�������)#B�'9�K]o#?��ͫ@@v
��8��8��8�.
 v���!3 EWi{�����:� ��ۨ��1��$MSKCFMAP  ��� ����(.�ONREoL  �!�9��EXCFEN�BE'
#7%^!FN�Ce/W$JOGOV�LIME'dO S"d��KEYE'�%��RUN�,�%��SFSPDTY�0g&P%9#SIGN|E/W$T1MOT�/�T!�_CE_G�RP 1p��#\x��?p��?�? �?�?�?O�?OBO�? fOO[O�OSO�O�O�O �O�O_,_�OP__I_ �_=_�_�_�_�_�_o�o�_:o�TCO�M_CFG 1qB	-�vo�o�o
Va__ARC_b"��p)UAP_CPL��ot$NOCHEC�K ?	+ �x�%7I[ m���������!�.+NO_WAIT_L 7%S2�NT^ar	+��s�_ERR_12s	)9�� ,ȍޏ���x���&��dT�_MO��t��, ��*oq�9�PA�RAM��u	+���a�ß'g{�� �=?�345678901��,��K� ]�9�i�������ɯۯ��&g�����C���cUM_RSPA�CE/�|����$?ODRDSP�c#6�p(OFFSET_�CART�o��DI�Sƿ��PEN_FILE尨!�ai��`�OPTION_I�O�/��PWORK� ve7s#  ��V�ؤ��p�4�p�	 ���p��<����RG_DSBOL  ��P#���ϸ�RIENTT5OD ?�C�� !�l�UT_SIM�_D$�"���V~��LCT w}��h�iĜa[�1�_PEsXE�j�RATv�Ш&p%� ��2^3j)TEX)TH�)�X d3����� ��%�7�I�[�m�� �������������!�3�E���2��u��� ������������c�<d�ASew� ��������썒^0OUa0o(ҿ�(����>u2, ���O ~H @D�  [?�aG?��cc��D][�Z�;��	ls��xoJ���������< ���� ��ڐH�(��H3k7H�SM5G�22G���Gp
͜��'f�/-,ڐC%R�>�D!�M#{|Z/��3�����4y H "�c/u/��/0B_���{�jc��t�!�/ �/�"t32�����/6  ���P%�Q%��%�|�T��S62�q?'e	'�� � �2I�� �  �=�+==��ͳ?�;�	�h	�0�I  ?�n @�2�.��Ov;��ٟ?&g9N�]O  ''�uDt@!� C�C�@F#�H!�/�O�O sb
����@�@�H�@�e0@B�QA�0Yv: �13Uwz$oV_�/z_e_�_�_�	��( �� -�2�1�1ta��Ua�c���:A-����.  �?�ff ���[o"o�_U�`oDX�0A8���o�j>�1'  Po�V(���e�F0�f�Y���L�?�����xb0@<�
6b<߈;�܍�<�ê<� <�&�,/aA�;r�@Ov0P�?fff?�0?&�ip�T@�.{r�?J<?�`�u#	 �Bdqt�Yc�a� Mw�Bo��7�"�[� F��j�������ُ� ���3����,����(�E�� E�~�3G+� F��a ��ҟ�����,��PP�;���B�pAZ� >��B��6�<OίD��� P��t�=���a�s���<��6j�h��7o��>�S��O��0���Fϑ�A�a�_���C3Ϙ�/�%?��?���������#	�Ę��P �N||CH���Ŀ�������@I�_�'�3�A�A�AR1�AO�^?�$��?�����±
�=ç>�����3�W
=�#�\ U��e���B��@���{����<����(�B��u��=B�0�������	�b�H�F�G����G��H��U`E���C��+��I#��I��HD��F��E��R�C�j=[�
�I��@H�!�H�( E<YD0߻������ ��� �9�$�]�H�Z� ��~������������� #5 YD}h� ������
 C.gR���� ���	/�-//*/ c/N/�/r/�/�/�/�/ �/?�/)??M?8?q? \?�?�?�?�?�?�?�? O�?7O"O[OmOXO�O |O�O�O�O�O�O�O�Ot3_Q(�������b��gUU���W_i_2�3�8�x�_�_2�4Mgs�_��_�RIB+�_�_�a���{�m iGo5okoYo�o}l��%P'rP�nܡݯ�o�=_�o�_�[R�?Q�u���  �p���o��/� �S��z
uүܠ�������ڱ�������8����  /�M��w�e��������l2 �F�$��Gb���t��a�`�p�S�C�y�@p�5�G�Y�۠�F� Dz��� F�P D�!�]����پ��ʯ�ܯ� ��~�?��W�@@�?�K��K���K���
 �|�������Ŀ ֿ�����0�B�TϸfϽ�V� ���{���1��$PAR�AM_MENU �?3���  DE�FPULSEr��	WAITTMO{UT��RCV��� SHELL�_WRK.$CU�R_STYL���	�OPT��P�TB4�.�C�R_DECSN���e�� ߑߣ���������� �!�3�\�W�i�{�����USE_PRO/G %��%����.��CCR���e�����_HOST �!��!��:���T �`�V��/�X��>��_TIME��^���  ��GDE�BUG\�˴�GI�NP_FLMSKĻ���Tfp����PG�A  ����)CyH����TYPE��������� �� -?hc u������� //@/;/M/_/�/�/ �/�/�/�/�/�/??�%?7?`?��WORD� ?	=	R}Sfu	PNSU�Ԝ2JOK�DR�TEy�]TRACECTL 1x3���� �`��`&�?�3�6DT �Qy3�%@�0Do � �c2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�Z� .O|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� �p����� *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o� $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������������(��$PG�TRACELEN�  )�  �_�(��>��_UP z����m�u�Y��n�>�_CFG �{m�W�(�~����PКӂ�DEFS_PD |��'ѶP��>�IN��T_RL }��(��8����PE_CO�NFI��~m�'�mњ��ղ�WLID����=�?GRP 1��W���)�A ����&ff(�A+3�3D�� D]� CÀ A@1�
�Ѭ(�d�Ԭ��0�~0�� 	 1�p�ح֚��� ´�����B�9�����O�9�s�(�>�T?�
5��������� =��=#�
����P;t _��������  Dz (�
 H�X~i�� ����/�/D/�//h/S/�/��
V�7.10beta�1��  A��E�"ӻ�Ay (�� ?!G��!/>���"����!����!BQ��!A\� �!���!2p����Ț/8?J?\?n?};� ���/��/�?}/�?�?OO :O%O7OpO[O�OO�O �O�O�O�O_�O6_!_ Z_E_~_i_�_�_�_�_ �_�_'o2o�_VoAo So�owo�o�o�o�o�o �o.R=v1�<�/�#F@ �y�} ��{m��y=��1� '�O�a��?�?�?���� ��ߏʏ��'��K� 6�H���l�����ɟ�� �؟�#��G�2�k� V���z��������o ��ίC�.�g�R�d� ���������п	��� -�?�*�cώ���� �������B�;� f�x�������DϹ��� ���������7�"�[� F�X��|������� ����!�3��W�B�{� f��������� ��� ��/S>wbt ������ =OzόϾψ��� �ϼ� /.�'/R�d� v߈߁/0�/�/�/�/ �/�/�/#??G?2?k? V?h?�?�?�?�?�?�? O�?1OCO.OgORO�O vO�O�O���O�O�O_ _?_*_c_N_�_r_�_ �_�_�_�_o�_)oT fx�to���/ �o/>/P/b/t/ mo�|���� ���3��W�B�{� f�x�����Տ����� ��A�S�>�w�b��� �O��џ������+� �O�:�s�^������� ͯ���ܯ�@oRodo �o`��o�o�o��ƿ�o ���*<N�Y�� }�hϡό��ϰ����� ���
�C�.�g�Rߋ� v߈��߬�����	��� -��Q�c�N�ﲟ�� ��l��������;� &�_�J���n������� ����,�>�P�:L ����������� �(�:�3��0iT �x�����/ �///S/>/w/b/�/ �/�/�/�/�/�/?? =?(?a?s?��?�?X? �?�?�?�?O'OOKO 6OoOZO�O~O�O�O�O �O*\&_8_r���_�_��$PL�ID_KNOW_�M  ��� Q�TSV ����P��?o"o4o�O�XoCoUo�o R�SM_GRP 1��Z�'0{`�@�`uf�e�`
�5� �g pk'Pe ]o�����������SMR�c�b�mT�EyQ}? yR ����������폯��� ӏ�G�!��-����� ������韫���ϟ� C���)���������`��寧���QST�a�1 1��)��v�P0� A 4� �E2�D�V�h������� ߿¿Կ���9��.� o�R�d�vψ��ϬϾϔ���2�0� Q�<3��3�/�A�S��4l�~ߐߢ��A5���������6
��.�@��7Y�k�}����8���������MAD  �)��PARNU/M  !�}o+���SCHE� S�
���f���S��UPD�f�x��_C�MP_�`H�� �'��UER_CHK-���ZE*�<RSr��_�Q_M�OG���_�X�__RES_G��!� ��D�>1bU �y�����/ �	/����+/ �k�H/g/l/��Ї/ �/�/�	��/�/�/� X�?$?)?���D?c?�h?����?�?�?�V� 1��U�ax�@c�]�@t@(@c�\�@�@D@c�[�*@��THR_INRr�J�b�U�d2FMASS?O �ZSGMN>OqCMO�N_QUEUE ���U�V P~P *X�N$ UhN�FV��@END�A��IEcXE�O�E��BE�@|�O�COPTIO�G���@PROGRAoM %�J%�@��?���BTASK_�IG�6^OCFG ���Oz��_�PDA�TA�c��[@Ц2=�DoVohozo�j 2o�o�o�o�o�o�);M jINFO
[��m��D�� ������1�C� U�g�y���������ӏ����	�dwpt�l �)�QE DIT ���_i��^WER�FLX	C�RGA�DJ �tZAЄ����?נʕFA��I�ORITY�GW�>��MPDSPNQ�����U�GD��OT�OE@1�X� _(!AF:@E� �c�Ч!tcp|n���!ud��>��!icm���?n<�XY_�Q�X�{��Q)� *�1�5��P��]�@� L���p��������ʿ ��+�=�$�a�Hυ�z��*��PORT)Q�H��P�E��_CARTREPP|X��SKSTA�H^�
SSAV�@�tZ�	2500H8�63���_x�
�'��*X�@�swPtS��ߕߧ���URGE��@B��x	WF��DO�F"[W\��������WRUP_DE?LAY �X��ԟR_HOTqX	B%��c���R_NOR�MALq^R��v�S�EMI�����9�Q�SKIP'��tUr�x 	7�1�1� �X�j�|�?�tU���� ����������$ J\n4���� ����4FX |j����� ��/0/B//R/x/�f/�/�/�/tU�$R�CVTM$��D��� DCR'����Ў!>s>.B<� >C^�>���r8�Y7){��:���YF����̮�&�w�:�o?�� <
6�b<߈;܍��>u.�?!<�&�?h?�? �?�@>��?O O2ODO VOhOzO�O�O�O�O�O �?�O�O__@_+_=_ v_Y_�_�_�?�_�_�_ oo*o<oNo`oro�o �o�o�_�o�o�o�o �o8J-n��_� ������"�4� F�X�j�U������ď ���ӏ���B�T� �x���������ҟ� ����,�>�)�b�M� �����������ïկ �Y�:�L�^�p����� ����ʿܿ� ���� 6�!�Z�E�~ϐ�{ϴ� ������-�� �2�D� V�h�zߌߞ߰����� ����
���.��R�=� v��k�������� ��*�<�N�`�r��� ������������� &J\?���� �����"4�FXj|��!GN_ATC 1�	;� AT&�FV0E0��ATDP/6/9�/2/9�AT�A�,AT�%G1%B960��+++�,��H/,�!IO_TYPE  �%��#t�REFP�OS1 1�V+O x�u/�n �/j�/
=�/�/�/Q? <?u??�?4?�?X?�?��?�+2 1�V+ �/�?�?\O�?�O�?�!3 1�O*O<OvO��O�O_�OS4 1��O�O�O_�_t_�_>+_S5 1�B_T_�f_�_o	oBo�_S6 1��_�_�_5o�o��o�oUoS7 1� lo~o�o�oH3l�oS8 1�%�_���SMA�SK 1�V/  q
?�M��XNOS/��r������!MO�TE  n��$��_?CFG ����q����"PL_RAN�G�����POWE/R ������SM_DRYPR/G %o�%�P���TART ���^�UME_PR�O-�?����$_EX�EC_ENB  y���GSPD��pՐݘ��TDB���
�RM�
�MT_�'�T����OB�OT_NAME �o����OB�_ORD_NUM� ?�b!�H863  ��կ���P�C_TIMEOU�T�� x�S23�2Ă1�� L�TEACH ?PENDAN��wƋ�-��M�aintenance Cons�䃌s�"���KC�L/Cm��

����t�ҿ No Use-��Ϝ�0��NPO�򁋁���.�CH_Lf������q	��~s�MAVAIL������糅��SPA�CE1 2��, j�߂�D��s��߂� �{S�8�?�k�v�k�Z߬� �ߤ��ߚ� �2�D� ��hߊ�|��`����� ������ �2�D� ��h��|���`�����P����y���2��� �0�B���f�����@{���3 );M_�������/� /4 4FXj|*/�� �/�/�/?(??=?5Q/c/u/�/�/G?�/ �/�?O�?$OEO,OZO6n?�?�?�?�?dO �?�?_,_�OA_b_I_w_7�O�O�O�O�O �_�O_(oIoo^oofo�o8�_�_�_�_ �_�oo6oEf){���G �No� ���
M� ���*�<�N� `�r�������w���o �収���d.�� %�S�e�w��������� ��Ǐَ���Θ8�+� =�k�}�������ůׯ ͟����%�'�X�K� ]���������ӿ�������#�E�W� `� @����� ��x�����\�e��� ��������R�d߂� 8�j߬߾߈ߒߤ��� �������0�r��� X������������8����
�ύ�_MODE  �{^��S ��{|�2�0�����3��	S|)CWOR�K_AD��q��+R  �{��`� �� _INT�VAL���d���R_OPTION�� ��H VAT_GRP 2��uwp(N�k|��_ �����/0/B/ ��h�u/T� }/�/�/ �/�/�/�/?!?�/E? W?i?{?�?�?5?�?�? �?�?�?O/OAOOeO wO�O�O�O�OUO�O�O __�O=_O_a_s_5_ �_�_�_�_�_�_�_o 'o9o�_Iooo�o�oUo �o�o�o�o�o�o5 GYk-���u �����1�C�� g�y���M�����ӏ� ��	��-�?�Q�c��� �������������ǟ�;�M�_����$�SCAN_TIM��_%}�R ��(�#((�<}04d %d 
!D�ʣ��u�/�����+U��25���@�d5�P�g��]	���������dd��x�  P���w� ��  8� �ҿ�!���D�� $�M�_�qσϕϧϹπ�������ƿv��F�X��/� �;�ob��p�m��t�_D�iQ̡  � l�|�̡ĥ������ �!�3�E�W�i�{�� ������������� /�A�S�e�]�Ӈ��� ����������) ;M_q���� ���r���j� Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�%�/  0��6��!?3? E?W?i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O*�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo�O�OJ�o �o�o�o�o�o�o  2DVhz��������
�7?  ;�>�P�b�t����� ����Ǐُ����!� 3�E�W�i�{�������ß �ş3�ܟ� �&�8�J�\�n������������ɯ���;�,� �+��	123456{78�� 	� =5���f�x�������������
�� .�@�R�d�vψϚ�� ����������*�<� N�`�r߄߳Ϩߺ��� ������&�8�J�\� n�ߒ��������� ���"�4�F�u�j�|� �������������� 0_�Tfx�� �����I >Pbt���� ���!/(/:/L/ ^/p/�/�/�/�/�/�/�2�/?�#/9?�K?]?�iCz  �Bp˚   ��h2��*�$SC�R_GRP 1��(�U8(�\x�d�@� � ��'�	 �3�1�2�4(1*� &�I3�F1OOXO}m7��D�@�0�ʛ)���HUK�L�M-10iA 890?�90;��F;�?M61C D�:��CP��1
\&V �1	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^� oOUO>oPo#G�/血��o'o�o�o�o�oB�0�rtA9A�0*  @�BuD&Xw?��ju�bH0�{UzAF@ F�`�r��o��� ��+��O�:�s��m�Bqrr����������B�͏b����7�"�[� F�X���|�����ٟğ ���N���AO�0�B��CU
L���E�jqBq=g��Ҕ�$G@�@pnϯ B���G��I
E�0EL_DE�FAULT  ~�T��E���MIPOWE?RFL  
E*���7�WFDO�� *��1ERVENT 1���`�(�� L!DU�M_EIP��>���j!AF_IN�E�¿C�!FT$������!o:�� ��a�!RPC_MAINb��DȺPϭ�t�VIS�}�Cɻ����!TMP��PU�ϫ�d���E�!
PMON_�PROXYF߮�e 4ߑ��_ߧ�f�����!RDM_SR�V�߫�g��)�!�R�Iﰴh�u�!%
v�M�ߨ�id����!RLSYNC���>�8���!gROS��4��4�� Y�(�}���J�\����� ��������7��[ "4F�j|�� ��!�Eio��ICE_KL ?�%� (%S?VCPRG1n>���3��3���4//�5./3/�6V/[/�7~/�/�H�D�/�9�/�+� @��/��#?��K? ��s?� /�?�H/ �?�p/�?��/O� �/;O��/cO�?�O �9?�O�a?�O��? _��?+_��?S_� O{_�)O�_�QO�_ �yO�_��Os�� ��>o�o}1�o�o�o �o�o�o�o;M 8q\����� ����7�"�[�F� �j�������ُď�� �!��E�0�W�{�f� ����ß���ҟ�� �A�,�e�P���t���������ί�y_D�EV ���MC:�@`]!�OUT���2��REC 1��`e�j� �	 �����˿���8ڿ��
 �`e�� �6�N�<�r�`ϖτ� ���Ϯ�������&�� J�8�n߀�bߤߒ��� ��������"��2�X� F�|�j�������� ������.�T�B�x� Z�l������������� ,P>`bt ������( L:\�d�� ��� /�$/6// Z/H/~/l/�/�/�/�/ .��/?�/2? ?V?D? f?�?n?�?�?�?�?�? 
O�?.O@O"OdORO�O vO�O�O�O�O�O�O_ _<_*_`_N_�_�_x_ �_�_�_�_�_oo8o o,ono\o�o�o�o�o �o�o�o�o "4 jX������ ����B�$�f�T� v������������؏ ��>�,�b�P�r����p�V 1�}� P�
�ܟ� G��T�YPE\��HEL�L_CFG ��.��͟  x	�����RSR�� ����ӯ������� ?�*�<�u�`������������  �%�3�E��Q�\���M�o�p�S�d��2��d]�|K�:�HK 1�H� u������� A�<�N�`߉߄ߖߨ� ����������&�8���=�OMM ��H���9�FTOV_�ENB&�1�OW_REG_UI��~�IMWAIT��a���OUT�������TIM������VAL����_�UNIT��K�1�M�ON_ALIAS� ?ew� ( he�#���������� ����);M��q ����d�� %�I[m� <������!/ 3/E/W//{/�/�/�/ �/n/�/�/??/?�/ S?e?w?�?�?F?�?�? �?�?�?O+O=OOOaO O�O�O�O�O�OxO�O __'_9_�O]_o_�_ �_>_�_�_�_�_�_�_ #o5oGoYokoo�o�o �o�o�o�o�o1 C�ogy��H� ���	��-�?�Q� c�u� �������Ϗ� ����)�;��L�q� ������R�˟ݟ�� ���7�I�[�m��*� ����ǯٯ믖��!� 3�E��i�{������� \�տ�����ȿA� S�e�wω�4ϭϿ��� �ώ����+�=�O��� s߅ߗߩ߻�f����� ��'���K�]�o�� ��>���������� #�5�G�Y��}����������n��$SMO�N_DEFPRO ������ *�SYSTEM* � d=��REC�ALL ?}�� ( �}��>Pbt�� ,�� ���;M_ q��(���� //�7/I/[/m// �/$/�/�/�/�/�/? �/3?E?W?i?{?�? ? �?�?�?�?�?O�?/O AOSOeOwO�OO�O�O �O�O�O__�O=_O_ a_s_�_�_*_�_�_�_ �_oo�_9oKo]ooo �o�o&o�o�o�o�o�o �o5GYk}� "������� 1�C�U�g�y������ ��ӏ���	���-�?� Q�c�u�����,���ϟ�������&co�py mc:di�ocfgsv.i�o md:=>i�nspiron:5072�e�w������0.�frs:o�rderfil.�dat virt:\temp\E��������(��*.d¯Ԩׯh�z������xyzrate 61ϭH�Z�����Ϣ�3����mpbackίb�tφ�n�� }*.�db6�*C�U�Y�����ߡ��3�=���2636  ��p߂ߔ�'�9�S�W�P����
�� �� ����n��勵��Z� H�Z������"�4߽� U�a�s�������E�T�`Y�����!�.x.�:\��8 O���n��%�/.a6H�� ^�&�8����� m�������Z� �/"4�Xi/{/ �/��C/��/�/? 0BTe?w?�?���I?��?�?OO��$SNPX_AS�G 1�����9A� P� 0 '%�R[1]@1.1,O 9?�#3%dO�O sO�O�O�O�O�O�O _ _D_'_9_z_]_�_�_ �_�_�_�_
o�_o@o #odoGoYo�o}o�o�o �o�o�o�o*4` C�gy���� ���	�J�-�T��� c�������ڏ���� �4��)�j�M�t��� ��ğ������ݟ�0� �T�7�I���m����� ���ǯٯ���$�P� 3�t�W�i�������� ÿ����:��D�p� Sϔ�wω��ϭ��� � ��$���Z�=�dߐ� sߴߗߩ������� � �D�'�9�z�]��� �������
����@� #�d�G�Y���}����� ��������*4` C�gy���� ��	J-T� c������/ �4//)/j/M/t/�/ �/�/�/�/�/�/?0?�4,DPARAM ��9ECA W�	��:P�4�0�$HOFT_KB_CFG  p3�?E�4PIN_SI/M  9K�6�?��?�?�0,@RVQS�TP_DSB�>��21On8J0SR }��;� & =O�{Op0�6TOP_�ON_ERR  �p4�9�APTN� �5�@�A�BRING_�PRM�O J0V�DT_GRP 1y�Y9�@  	�7 n8_(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 Dkhz���� ���
�1�.�@�R� d�v���������Џ�� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\������� ����ȯگ����"� I�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� tߛߘߪ߼������� ��(�:�a�^�p�� ���������� �'� $�6�H�Z�l�~��������������3VPRG_COUNT�6���A�5ENB��OM=�4J_U�PD 1��;8  
p2��� ��� )$6H ql~����� /�/ /I/D/V/h/ �/�/�/�/�/�/�/�/ !??.?@?i?d?v?�? �?�?�?�?�?�?OO AO<ONO`O�O�O�O�O �O�O�O�O__&_8_�a_\_n_�_�_�_Y?SDEBUG" � ��Pdk	�PSP_�PASS"B?~�[LOG ��+m�P�X�_�  �g�Q
M�C:\d�_b_M�PCm��o�o��Qa�o �vfSAV �m:dUb�U�\gSV�\TE�M_TIME 1�� (����W�T1SVGUNYS} #'k�sp�ASK_OPTICON" �gosp�BCCFG ���| �b��z`����4��X�C� |�g�����ď֏���� ��	�B�-�f�Q�c� ���������ϟ�� ,�>�)�b��YR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz��rBr�|�|� ���z� �%��I� 4�m�X���|������� �֏���3��W�B� g���x�����՟���� ����S�>�w�b� ����'2A ��ʯܯ�� ����E�0�i�T��� x���ÿտ翢���� /��?�e�1�/���/ �ϜϮ��������,� �P�>�`߆�tߪߘ� �߼��������L� :�p�^������� ����� �6�H�>/`� r�������������� �� 0Vhz8 ������
 .�R@vd�� �����//</ */L/r/`/�/�/�/�/ �/�/�/�/?8?&?\? J?�?n?�?�?�?�?�� �?OO�?FO4OVOXO jO�O�O�O�O�O�O_ _�OB_0_f_T_v_�_ �_�_z_�_�_�_oo >o,oboPoroto�o�o �o�o�o�o(8 ^L�p���� ���$��H�6�l� ~�(O����f�d��؏ ���2� �B�D�V��� ����n����ԟ
��� .�@�R�d����v��� �����Я���*�� N�<�^�`�r�����̿ ���޿��$�J�8� n�\ϒπ϶Ϥ����� ��ߊ�(�:�L���|� jߌ߲ߠ��������� �0�B�T��x�f�� ������������,� �P�>�t�b������� ��������:( JL^����� � �6$ZH ~l��^���d� � //D/2/h/V/x/ �/�/�/�/�/�/�/? 
?@?.?d?v?�?�?T? �?�?�?�?�?OO<O *O`ONO�OrO�O�O�O �O�O_�O&__6_8_ J_�_n_�_�_�_�_�_ �_�_"ooFo��po �o,oZo�o�o�o�o �o0Tfx�H �������,� >��b�P���t����� ����Ώ��(��L� :�p�^�������ʟ�� �ܟ� �"�$�6�l� Z���~�����دꯔo ��&�ЯV�D�z�h� ������Կ¿��
�� .��R�@�v�dϚτ��  ���� ��������$TBJ�OP_GRP 2�ǌ�� � ?������������_xJBЌ���9� �< ��X���� @����	 �C��} t�b  C��<��>��͘Ր���>̚йѳ33�=�CLj�f�ff?��?�ff�BG��ь�����t��ކ�>�(�\�)�ߖ�E噙�;���hCYj�� � @h��B�  �A����f��C�  Dhъ�1���O�4�N����
:���Bl^���j�i�l�l����A�ə�A�"��D9��֊=qH����нp�h�Q�;�A�j��o��@L��D	2��������$�6�>B��\��T���Q�ts>x�@33@���C���y�1�����>��Dh�����x�����<{�h�@i� ��t ��	���K& �j�n|��� p�/�/:/k/������!��	V�3.00J�m61cI�*� IԿ���/�' Eo���E��E����E�F���F!�F8���FT�Fqe�\F�NaF����F�^lF����F�:
F��)F��3G��G��G���G,I�!CH�`�C�dTDU��?D��D���DE(!/E\��E��E��h�E�ME���sF`F+�'\FD��F`�=F}'�F���F�[
F���F��M;��;Q�T,8�4`� *�ϴ?�2����3\�X/O��ESTPARS  ���	���HR@ABL/E 1����0�É
H�7 8��9
GB
H
H����
G	
HE

H
HYE��
H�
H
H6FRD	IAO�XOjO|O�O�O�ETO"_4[>_P_�b_t_�^:BS _�  �JGoYoko}o�o�o�o �o�o�o�o1C Ugy����`#o RL�y�_�_�_�_�O�O��O�O�OX:B�rNUoM  ���P��� V@P:B_CFG ˭��Z�h�@��IMEBF_TT%AU��2@��VERS�q���R 1���
 �(�/����b�  ����J�\���j�|��� ǟ��ȟ֟����� 0�B�T���x�������R2�_���@�
��MI_CHAN��� � ��DBGL�V���������E�THERAD ?U��O������h�����ROUT6�!��!����~��SNMASKD�|�U�255.���#�����OOLO_FS_DI%@�u�.�ORQCTRL �����}ϛ3r� �Ϲ���������%� 7�I�[�:���h�z߯��APE_DETA�I"�G�PON_S�VOFF=���P_?MON �֍��2��STRTCH/K �^������VTCOMPAT���O�����FPRO�G %^�%  BCKEDT-Q�<��9�PLAY&H��_INST_Mްe ������US��q��LCK���Q?UICKME�=�ރ�SCREZ�>G�tps� �� �u�z����_��@@�n�.�SR_GRP� 1�^� �O����
��+ O=sa�쀚 �
m������L/ C1gU�y �����	/�-/�/Q/?/a/�/	1?234567�0�/��/@Xt�1���
� �}ipnl�/� gen.htm�? ?2?D?V?`�Panel _setupZ<}P���?�?�?�?�?�?  �??,O>OPObOtO�O �?�O!O�O�O�O__ (_�O�O^_p_�_�_�_ �_/_]_S_ oo$o6o HoZo�_~o�_�o�o�o �o�o�oso�o2DV hz�1'�� �
��.��R��v����������ЏG���U�ALRM��G ?9� �1�#�5� f�Y���}�������џ�ן���,��P��S�EV  �����ECFG ���롽�A�� :��Ƚ�
 Q��� ^����	��-�?�Q��c�u�����������Ԇ� �����I2��?���(%D�6�  �$�]�Hρ�lϥϐ� �ϴ�������#��Gߌ��� �߿U�I�_Y�HIST 1}��  (��� ��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1����(�:�� ����962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V