��   I�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETGY��ETH_FLT�R.  $��   ��FTP_CTRL�. @ $L�OG_8	�CMO�>$DNLD_�FILTE� � S�UBDIRCAP~�  �HO��NT. 4� H�_NAME �!ADDRTY�PA H_LEN�GTH' ��z +LS D� $ROBOTyIG PEER^ބ MASKMR�U~OMGDEV�#	� RDM*~�DISABL&}���TCPIG�/ 3 $ARP�SIZ&_IP=F'W_MC��oF_IN� FA~�LASSs�HO�_� INFO��wTELK PV�b	 WOR�D  $AC�CESS_LVL�?TIMEOUT�uORT � �I�CEUS= �   ��$#  �����!�� � � V?IRTUAL�/�!�'0 �%
�*��F�����$�%����+ �����$�� �-�2%;�SHARE�D 1�) � P!�!�?���! |?�?�?�?�?O�?%O �?1OOZOOBO�OfO �O�O�O�O_�O�OE_ _i_,_�_P_�_t_�_ �_�_o�_/o�_Soo Lo�oxo�opo�o�o�o �o�o*Os6 �Z�~���� �9��]� ���D�V� ��z�ۏ����#�� �Y�H�}�@���)7z �_LIST 1�=x!1.ܒ0Ȫ�d�ە1�d�2�55.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H� ��	��-�O�5I��@��o�������O�6����8������ �$���-� ���-@�!�%�%��&!Ò�)�0H!� ����rj3_tp�d���! � �!!KC� e�0ٙ��&W�!Cm ��w����S�!CON� ��1�=�smo	n��W�