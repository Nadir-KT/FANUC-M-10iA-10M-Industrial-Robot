��   ��A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����DRYRUN�_T   � �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �   &J_ � 4 $T�YPENFST_�IDX��_IC�I�MIX_BG�-�� G_NA�Mc %$MOD�c_USdCIFoY_TI< #�MKR-  �$LINc  { x_SIZa�#� .  �$USE_FL�GA�l�i�S�IMA�Q�QB��SCANRAX��IN�I��_C7OUNrRO�_�!_TMR_VA�gyh>� i�p'` ���H��!^%�$$CLA�SS  �����!��5��5� VIRTUR �/� '|/ �%5���U����8� ��!2�%I1�+ �M?_?q?�?�?�?�? �?�?�?OO%O7OIO`[OmO��+6W?�%{�! ��0�O�O�O��,E)1%� 1�+ 4%zO*_��11_]_ <_�_�_r_�_�_�_�_ �_�_#oooYo8oJo �ono1�C���-5�4�� �b1�d,1�!�a�o.@ Rdv����� ��?~c�a1&�8� J�\�n���������ȏ�ڏ�����!�C�1}�)  U�g�y���������ӟ ���	��-��G�`� r���������̯ޯ� ��&�8�C�\�n��� ������ȿڿ���� "�4�F�Q�j�|ώϠ� ������������0� B�M�_�xߊߜ߮��� ��������,�>�P� [�t��������� ����(�:�L�^�i� ��������������  $6HZe�w�� ������  2DVh�F