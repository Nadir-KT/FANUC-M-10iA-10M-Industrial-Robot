��   9�A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���P�ASSNAME_�T   0 }$+ $'�WORD  ? L�EVEL  w$TI- OUTT�RO&F/d� $SETUP�JPROGRAM�JINSTALL�JY  $C�URR_O�US�ER�NUM�S�TPS_LOG_ZP N��$�T��N�  6 CO�UNT_DOWN��$ENB_PCMPWD � �DV�IN!s$C� CRE�OPARM:� T:DIAG:)��LVCHK!F�ULLM0�YX=T�CNTD��MENU!AUT�O, �$$C�L(   �������	��	�V�IRTUA� ���$DCS_COD�@�����  {W'_S  *%�! T&�A9�1&"!. 
 $���~-�/�/ �/�/�/�/�/??0? >?T?b?x?�?�?�?�?\��`#SUP� l+0�?�?`#F�?O|FO��  sL�pA���O z �� �V�[t&��j�� mBO�O��H�G�O��XU 