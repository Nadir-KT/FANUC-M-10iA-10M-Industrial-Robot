��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�H UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2�X�D�#
 d �$CARD_E�XIST4$FSSB_TYP~uAHKBD_S�B֒1AGN Gn �$SLOT_N�UMJQPREV�,DBU� g1G ;1_�EDIT1 �� 1G=� S<�0%$EP�O$OP�A�ETE_OKRU�S�P_CRQ�$;4�V� 0LACIw1�RAPk �1�x@ME@$D�V�Q�Pv�A{�oQL� OUzR A,mA�0�!� B� OLM_O�^eR�"�CAM_;1 �xr$ATTqR4NP� ANN�@�5IMG_HEI�GHQ�cWIDTMH4VT� �UU0F_ASPECQw$M�0EXP�v�@AX�f�CFT� X $GR�� � S�!�@B@N�FLI�`t� UI�RE 3dTuGITC�HC�`N� S�d_�L�`�C�"�`ED(lpE� J�4S�0� ��zsa�!ip;G0� � 
$WARNM�0f�!,P� �s��pNST� CORyN�"a1FLTR�u�TRAT� T�p H0ACCa1��8�{�ORI
`"S�={RT0_S�B@_�CHG,I1 [ Tp�"3I9�TY�D,P*2 �`w@� �!R*�HD�cJ* C��2���3��4��5��6���7��8��94:�qO�$ <� �$6xK3 1w`O_M|�@�C t � �E#6NGP�ABA� �c��ZQ���`����@nr��� ��P��0����x�p��PzPb26����"J��_R��BC�J��3�JVP��tB�S��}Aw��"�tP_�*0OFSzR @�� RO_K8���aIyT�3��NOM_�02�1ĥ3"��T� �� $���AxP��K}EX�� �0g0�I01��p�
$TF�a��C$MD3��T�O�3�0U� �� K�Hw2�C1|�	EΡg0wE{vF�vF�40CPp@�a2 m
P$A`PU�3N)#�dR*��AX�!sDETAI�3BUFV��p@1� |�p۶�pPIZdT� PP[�MZ��Mg�Ͱj�F[�SIMQSI�"0��A.�Ψ��'��lw 	Tp|zM��P�B��FACTrbHPE�W7�P1Ӡ��v��M]Cd� �$*1�JB�p<�*1DEC�Hښ�H�V��b� �� +PNS_E;MP��$GP���B,P_��3�p�@Pܤ��TC��|r��0�s ��b�0�� �B���!
����JR� ��SEGKFR��Iv �aR��TkpN&S,�PVF�4��� & k�Bv�u�cu��aE�� �!2��+�MQ��E�SI!Z�3����T��P������aRSINF �����kq���������LX�����F�C3RCMu�3CClpG� �p���O}���b�1��������2�V�DxIC��C���r����P��L{� EV �zF�_��F�pNB0��?������A�! �r�Rx����V�lp��2��aR�t�,�g��qRTx @#�5�5"2��uAR��:�`CX�$LG�p���B�1 `s�P�t�aA�0{�У+0R���t�ME�`!BupCrRA 3tAZ�л�pc�OT�FC�b�`�`�FNp���1��ADI+�a%��b�{�@�p$�pSp�c�`S�P���a,QMP6�`Y$�3��M'�pU��a�U  $>�TITO1�S�S�!��$��"0�DBPXWO���!��$SK4��2�@DB��"�"@�PR8� �
� ���# l>�q1$��$��
+�L9$?(�V�)%@?R4C&_?R4gENE��'~?�(�� RE�pY2(�H �OS��#$L�3$$3R�h�;3�MVOk_D@!V�ROScrr�w�S����CRIGGER�2FPA�S��7�ET�URN0B�cMR_���TUː[��0EkWM%���GN>`���RLA���Eݡ<�P�&$P�t�'�@4a��C�DϣV��DXQ��4�1��MVG�O_AWAYRM�O#�aw!� CS�_)  `IS#� �� �s3S�AQ汯 4Rx�ZSW��AQ�p�@1UW��cTNTV)�5RV
a��� |c�éWƃ��JB��<x0��SAFEۥ�V�_SV�bEXCL�UU�;��ONLĆ�cYg�~az�OT<�a{�HI_V? ��xR, M�_ *�0�� ��_z�2� ��QSGO  + �rƐm@�A�c~b����w@��V�i�b�fAN�NUNx0�$�dIDY�UABc�@Sp�i��a+ �j�f	�!�pO�GIx2,��$F��b�$ѐOT�@A� $DUMMY ��Ft��Ft±� 6�U- ` !�HE�|s��~bc�B@ �SUFFI��V4PCA�Gs5Cwu6Cq �!MSWU�. 8!�KEYI��5�TM�1�s�qoA�vINޱE��!, �/ D��HOST�P!4���<���<�0°<��p<�EM'����Z�� SBL� UL>��0  �	�����DT�01� � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0QSp�����#��SAV� ����c�S< 9�`�f�P$�0E!� YN�_B�#2 0�`D�I�d�pO|�m��#�$F�R_IC� �ENC2_Sd3  ��< 3�9���� cgp����!4�"��2�A��ޖ5���`ǻ�@�Q@K&D-!�a�AV�ER�q����DSP
���PC_�q��"��|�ܣ�VALU�3�HE�(�M�I�P)���OPPm ��TH�*��SH" T�/�Fb�;�d�����d D��q�16� H(rLL_DU ǀ�a�@��k���֠COT�"U�/��~@@NOAUTO70�$}�x�~�@s���|�C ���C�� 2iaz�L�� �8H *��L � ���Բ@sv��`�  �� ÿ���Xq��cq��P�q���q��7��8���9��0���1�1� �1-�1:�1G�1�T�1a�1n�2|�2T��2 �2-�2:�U2G�2T�2a�2nʕ3|�3�3� �3�-�3:�3G�3T�3*a�3n�4|�R�����9 <���z�ΓKI����H硵Ba�FEq@{@: ,<��&a? P_P�?��>�����E@�@�� �QQ��;fp�$TP�$V�ARI����,�UP�2Q`< W�߃TD ��g���`��������_BAC�"= T2����$)�,+r³�p IFI��p�� �q M�P"�0�F�l@``>t ;h��6����ST� ���T��M ����0	��i���F����������kRt ����FOR�CEUP�b܂FL+US
pH(N��� ���6bD_CM�@E �7N� (�v�P��REM� Fa���j���
K�	N���EFF/���@3IN�QOV���OVA�	TROV� DT)��DTMX:e �P:/���Pq�vXpCL�N _�p��@ ��	_�|��_T: �|�J&PA�QDI����1��0�Y0RQDm�_+qH���M���CL�d#�RIV�{�ϓN"EAR/�I�O�PCP��B�R��CM�@N 1b =3GCLF��!�DY�(��a�#5T��DG���� �%�?'�FSS� )��? P(q1�1��`_1"811�E�C13D;5D6�GSRA���@�����PW�ON2EBUG�S�2�C`g�ϐ_E A ���?����TERM�5B�5X��ORI�w�0C�6C`SM_�-`���0D�5���T�A�9E�5���UP>��F� -Qϒ�A�P�3�@B$S�EGGJ� EL�UU�SEPNFI���pBx��1@��4>DC$sUF�P��$����Q�@C���G�0T������SNSTj�P�ATۡg��APTH	J�A�E*�Z%qB\`@F�{E��F�q�pARxP<Y�aSHFT͢qA|�AX_SHOR$��>��6 @$GqPE���OVR���aZP�I@P@$U?r *aAGYLO���j�I�"���Aؠ��ؠERV ��Qi�[Y)��G�@R���i�e�i�R�!P�uASYM���uqA#WJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P���WkOR�@M��k0�SMT��G��GR��3�aPA�@��p|5�'�H � j��A�TOCjA7pP<]Pp$OPd�O�P�C�%�p�O!���RE.pR�C�AOX�?��Be5pR�E�ruIx'QG�e$PW�R) IMdu�RR_p$s��5��B Iz2�H8�=�_ADDR~H�H_LENG�BP�q�q:�x�R��So�mJ.�SS��SK������ ��-�SEh*���rSN�MN1K	�j�5�@r�֣OL��\�WpW�Q�>pACRO�p���@�H ����Q� ��OSUPW3�b_>�I��!q�a1�������� |��������-���X:���iIOX2S=��D�e��]���L� $��p�!_OFyF[r_�PRM_�{�aTTP_��H��M (�pOB�J�"�pG�$H�L�E�C��ٰN �s 9�*�AB_��T��
�S�`�S��L�V��KRW"duHIoTCOU?BGi�LO�q����d�0 Fpk�GpSS� ��G�HWh�wA��O.�}�`INCPUX2VISIO��!���¢.�á<�á-� ��IOLN)�P 8�7�R'�[p$SLz�bd PUT_��$dp�Pz ��^� F_AS2Q/�$LD���D�aQT U�0]P�A������PHYG灱Z���5�sUO� 3R `F� ��H�Yq�Yx�ɱvpP�Sdp���x��ٶ�E  �UJ��S����NE�WJOG��G �DIS��&�K�Ġ��3T |��AV8��`_�CTR!S^��FLAGf2&�LG�dU �n�:��3?LG_SIZ��`�ň��=���FD��I����Z �ǳ��0�� ��@s��-ֈ�-�=�-����-��0-�ISCH�_��Dq��N?���V
��EE!2�C��"n�U�����`L�Ӕ�7DAU��EA��Ġt����GHr��I��BOO)�WL ?`�� ITV���0�\�REC�SCR�f 0�a�D^�����MARG��`!P�)�T��/ty�?I�S�H�WpW�I���T�JGM���MNCH��I�FN�KEY��K��PR�G��UF��P��F�WD��HL�STP��V��@�����RSS�H�` �Q�C��T1�ZbT�R ���U �����|R��t�i���G��8PPO��6�F�z1�M��FOCU���RGEXP�TUI��IЈ�c��n ��n����ePf���!p�6�eP7�N���CAN�AI�jB��VAIL杆CLt!;eDCS�_HI�4�.��O��|!�S S�n�R��_BUFUF1XY��PT��$�� �v��f�(L6q1YY��P ������pOS1�2��3��1� 0Z �  ��aiE�\*��IDX�dP�R�hrO�+��A&STʠ�R��Yz�<! /Y$EK&CK+����Z&m&�5�0[ L��o�0��]PL�6p�wq�t^����w��7�_ \ �����а�7��#�0C��] =��CLDP��;eTRQLI�jd.�094FLGz�0r1�R3�DM�R7��LD8R5<4R5ORG.��� e2(`���V�8.��T<�4�d^ �q�<4��-4R5S�`T00m��0�DFRCLMC�!D�?�?3I@��MI�C��d_ d���R�Qm�q�DSTB�	�  �Fg�HA�X;b �H�LEXGCESZr�rBMup
�a`��B;d�!rB�`��`a��F_A@�J��$[�O�H0K�d�b \��ӂS�$M�B��LIБ}SREQUIR�R>q�\ÁޕXDEBU��DIW�ML� MP�c�b�a��P؃ӂ!BoAND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@q��o���RPST�8� e�rLOCf�RI�p�EX�f�A�p��AoAODA�QP�f X��ON��[rMF�����f)��"I��%�e��T���F�X�@IGG� g �q��"E�0��#4���$R�a%;#7y���Gx��VvCPi�DATAw�pE:�y�[��Eѭ�NVh t �$MD�qIё) �v+�tń�tH�`�P��u�|��sANSW�}��t�?�uD�)p�b�	@Ði �@�CU��V�T0�eR;R2�j Dɐ�Q�ނ�Bd$CALI��@F�G�s�2�R�IN��v�<��NT	E���kE���,��b,����_Nl��ڂЍ�kDׄRm�DI�ViFDH�@ـn��$V��'c!$��$Z������~�[��oH �$BELTbʾ�!ACCEL+8��ҡ��IRC�t�����T/!��$P)S�@#2LPq�Ɣ�83������� ��PACTH��������3̒Vp�A_�Q�.�4�Br�Cᐈ�_MGh�$DDQ���G�$FWh��p��m���숒b�DE��PPA�BNԗROTSPCEED����00J���8��@��P$U'SE_��P��sƣSY��c�A kqY�Nu@Ag��OFF��q�MOUN�NG�g�K�OL�H�INC*��a��q��Bj�L@�BENCS��q�B�đ���D��IN#"I`(���4�\BݠVEO�|w�Ͳ23_UPE�^߳LOWL���00����D���BwP���� �1RCʀƶMgOSIV�JRMO����@GPERCH  �OV��^�� i�<!�ZD<!�c��d@�P��V1�#P͑���L���EW��ĸU�P������TRK|r�"AYLOA'a �� Q-�(�<�1Ӣ`0 ���RTI$Qx�0 MO���МB R�0J��D���s�H����b�D�UM2(�S_BC?KLSH_C(��� >�=�q�#�U��ԑ���x2�t�]ACLALv�Ų�1n�P�CHKt00'%SD�RTY4� k��y�1�q_6#2�'_UM$Pj�Cw�_��SCL��ƠLMT�_J1_LO��@���q��E������8���幘SPC��7�������PCo���H�� �PU�m�C/@�"X�T_�c�CN_��N���e���SFu���V �&#����9�(���=�C�u�SH6#��c� ���1�Ѩ�o�0�͑
̨�_�PAt�h�_Ps�W�_10��4�R�01(D�VG�J� L�@J��OGW���TORQU��ON*�Mٙ�`sRHљ��_W��-�_=��C��I��UI�I�II�F�`��JLA.�1[�VC"��0�D�BO1U�@8i�B\JRKU���	@DBL_SMtd�BM%`_DLC�BGRV��C��I��H_� �*�COS+\�(LN �7+X>$C�9)I�9) u*c,)�Z2 H�ƺMY@!�( "TH|&-�)THET0�NK23I��"=�A [CB6CB=�C�A��B(261C�616SqBC�T25GTS QơC��aS$" �4xc#�7r#$DUD� EX�1s�t��B�6���A9Q|r�f$NE�DpAIB U�\B5��$!��!A�%E(G%(!�LPH$U�2׵�2S XpCc%pCr%�2�&�C(�J�&!�VAHV6H3��YLVhJVuKV�KV��KV�KV�KV�IH�AHZF`RXM��wXuKH��KH�KH�KH�KH*�IO2LOAHO�YWNUOhJOuKO�KO�KUO�KO�KO�&F�2�#1ic%�d4GSPBALANCE_�!��cLEk0H_�%S�P��T&�bc&�br&PFULC�hr�gr�r%Ċ1ky�UTOy_?�jT1T2Cy��2N&�v�ϰctw�@g�p�0Ӓ~���T���O���� INSE9Gv�!�REV�v!����DIF��1ll�w�1m
�OB�q
����MIϰ1��?LCHWAR�����AB&u�$ME�CH,1� :�@�U�AX:�P��Y�G$�8p�n 
Z��|���ROBR�CR��N�=��MSK_�`f�_p P Np_��AR����΄ݡ�1��ҰТ΀ϳ��΀"�I�N�q�MTCO�M_C@j�q � L��p��$N'ORE³5���$�or 8� GR��E�SD�0ABF�$XYZ_DA5A<���DEBU�qI���Q�s �`$�C;OD�� ��k��F���$BUF/INDXР�����MOR��t $-�U��)��r�B���������Gؒu �� $SIMUL�T ��~�� ���OB�JE�` �ADJUyS>�1�AY_Ik§�D_����C�_F-IF�=�T� �� Ұ��{��p� �����pt�@��D�FRI�ӚӥT��RO� ��E��{���OPWOܭŀv0��SY�SBU�@ʐ$SO!P����#�U"��p�PRUN�I�PA��DH�D����_O�U�=��qn�$^}�IMAG��ˀ��0P�qIM����I�N�q���RGOVCRDȡ:���|�P~���Р�0L_6p���Li��RB���0��M���EDѐF� ���N`M*���}'��˱SL�`ŀw� x $OVS�L�vSDI��DEXm�g�e�9w�����	V� ~�N���w���ІÛǖȳ�M���q<��� x �HˁE�F�ATUS
���C�0àǒ�çBTM����If�¿�4����(�ŀy �DˀEz�g���PE��r�����
���EXE��V��E�Y�$Ժ �ŀz @ˁ��UP�{�h�$�p��XN����9�H� ��PG"�{ h �$SUB��c�@_���01\�MPWAI2��P����LO��<��F�p�$RCV?FAIL_C�f��BWD"�F���DE�FSPup | Lˀ`�D�� U�UNI��S���RX`���_L�pP��̐���ā}��� B��~���|��`ҲN�`KSET��y���P� �$�~���0SIZAE�ଠ{���S<��OR��FORMA�T/p � F���rEeMR��y�UX������PLI7�ā�  $�P_GSWI�������_PL7�AL_ S�ސR�A��B��(0C��Df�$E�h����C_=�U�� � � ���~�J3�0�����TIA4��5��6��MOM������h �B�AD��*��* PU70NRW��W �U������ A$PI�6���	�� )�4l�}69��Q����c�SPEED�PG q�7�D�>D�� ��>tMt[��SAM�`痰>��MOV���$��p �5��5�D�1�$2�������{�Hip�IN?,{� F(b+=$�H*�(_$�+�+GAMM�f�1{�$GET��ĐH��D����
^pLIB�R�ѝI��$HIB��_��Ȑ*B6E��b*8A$>G086LW= e6\<G9�686��R���ٰV��$PGDCK�Q�H�_����;"��z�.%�7��4*�9� �$IM_SRO��D�s"���H�"�LE��O�0\H��6@�qR� �ŀ�P�q?UR_SCR�ӚA�Z��S_SAVEc_D�E��NO��CgA�Ҷ��@�$��� �I��	�I� %Z[�  ��RX" ��m���" �q�'"�8�H ӱt�W�UpS���v�
U�M��O㵐.'}q ��Cg���@ʣ�����S�M�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PLM���	� 0h�H�{�%X��O��z�Z�eT�M���� pS��C��O__0_B_�a:��_%�� |S��� �@	�v��v �@��ȯw�v��EM��% (�fr�B�ː��ft�P��PM��QU.� �U�Q��A�f�QTH=�HOLޫ�QHYS�ES��,�UE��B��O.#��  -�P0�|��gAQ���ʠu���O��ŀ�ɂv�-�A;ӎ�ROG��a2�D�E�Âv�_�ĀZ�INFO&��+�����b�A��킍 ((@SLEQ/�#@������o���S`�c0O�0�01E�Z0NUe�_�AUT<�Ab�COPY���(��{��@M��N������1�P�
� ��RG4I�����X_�Pl�C$�����`�W���P��j@�G���E�XT_CYCtb����p����h�_NA�!$�\�<��RO�`]�� �s m��POR�㸅����SRVt�)l����DI �T_l� ��Ѥ{�ۧ��ۧ �ۧU5٩6٩7٩8��Ҝ�S�B쐒��$R�F6���PL�A�A^�TAR��@E �`�Z�����<��d� ,(@FLq`h��@SYNL���M�C���PWRЍ�쐔�e�DELAѰ�Y��pAD#qX� �Q�SKIP�� Ĵ��x�O�`NT!� ��P_x���ǚ@ �b�p1�1�1Ǹ� ?� �?��>��>�&��>�3�>�9�J2�R;쐖 4��EX� TQ����ށ�Q����[�KFд�w�R;DCIf� �U`�X}�R�#%M!*�0��)��$RGEAR_�0IO�TJBFLG��igpERa��TC�݃������2TH2yN��� 1�b���Gq T�0 �$���M���`Ib���v�REF�1��� l�h��ENAB��lcTPE?@��� !(ᭀ����Q�#�@~�+2 H�W���2������"�4�F�X�j�3�қ{��������j�4�Ҝ��
��P.�@�R�j�5�ҝu�@����������j�6�����(:Lj�7�ҟo�����j�8�Ҡ���"4F ��SWMSK�����a���E�A��REM�OTE�����`�@ "1��Q�IO�5�"%I��P��PO9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C���t_RS232%�Sb��iDEVICEU�S#�R�RPARI�T�!OPBIT��Q��OWCON�TR��Q�ѓ�RC�U� M�SUXTA�SK�3NB��0�$TwATU�P�"�@@쐦F�6�_�PC�}�$FREEF�ROMS]p�ai�GsETN@S�UPDl��ARB�SP%0����� !m$U�SA���az9�L�EcRI�0f��pRY�5~"_�@f�P�1�!�6'WRK��D9�F�9ХFRIEND��Q4bUF��&�A@T�OOLHFMY5��$LENGTH_;VT��FIR�pqC��@�E� IUFI�N�R���RGI<�1�AITI:�xG�X��I�FG2�7G�1a����3�B�GPRR�DA��O_� o0e�I1RER�đ�3&����TC���AQJV �QG|�.2���F��1 �!d�9Z�8+5K�+5���E�y�L0�4�X ��0m�LN�T�3H@z��89��%�4�3G��IW�0�W�RdD� Z��Tܳ��K�a3d��{$cV 2��H�1��I1H�02K2sk3K3Jci�a I�i�a�L��SL��RS$Vؠ�BV�EVk�(]V*R��� �,6Lc ���9V2F{/P:B��kPS_�E��$rr8�C�ѳ$A0��wCPR���v�U�cSk��� {�@#�2��� 0����VX`�!�tX`���0P�Ё�
�5S^K!� �-qR���!0���z�NJ A)X�!h�A�@LlA��^A�THIC�1��8�����1TFE���q>>�IF_CH�3A�aI0�����G1�x�������9�Ɇ_�JF҇PR(����RVAT�� ��-p��7@����DO��E��COU(��A�XIg��OFFS=E+�TRIG�SK���c���Ѽ�e�[�K�Hxk���8�IGMAo0�A-��ҙ�ORG�_UNEV��� ��S�쐮d ӎ$������GR3OU��ݓTO2��!�ݓDSP��JOG�'��#	�_P'�2O�R���>P6KEPFl�IR�0�PM�R&Q�AP�Q��E�0q�e���SYSG��"��;PG��BRK*Rd�r�3�-�������ߒ�<pAD��ݓJ�BS�OC� N�DU�MMY14�p\@S}V�PDE_OP3�SFSPD_OVR��ٰCO��"��OR-��N�0.�F�r�.��OV�SFc�2�f��F��!4��S��RA�"LCHD}L�RECOV��0�W�@M�յ�#RO3��_�0�� @�ҹ@VER�E�$OFS�@CV� 0BWDG�ѴC���2j�
�TR�!|��E_FDOj��MB_CM��U�B �BL=r0�w�=q�t�VfQ��x0sp��_�Gxǋ�AM��k�J0������_M��2{�#�8$CA�{Й�>��8$HBK|1c��IO��.�:!aPPA"�N�3�^�F����:"�DVC_DB�C��d�w"����!"��1���ç�3����/ATIO� �q0��UC�&CAB �BS�PⳍP�Ȗ���_0c�SUBCPUq��S�Pa a� ��}0�Sb��c��r"ơ?$HW_C��� �:c��IcA�A-�l$�UNIT��l��A�TN�f����CYC=LųNECA��[��FLTR_2_F�I���(��}&��LPx&�����_SCT@SF_��F����G����FS|!�¹�CHA�A/����2��RS�D�x"ѡb�r�: _T��PRO��O�� KEM�_��8u�q u�q��D�I�0e�RAILAiC��}RMƐLOԠdC��:anq��wq��V��PR��SLQ�p�fC�ѷ 	��FUsNCŢ�rRINkP`+a�0 ��!RA� >R 
Я�ԯgWAR�BLFQ���A�����D�A�����LD@m0�aB9��nqBTIvrbؑ���PgRIAQ1�"AFS�P�!�����`%b����M�I1U�D�F_j@��y1°LM�E�FA�@HRDY4�4��Pn@RS@Q�0|"�MULSEj@xf�b�q �X���ȑ���$.A-$�1$c1Ó����� x~�EaG�0ݓ�q!AR����09>B�%��wAXE��ROB���W�A4�_�-֣SYЯ��!6��&S�'WR䩐�-1���STR���5�9�E�� !	5B��=QB90��@6������OT�0vo 	$�ARY8��w20���	%�FI���;�$LINK(�H��1�a_63��5�q�2XYZ@"��;�q�3@��1�2J�8{0B�{D0��� CFI��6G`��
�{�_J�p�6��3aOP_O42Y;5�QTBmA"2�BC
�z�DU"�6=6CTURN3�vr��E�1�9�ҍGFL��`���~ �@�5<:7��� 1�?0K�Mc�68Cb�vrb�4�ORQ��X� >8�#op������wq�Upf�����TOVE�Q��M;�E#�UK#�UQ"�VW�ZQ�W���T υ� ;����QH�!` �ҽ��U�Q�WkeK#keLcXER��	G!E	0��S�dAWaǢ�:D���7!�!AX�rB!{q��1u y-!y�pz�@z �@z6Pz\Pz� z 1v�y�y�+y �;y�Ky�[y�ky��{y��y�q�yDEBU��$�����L�!º2WG`  AB�!�,��SV���� 
w���m���w��� �1���1���A���A�� 6Q��\Q���!�m@�\�2CLAB3B�U������S w'��SER���� O� $�@� Aؑ!p�PO��Z��q0w�Ða�_MRA�ȑ� d  T�ĴERR��STYz�B�I�V3@��cΑTOQ�d:`L0� �d2� ��˰�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	^�FZN_C;FG_!� 4��?� ��|�ų����@�ȲW� p ��\$� � n���Ѵ��9c�Q��(��FA�He�,�XE�DM�(�����!s��Q�g�P{RV HEL}Lĥ� 56��B_BAS!�RSQR��ԣo �#S��T[��1r�%��2ݺU3ݺ4ݺ5ݺ6ݺ�7ݺ8ݷ��ROO0I䰝0�0NLK!�C�AB� ��ACK��IN��T:�1�@p�@ z�m�_PU!�CO� ��OU��P�� Ҧ) ��޶��T�PFWD_KAR�ӑ��RE~��P8��(��QUE������P
��CSTOPI_AL�����0&p���㰑�0SEMl�db�|�M��d�TY|�3SOK�}�DI����p�(���_TM\�MANRQ�ֿ0E�+�|�$KEYSWITCH&	����HE
�BEAT4����E� LEҒ��
�U��FO�����_O_HOM�O�7REF�PPRz�(�!&0��C+�OA��ECO��B�rIGOCM�D8׵��@8��8�` � D�1����U��&�MH�»P��CFORC��� ����OM�  G� @V��|�U,3EP� 1-�`� 3-��4��NPX_A�SǢ� 0ȰAD�D����$SIZ>��$VARݷ �TIP]�\�2�A򻡐���]�_� ��"S꣩!Cΐ��F'RIF⢞�S�"�c���NF��V ��` �� x�`SI�TqES�R6SSGL(	T�2P&��AU�� �) STMTQZP�m 6BW�P*SHsOWb��SV��\$�� ���A00P�a�6�@�J�T�5�	6��	7�	8�	9�	A �	� �!�'��0�F�0u�	f0u �	�0u�	�@u[PTu%121?1LU1Y1f1s2�	U2�	2�	2�	2�	U2�	2�	22U2%222?2LU2Y2f2s3P)U3�	3�	3�	3�	U3�	3�	33U3%323?3LU3Y3f3s4P)U4�	4�	4�	4�	U4�	4�	44U4%424?4LU4Y4f4s5P)U5�	5�	5�	5�	U5�	5�	55U5%525?5LU5Y5f5s6P)U6�	6�	6�	6�	U6�	6�	66U6%626?6LU6Y6f6s7P)U7�	7�	7�	7�	U7�	7�	77U7%727?7,iU7Y7Fi7sk]��VP�UPD��  ��|�԰���YSLOǢ� � z��и���o�E���`>�^t��АALU�ץ����CU���wF�OqID_L�ӿuH�I�zI�$FILcE_���t��$`�vJvSA��� h��~�E_BLCK��#�C,�D_CPU <�{�<�o����tJr���R ��
�PW O� ��L�A��S��������RUNF�Ɂ��Ɂ�����F�ꁡ�ꁬ��T�BCu�C� ��X -$�LEN@i��v������I���G�LOW_AXI��F1��t2X�M�����D�
 ��I�� 9��}�TOR��"��Dh��� L=�������s���#�_MA�`�ޕ��ޑTCV����T���&��@ݡ����J�����J����Mo���J�Ǜ ��)�����2�Ѓ �v�����F�JK��V�Ki�Ρv�Ρ3��J�0�ңJJڣJJ�AALң�ڣ���4�5z�&�N1�-�9���␅�L~�_�Vj�������{ ` �GROU�p�D��B�NFLI�C��REQUI;REa�EBUA��p����2¯����x�c�� \��/APPR��C����
�EN�CLOe��S_M v�,��
���� ���MC�&���g�_MG�q�C� �{ȸ9���|�BRKz�N�OL��|ĉ R��_CLI|��Ǫ�k�J����P
���ڣ�����&���/���6��6���8��r����# ��8�%�W�2�e�PATHa�z�pӠz�=�vӥ�ϰ�x�CN=�CA�����p�IN�UC��bq��-CO�UM��YZ������qE%���2����~��PAYLOA���J2L3pR_AN��<�L��F�B�6�R��{�R_F2LSHR��|�LOG��р���ӎ���ACRL_@u�������.���H�p��$H{���FL�EX
��J�� :�/�����6�2�����;�M�_�F16����n���������ȟ��Eҟ���� �,�>�P�b���d� {������������5���T��X��v��� EťmFѯ��� ����&�/�A�S��e�D�Jx�� � �������j�4pATر���n�EL  ԁ%øJ���ʰJEΧ�CTR�Ѭ�TN���F&��HAND_VB[
�pK�7� $F2{�6�, �rSWi�ED�U��� $$Mt�h�R��08��@<b 35��^6A�p3�k��q{9�t�A�̈p��A��A��ˆ0��U���D��Dʴ�P��G��ISTЙ�$A��$AN��DY ˀ�{�g4�5D���v� 6�v��5缧�^�@��P�����#�,��5�>�+p�K�� �&0�_�ER!V9�SQA'SYM��] ������x��ݑ���_SH l�������sT�(����(�:�JA���S�c�ir��_VI�#�Oh9�``V_UNI��td�~�J���b�E �b��d��d�f��n�@��������uN����2�H�������"CqEN� a�DI��>�Obt D�Dpx��� ��2IxQA ����q��-��s �� �s����� ��OMME��rr/�TVpPT�P ���qe�i����P�x ���yT�Pj� $�DUMMY9�o$PS_��RFq�vsp$:� s�8��!~q� X�����K�STs�ʰSB}R��M21_Vt�8$SV_ERt�qO��z���CLRx�EA  O�r?p? Oր� � D $�GLOB���#LO ��Յ$�o��P�!wSYSADR�!�?p�pTCHM0 �� ,����W_NA��/�e�$%�SR��l (:]8:m�K6�^2 m�i7m�w9m��9���� ���ǳ���ŕߝ�9ŕ ���i�L���m���_�_�_�TD�XSCSRE�ƀ�� ��3STF���}�pТR6�sq] _v AŁ�� T����TYP �r�K��u�!u����O�@IS�!���tD�UE{t�# ����H�S���!�RSM_�XuUNEXCEPWv��CpS_��{ᦵ�ӕ���8÷���COU ���� 1�O�UE�T�փr���PRO�GM� FLn!$CU��PO*q��c��I_�pH;� �s 8��N�_HE
p���Q��pRY �?���,�J�*���;�OUS�� �� @d���$BU�TT��R@���CO�LUM�íu�SE�RVc#=�PANE|v Ł� � �P'GEU�!�F��9�?)$HELP��WR/ETER��)״� ��Q������@`� P�P �INЊ�s�PNߠw v�1������ �v��LN�� ���r�_��k�$H�ЎM TEX�#����F�LAn +RELVB��D4p�������M��?,��ӛ$�����P=�USRVwIEWŁ� <d���pU�p0NFI<n i�FOCU��i�7PRI# m+�qއ�TRIP)�m��UNjp{t� xQP��XuWARNWu�d�SRTOLS��ҕ�����O|SOR�N��RAUư��T���%��VI|�zu�� $�PA�THg��CACH�LOG6�O�LI�MybM���'��"�HwOST6�!�rz1�R�OBOT5����IMl� D�C� �g!��E�L���i�V�CPU_AVAIYLB�O�EX7�!BQNL�(���A�� Q���Q ��ƀ� � QpC���@$�TOOL6�$�_wJMP� �I�u$SS�!&; �SHIF��|s�AP�p�6�s���R�^��OSURW�p�RADIz��2�_ �q�h�g! �q)��LUza$OUT?PUT_BM��IML�oR6(`)�@wTIL<SCO�@Ce�;��9��F ��T��a��o�>� 3�����w�2u�b��V�zu��%�DJ�U��|#�WAIET������%O{NE��YBOư� �� $�@p%�C�SBn)TPE��NEC��x"�$�t$���*B_T��R���%�qR� ���sB�%�tM�+��t�.耰F�R!݀��OPm�M�AS�_DOG�
OaT	�D����C3S�|	�O2DELAY���e2JO��n8E��S s4'#J�aP6%�����Y_��O2� �2����5��`? ���ZABCS�� � $�2��J�
�sp�$$CLAS>�����Aspx�0'@@VIRT��O.@ABS�$�1� <E� < *A tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R��d�v�����M@[�AX�Lր�&A�dC  ����IN��ā��P#RE������LARMRECO�V <I䂥�N�G�� \K	 �A   J�\�M@PoPLIC�?<E��E�Ha�ndlingTo�ol �� 
V�7.50P/28~[�  ������
�_SW�� �UP*A� ��F�0ڑ����A�0��� 20��*A��:���X��FB 7DA�5�� N'@ω�@����No�ne������ ���T��*A4_y�xl�_���V����g�UT�OB�ค����HGAPON8@��LA�ѽU��D 1<EfA����������� Q 1שI Ԁ��Ԑ�:��i�n����#B�)B ���\��HE�Z�r�HTTHKY��$BI�[�m� ����	�c�-�?�Q� o�uχϙϫϽ����� ���_�)�;�M�k�q� �ߕߧ߹�������� [�%�7�I�g�m��� �����������W�!� 3�E�c�i�{������� ��������S/A _ew����� ��O+=[a s������� K//'/9/W/]/o/�/ �/�/�/�/�/�/G?? #?5?S?Y?k?}?�?�? �?�?�?�?COOO1O OOUOgOyO�O�O�O�O �O�O?_	__-_K_Q_���(�TO4�s���DO_CLEAN��|e��SNM  9� �9oKo]ooo��o�DSPDRY�R�_%�HI��m@ &o�o�o#5GY k}����"����p�Ն �ǣ�qX�Մ��ߢ��g�PLU�GGҠ�Wߣ��PRUC�`B`9��o��=�OB��oe�SEGF��K������o %o����#�5�m���LAP�oݎ������ ����џ�����+��=�O�a���TOTA�L�.���USENUʀ׫ �X���R�(�RG_STRI�NG 1��
��M��Sc��
��_ITEM1 �  nc��.�@� R�d�v���������п �����*�<�N�`��r�I/O S�IGNAL���Tryout M�ode�Inp���Simulat{ed�Out��OVERR�`� = 100�In cycl����Prog A�bor�����S�tatus�	H�eartbeat���MH FauylB�K�AlerU� ��s߅ߗߩ߻�����8���� �S�� �Q��f�x���� ����������,�>��P�b�t�������,�WOR������V��
 .@Rdv�� �����*8<N`PO��6� ���o����� //'/9/K/]/o/�/ �/�/�/�/�/�/�/�DEV�*0�?Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO��O�O�OPALT B��A���O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:o�OGRI�p��ra�OLo �o�o�o�o�o�o *<N`r��� ���`o��RB�� �o�>�P�b�t����� ����Ώ�����(��:�L�^�p����PREG�N��.������ ��*�<�N�`�r��� ������̯ޯ����&����$ARG_���D ?	����i�� � 	$��	+[}�]}���Ǟ��\�SBN_CON?FIG i��������CII_SAVE  ���۱Ҳ\�TCEL�LSETUP �i�%HOME�_IO�͈�%M�OV_�2�8�RE�P���V�UTOB�ACK
�ƽFRA:\��� �Ϩ���'`�!��������� ����$�6�c�Z�8lߙ��Ĉ������ �������!凞��M� _�q����2����� ����%�7���[�m� �������@�������`!3E$���J�o�������I�NI�@��ε~��MESSAG�����q��ODE_!D$���O,0.ޜ�PAUS�!�~i� ((Ol� ������� / �//$/Z/H/~/l/�/�'akTSK � q�����UP3DT%�d0;�WSM_CF°�i�еU�'1GRgP 2h�93 |��B��A�/S�XSC�RD+11
1; 	����/�?�?�?  OO$O��߳?lO~O �O�O�O�O1O�OUO_  _2_D_V_h_�O	_X�>��GROUN0O��SUP_NAL��h�	�ĠV_ED�� 11;
 �%�-BCKEDT�-�_`�!oEo%����a��o����,�ߨ���e2no_��o�o�b���ee�o"�o�oED3�o��o ~[�5GED4�n#�� ~�j���ED5Z��Ǐ�6� ~���}���ED6����k�ڏ ~G���!�3�ED7��Z���~� ~�V�şןEDa8F�&o��Ů}p����i�{�ED9���W�Ư
}3�����CRo�����3��տ@ϯ����P�PNO�_DEL�_�RGE?_UNUSE�_�T�LAL_OUT �q�c�QWD_ABOR� �΢Q��ITR_RTN�=���NONSe����CAM_PARAM 1�U�3
 8
SO�NY XC-56� 2345678�90�H � �@���?���(O АV�|[r�u�~�X�HR5k�p|U�Q�߿�R57�����Aff��K�OWA SC31�0M|[r�̀�d @6�|V�� _�Xϸ���V��� ����$�6��Z�l��CE�_RIA_I8j57�F�1��tR|]��_LIO4YW=� ��P<~��F<�GP 1�,���_GYk�*C*  ��CU1� 9� @� G� Z�CLC]� d� l� s�R� ��U[�m� v� � }�� �� C�� ő"�|W��7�HEӰONFI� ��<�G_PRI 1�+P�m®/���������'CHK�PAUS�  1E� ,�>/P/:/ t/^/�/�/�/�/�/�/ �/?(??L?6?\?�?"O�����H�1�_MOR�� =�XaBiq-���5 	 �9 O�?$O@OHOZK�2	���=$9"�Q?55��C�P)K�D3P������a�-4�O__|Z
�OG_�7�PO��� ��6_��,xV�AD�B���='�)
m�c:cpmidb�g�_`��S:�)�����Yp�_)o�S`	�BBi�P�_mo8j�)�Koo�o9i+�)��og�o�o
�m�of�oGq:I~�ZDEF f8���)�R6pbuf.txtm�]n�@�����# 	`)ЖޕA=L���zMC�21�=��9����4�=�n׾�Cz�  BHBCCPU�eB�_B�y�;��>C����CnSZE@E�?{hD]^Dْ?r�����D��^��G	���F��F���Cm	fF�O��F�ΫSY����vqG���Em�J)�.���1)��<�Lq�G�x2��Ң ��� a�D�j���E��e��X�EQ��EJP F�E��F� G����F^F E��� FB� H,�- Ge��H3�Y���  >�?33 ���xV�  n2xQ@��5�Y��8B� A�AST<7#�
� �_'��%��wRSMOFSb���~2�yT1�0�DE �O c
��(�;�"�  (<�6�z�R���?��j�C4��SZm� �W��{�m�C��B�-G�C�`@$�q���T{�FPROG� %i����c�I���� �Ɯ�f�KEY?_TBL  �vM��u� �	
��� !"#$%�&'()*+,-�./01c�:;<=>?@ABC�p�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������p��������������������������������������������������������������!j�L�CK��.�j���ST�AT���_AUT/O_DO���W/��INDT_ENB�߿2R��9�+�T2<w�XSTOP\߿2�TRLl�LETE�����_SCRE�EN i�kcsc��U��MMENU 1 i?  <g\�� L�SU+�U��p3g�� ����������2�	� �A�z�Q�c������� ��������.d ;M�q���� ��N%7] �m���/� �/J/!/3/�/W/i/ �/�/�/�/�/�/�/4? ??j?A?S?y?�?�? �?�?�?�?O�?O-O fO=OOO�OsO�O�O�O �O�O_�O_P_Sy�_MANUAL���n�DBCOU�RI�G���DBNUM��p��<���
�QP�XWORK 1!R�ү�_oO.o@o|Rk�Q_AWAY�S���GCP ��=��df_AL�P�dbB�RY�������X_�p� 1"�� , 
�^���o xvJf`MT�I^�rl@��:sONTIM��M����Zv�i
õ��cMOTNEND����dRECORD 1(R�a��ua�O��q��sb� .�@�R��xZ������ �ɏۏ폄���#��� G���k�}�����<�ş 4��X���1�C��� g�֟��������ӯ� T�	�x�-���Q�c�u� ���������>��� �)Ϙ�Mϼ�F�࿕� �Ϲ���:�������%� s`Pn&�]�o��ϓ�~� ����8�J�����5�  ��k����ߡ��J� ����X��|��C�U� ���������0������	��dbTOLEoRENCqdBȺb�`L�͐PCS_?CFG )�k)wdMC:\O �L%04d.CS�V
�`c�)sA V�CH� z�`�)~���hMRC_�OUT *�[��nSGN +��e�r��#�10�-MAY-20 �09:26*V15�-JANj10:�51�k P/�Vt��)~�`�pa�m��P�JPѬVERSION S�V2.0.8�.|EFLOGIC� 1,�[ 	�DX�P7)�PF."PROG_ENB�o\�rj ULSew �T��"_WRSTJ�NEp�V�r`dEMO�_OPT_SL �?	�es
 	R575)s7)�/�??*?<?'�$TO�  �-��?&V�_@pEX�Wd�u��3PATH ASA\�?�?O/{�ICT�aFo`-��gdse�gM%&ASTBF_TTS�x�Y^C��StqqF�PMAU� \t/XrMSWR.�i��a.|S/�Z! D_N�O0__T_C_x_�g_�_�tSBL_F�AUL"0�[3wTDIAU 16M�ap��A1234567890gFP?BoTofoxo �o�o�o�o�o�o�o�,>Pb�S�pP�_ ���_s� � 0`�����)� ;�M�_�q����������ˏݏ��|)UMP��!� �^�TRp�B�#+�=�PMEfE~I�Y_TEMP9 È�3@�3A v��UNI�.(YN_?BRK 2Y)�EMGDI_ST�A�%WЕNC2_�SCR 3�� 1o"�4�F�X�fv����������#��ޑ14 ����)�;�����:ݤ5����� x�f	u�ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� �P�b�t�� ��xߞ� ����������
��.� @�R�d�v����� ��������*�<�N� ��r������������� ��&8J\n �������� "`�FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/4?,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O?�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �O�O�o�o�o
. @Rdv���� �����*�<�N� `�r����o����̏ޏ ����&�8�J�\�n� ��������ȟڟ�����H�ETMODE� 16���+ ��ƨ
R�d��v�נRROR_P�ROG %A�%��:߽�  ��TA�BLE  A�������#�L�RRS�EV_NUM  y��Q��K��S���_AUTO_?ENB  ��I��Ϥ_NOh� 7�A�{�R�  *U�������������^�+��Ŀֿ迄�H�ISO���I�}�_A�LM 18A� e�;�����+鿀e�wωϛϭϿ��_\H���  A����|��4�TCP_V_ER !A�!�����$EXTLOGo_REQ��{��V�SIZ_�Q�TOoL  ��Dz���A Q�_BW�D����r���n�_D�I�� 9���}�z���m���STE�P����4��OP_�DO���ѠFA�CTORY_TU�N�dG�EATU�RE :�����l�Hand�lingTool� ��  - C�English� Diction�ary��ORDE�AA Vis��� Master����96 H��n�alog I/O����H551��u�to Softw�are Upda�te  ��J��m�atic Bac�kup��Part�&�groun�d Edit�� � 8\apC_amera��F���t\j6R�ell����LOADR�o�mm��shq��T7I" ��co���
! o���pa�ne�� 
!���tyle se�lect��H59��nD���onit�or��48����t�r��Reliab����adinDiagnos"�����2�2 ual �Check Sa�fety UIF� lg\a��ha�nced Rob� Serv q �ct\��lUse�r FrU��DI�F��Ext. D�IO ��fiA �d��endr E�rr L@��IF��r��  �П�9�0��FCTN M�enuZ v'��7}4� TP In���fac  SU_ (G=�p��_k Excn g��3��High-S�per Ski+� � sO�H9 � mm�unic!�onsg�teur� �����V����coknn��2��EN���Incrstr�u���5.fd�KAREL C�md. L?ua�A� O�Run-;Ti� Env����K� ��+%�s#�S�/W��74��Li�censeT� � (Au* ogB�ook(Sy��m�)��"
M�ACROs,V/�Offse��ap���MH� ����pf�a5�MechStop Prot��� d�b i�S�hif���j54�5�!xr ��#��,���b ode �Switch��mK\e�!o4.�&� pro�4��g���Multi-�T7G��net.�Pos Re�gi��z�P��t� Fun���3 9Rz1��Numx ������9m�1�  A�djuj��1 J�7�7�* ����6t�atuq1EIKoRDMtot��_scove�� ���@By- }ues�t1�$Go� � U5\�SNPX b�"���YA�"LibAr����#�� �$�~@h�pd]0�Jt�s in VCC!M�����0�  �u!Ξ�2 R�0�/I��08��TMIL{IB�M J92�@�P�Acc>�F�9=7�TPTX�+�B�RSQelZ0�M8� Rm��q%��69�2��Unexce{ptr motnT  CVV�P���KC����+-��~K�  II)�VSP� CSXC�&.c��� e�"�� t�@�Wew�AD �Q�8bvr nmeYn�@�iP� a0�y�0�pfGrid~Aplay !� �nh�@*�3R�1M-1�0iA(B2015 �`2V"  F����scii�loa�d��83 M��l�����Guar�d 'J85�0�mP'�L`����stuaPat�&]$Cyc���|0�ori_ x%Dat�a'Pqu���ch��1��g`� j� RLJam�5���I_MI De-B(\A^�cP" #^0C�  etkc^0a�sswo%q�)65�0�ApU�Xnt\��Pven�CTq�H�5�0YEL?LOW BO?Y���� Arc�0vis���Ch�Weld�Qcial4Izt��Op� ��gs�` �2@�a��poG yRjT1 NE�#3HT� xyWb��#! �p�`gd`����p\� =P��JPN� ARCP*PRx�A�� OL�pwSup̂fil�pp��J�� ��cro�6�70�1C~E�d��SuS�pe�tex�$Y �P� So7 t� /ssagN5 <Q�B�P:� �9 "0�Qr�tQC��P�l0dpn�笔�rpf�q�e��ppmasc�bin4psyn��' ptx]08�H�ELNCL V�IS PKGS �Z@MB &��B� J8@IPE �GET_VAR �FI?S (Uni�� LU�OOL: �ADD�@29.F�D�TCm���E�@D�Vp���`A�ТNO� WTWTEST� �� ��!��c�F�OR ��ECT ��a!� ALSE �ALA`�CPMO�-130��� b D�: HANG F�ROMg��2��R�709 DRAM� AVAILCH�ECKS 549���m�VPCS S�U֐LIMCHK���P�0x�FF P�OS� F�� q�8-12 CH�ARS�ER6�OG�RA ��Z@AVE�H�AME��.SV���Вאn$��9�m� "y�TRCv� �SHADP�UPD�AT k�0��ST�ATI��� MU�CH ���TIM�Q MOTN-0�03��@OBO�GUIDE DAUGH���b��@$Gtou� �@C� �0���PATH�_�M�OVET�� R6�4��VMXPAC�K MAY AS�SERTjS��CY�CL`�TA��BE COR 71�1�-�AN��RC O�PTIONS  ��`��APSH-1N�`fix��2�SO���B��XO򝡞�_TP��	�i��0j��du�{byz p wa���y�٠HI������U��pb XSPD T�B/�F� \hch�ΤB0���END�C�E�06\Q�p{ s>may n@�p�k��L ��traff#�	� ��~1�from sysvar scr�0qR� ��d�DJU����H�!A��/��S?ET ERR�D��P7����NDAN�T SCREEN� UNREA V�M �PD�D��PA����R�IO J�NN�0�FI��B���GROUNנD� Y�Т٠�h�S�VIP 53 QS���DIGIT V�ERS��ká�NE�W�� P06�@C�1IMAG�ͱ���8� DI`���p�SSUE�5��EP�LAN JON� gDEL���157QzאD��CALLI�ॡQ��m���IPN�D}�IMG N9� PZ�19��MN;T/��ES ���`wLocR Hol߀�=��2�Pn� PG:t��=�M��can������С: 3D �mE2view d3 X��ea1 �0�b�pof Ǡ"H�Cɰ�ANNOT� ACCESS �M cpie$Etn.Qs a� loMd�Flex)a:��w^$qmo G�sA9�a-'p~0��h0pa���eJ AUTO-�0��!ipu@Т<ᾡ�IABLE+� �7�a FPLN: �L�pl m� M�D<�VI�и�WI�T HOC�Jo�~1Qui��"��N���USB�@�Pt & remov����D�vAxis F�T_7�PGɰCP�:�OS-144� � h s 26�8QՐOST�p  �CRASH DU���$P��WORD�.$�LOGIN̈P��P:	�0�046 issueE��H�: Slow� st�c�`6Й���໰IF�IM�PR��SPOT:�Wh4���N1STY<��0VMGR�b�N�CAT��4oRR�E�� � 58t�1��:%�RTU!Pre -M a�SE:�@!pp���AGpL��9m@all��*0va�OCB WA����"3 CNT0 �T9DWroO0al�arm�ˀm0d �t�M�"0�2|� o�Z@OME<�� ���E%  #1-�SR�E��M�st}0g �    5KA�NJI5no M�NS@�INIS�ITALIZ'� E�f�we��6@� �dr�@ fp "~��SCII L�afails w�>�SYSTE[��i��  � Mq�1�QGro8�m n@�@vA����&��n᰼0q��RWRI O�F Lk��� \r�ef"�
�up� d�e-rela�Qd� 03.�0SSc}hőbetwe4�IND ex ɰTPa�DO� l�y �ɰGigE�s�operabil.`p l,��HcB�̚@]�le�Q0cf�lxz�Ð���OS� {����v4pfigi GLA�$�c2��7H� lap�0A[SB� If��g�2 l\c�0�/��E�� EXCE �㰁�P���i�� Do0��Gd`]Ц�fq��l lxt��EFal��#0�i�O�Y��n�CLOS��SR�Nq1NT^�F�U�FqKP�ANIO V7/ॠ1�{����DB �0��ᴥ�;ED��DET|�'�� �bF�NLINEb�BUG�T���C"RLIB��A���ABC JARK�Y@��� rkey��`IL���PR��N\��ITGAR� D$��R �Er *�T���a�U�0��h�[�Z�E V� TAS�K p.vr�P�2" .�XfJ�srn8�S谥dIBP	c�v��B/��BUS��UNN� j0-�{�d�cR'���LOE�wDIVS�CULs0$cb����BW!���R~�W`P�����ITd(঱tʠ�OF���UNEXڠ+���p��FtE��SVEM�G3`NML 50�5� D*�CC_SAFE�P*� �ꐺ� PET��'P�`�gF  !���IR����c i S>� K���K�H GUN�CHG��S�MEKCH��M��T*��%p6u��tPORY_ LEAK�J����SPEgD��2Vw 74\GRI�x�Q�g��CTLN��TRe @�_�p ���EN'�IN�����0�$���r��T3)�iԗSTO�A�s�L���͐X	���q��Y� ��TO2�J m���0F<�K����DU��S��O��3 �9�J F�&���SSVGN-1#I���'RSRwQDAU�Cޱ � �T6�g��� 3�]�~��BRKCTR/"� �q\j5��_�QܺS�qINVJ0D ZO�Pݲ���s��г��Ui ɰ̒�a�DU{AL� J50e��x�RVO117 AW�TH!Hr%�N�7247%�52��|�&aol ���R���at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���Md��Rǰt� \fosB�A�0Np�c�����{�U��ROP 2��b�pB��ITP4aM��b !AUt �c0< � plete��N@� z1^qR�635 (Acc_uCal2kA���I) "�ǰ�1a\�Ps��ǐ� bЧ0�P򶲊���ig\�cbacul "A3p_ �1��ն���_etaca��AT����PC�`�����_p�.pc!Ɗ��:�circB���5��tl��Bɵ�:�fm+�Ί�V�b�ɦ�r�?upfrm.����ⴊ�xed��Ί�~�'pedA�D �}b�ptlibB�� ߆_�rt��	Ċ�_0\׊ۊ�6�fm�݊��oޢ�e��̆Ϙ���c��Ӳ�5�j>�����tcȐ��	�r����emm 1��T�sl^0���T�mѡ�#�rm�3��ub Y�q�st�d}��pl;�&�c1kv�=�r�vf�䊰���9�vi����u�l�`�0fp�q �.yf��� daq; �i Data Ac_quisi��n��
��T`��1�8�9��22 DMCM RRS2Z��75��9 3 Rg710�o59pq5\?��T "���1 (D�T� n k@��������E Ƒȵx��Ӹ�etdmm F��ER����gE<��1�q\mo?۳ �=(G���[(

�2�` ! �@J�MACRO��Sk�ip/OffseP:�a��V�4o9� &qR662���Rs�H�
 6Bq8�����9Z�43 J�77� 6�J783�o ��n�"v��R5IKCBq2� PTLC�Zg� R�3 (�s,� �������03��	зJԷ\sfm�nmc "MNM�C����ҹ�%mnf�FMC"Ѻ0ª etmcr� �8����� ,���D�� �  874\prdq>,jF0����axisHPro�cess Axe�s e�rol^P�RA
�Dp� 56 �J81j�59� 5�6o6� ���0w�6�90 98� [!IDV�1��2(x2��2ont�0�
�����m2���?C��etis "ISD��x9�� FpraxRA�M�P� D��de�fB�,�G�isb/asicHB�@޲�{6�� 708�6
��(�Acw:�����@�D
�/,��AMOX��  ��DvE��?;T��>Pi� RAFM';�]�!PAM�V�W�Ee�U0�Q'
bU�75�.��ceNe� nterface^�1' �5&!54�K��b(Devam±�/�#��Э/<�Tane`"D�NEWE���btpd/nui �AI�_s~2�d_rsono����bAsfjN��bdv_arFvf�xhp�z�}w��hkH9xs�tc��gAponlGzv{�ff��r ���z�3{q'Td~>pchampr;re�p� ^5977� �	܀�4}0��mɁ�/������lf�!�pcc7hmp]aMP&B<�� �mpev������pcs��YeS~�� Macro�O	D��16Q!)*�:$��2U"_,��Y�(PC ��$_;������o|��J�gegemQ@�GEMSW�~ZG�g�esndy��OD�n�dda��S��syT�Kɓ�su^Ҋ����n�m���L��  �	��9:p'ѳ޲���spotplus�p���`-�W�l�J�s⽱t[�׷p�key �ɰ�$��s�-Ѩ�m�~��\featu 0�FEAWD�oolo�srn'!2 �p���a�As3��tT�.� (N. A.)��!e!�J# (j�,��oBIB�o�D -�.�n��k9�"K��u[-�_���}p� "PSEq�W����wop "sEЅ�&�:�J����� �y�|��O8��5��R ɺ���ɰ[��X�� �����%�(
ҭ�q HL�0k�
�z�a !�B�Q�"(g�Q �����]�'�.����ɀ&���<�!ҝ_�#��tpJ�H�~Z��j����� y������2��e��� ���Z����V��!%���=�]�͂��^2�@i[RV� on�QYq͋JF0� 8ހ�`�	�(^�dQueue���X\1�ʖ`�+F1�tpvtsn��N�&��ftpJ0v �R�DV�	f��J1 Q4���v�en��k/vstk��mp��~btkclrq���get�����r��`kack8�XZ�strŬ�%��stl��~Z�np:!�`���q/��ڡ6!l�/Yr�mc�N+v3�_� ���l�.v�/\jF��� �`Q�΋ܒ��N50 (FRA���+��͢frap�arm��Ҁ�} 6��J643p:V�E�LSE
#�VA�R $SGSYS�CFG.$�`_U?NITS 2�DG0~°@�4Jgfr��4A�@FRL-��0ͅ�3 ې���L�0NE�:� =�?@�8�v�9~Qx3�04��;�BPRS�M~QA�5TX.$VNUM_OL��85��DJ507��l�? Functʂ"q�wAP��琉�3 HH�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6 N�kAP����S��"TPPR���Q.A�prnaSV�ZSx��AS8Dj510U�-�`cr�`8 ��ʇ��DJR`jYȑH � �Q �PJ�6�a21��48AAVM 5�Q�b0 lB�`TUP� xbJ5459 `b�`616���0VCAM 9��CLIO b1��5 ���`M�SC8�
rP R`\�sSTYL �MNIN�`J62�8Q  �`NRExd�;@�`SCH ���9pDCSU Me�te�`ORSR �Ԃ�a04 kR_EIOC �a5�`542�b9vpP<� nP�a�`�R�`7�`��MASK H�o�.r7 �2�`O'CO :��r3��p�b�p���r0X��a�`�13\mn�a39 HRM"�q�q�ҿLCHK�uO�PLG B��a03� �q.�pHCR �Ob�pCpPosi��`fP6 is[rJ�554�òpDSWĤbM�D�pqR�a37� }Rjr0 �1�s4i �R6�7��52�rs5 �2�r7 1� �P6���Regi��@T�uFRDM��uSaq%�4�`93�0�uSNBA�uSwHLB̀\sf"p�M�NPI�SP{VC�J520���TC�`"MNрT�MIL�IFV�P�AC W�pTPT�Xp6.%�TEL�N N Me�0�9m3UECK��b�`UFR�`��V�COR��VIPL:pq89qSXC�S�`�VVF�J�TP ��q��R626l�u� S�`Gސ�2�IGUI�C��PG�St�\ŀH863`�S�q�����q34sŁ684���a��@b>�3 :B��1 \T��96 .�+E�g51 y�q53�3f�b1 ���b1 n��jr9 ���`VAT9 ߲�q75 s�F�<�`�sAWSM��`�TOP u�ŀR582p���a80 
�ށgXY q���0 ,b��`885�QXрO�Lp}�"pE࠱tp��`LCMD��ET3SS���6 �V��CPE oZ1�V�RCd3
�NLH�h���001m2Ep��3� f��p��4 /1�65C��6l���7zPR��008 tB~��9 -200�`�U0�pF�1޲1 ��޲2L"���p��޲y4��5 \hmp~޲6 RBCF�`0ళ�fs�8 �Ҋ���~�J�7 rbc	fA�L�8\PC�����"�32m0u�n�K�R�ٰn�5 5EW�
n�9 z��40Y kB��3 ��6ݲ��`00iB/��6$�u��7�u��8 µ������sU0�`�t �1 05\rb��2 E���K���j�2��5˰��60��a�HУ`:�63�jAF�_����F�7 ڱ݀H�80�eHЋ��cU0��I7�p��1u��8u��9 73�������D7� ��5t�9+7 ��8U�1��2J��1�1:���h���1np�"��8(�U1��\pyl��,࿱�v ��B�854��1hV���D�4��im�с1�<���>br�3�pr�4@pGPr�6 !B���цp��1�����1�`͵155ض1g57 �2��62�S����1b��2����1Π"�2���B�6`�1<c�4 L7B�5 DR��8_�{B/��187 u�J�8 06�90� rBn�1 (��202 0EW,ѱ�2^��2��90�U2��p�2��2 b��4:��2�a"RB����9\�U2�`w�l���O4 60Mp��7��`����b�s
5 ���3����pB"9 3a ����`ڰR,:�7 �2��V�2��5@���2^��a^9��B�qr����n�5����5᥁"�8a�Ɂ}Չ5B���5����`U�A���� ��86 �6 S�0��5�p�2�#�529 �2^�Tb1P�5~�2`P���&P5��8��5��u�!�5��ٵ5+44��5��R�ąPa nB^z�c (�a4�����U5J�
V�5��1�1^��%������5 b21���gA��58W8-2� rb��5N�E�G5890r� 1�95 �"������c 8"a��|�L ���!J"E5|6��^!�6���B�"8�`#��+�8�%�6B�AME�"1w iC��622�B�u�6V��d� 4��8�4�`ANRSP�e?/S� C�5� �6� ��� \� �6� ��V� 3t��� TG20CA�R��8� pHf� 1DH�� AOE�� �� ,�|�� �0\�� �!64K��ԓrA� �1� (M-7�!/50T�[PM��P�Th:1�C�#Pe� �3��0� 5`M75T1"� �D8p� �0Gc�� u�4��i1-710i�1� Skd�7j�z�?6�:-HS,�  �RN�@�UB�f�X�=m75sA*A6a�n���!/CB�B2.6A �0;A�CIB�A�2P�QF1�UB2�21� �/70�S� �4��� �Aj1�3p���r�#0 B2\m*A@C@��;bi"i1K�u"A~A�AU� imm7c7@��ZA@I�@�Df�Ab�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5*A��EA�5B�4>\77
B7=Q�D�2�Q$B�E)7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E"l7�@7�A
1�E�V~`��W2%Q�R9ї@0L_�#����"A����b��H3s=rA/2 �R5nR4�74rNUQ1�ZU�A�s\m9
1M�92L2�!F!^Y�ps�� 2ci��-?�qhimQ�t  w043�C�p�2�mQ�r�H_ �H20��Evr�QHsXBSt62�q`s����� ��P�xq350_*A3I)�2�d�u0�@� '4kTX�0�pa3i1�A3sQ25�c��s�t�r�VR1%e�q0 
��j1��O2 �A �UEiy�.�‐ �0C2h20$CXB79#A�����M Q1]�~�� 9 �Q��?PQ��qA!Pvs � 5	15aU���?P�Ņ���ဝQ9A6�zS*�7�qb5�1��8��Q��00P(��V7]u�aitE1���ïp�?7� !?�z��rbUQRB1PM=�Qa9p��H��QQ�25L��@�����Q��@L���8ܰ��y00\r�y�"R2BL�tN�  ��� �1D�ʑ2�qeR�5���_b�3�X]1/m1lcqP1�a�ED�Q� 5F����!5���@M-16Q�� f� ��r��Q�e� ��� PN�LT_�1��i1��9453��@�e�|�b1l>F1u*AY2�
��R8�Q���RJ�J3�D}T� 85
Qg�/0��*A!P� *A�Ð𫿽�2ǿپ6t�6=Q���P�X���� AQ� g� *ASt]1^u�ajrI�B ����~�|I�b��yI�\m�Qb�I�uz�A��c3Apa9q� B6S���S��m���}�85�`N�N�   �(M���f1���6��P��161��5�s`҃SC��U��A����5\set06c��f��10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C����5�B��B��h`�F��� X0���A:���C�M��!AZ��@��4�6i����� e�O�-	���f 1��F �ᱦ�1F�8Y	���T6HL3��BU66~`���U�dU�9D20Lf0��Qv�  ��fjq��N������ 0v
� ��i	�	��72lqQ2�������� \chngmOove.V��d��|��@2l_arf 	�f~��6���� ��9C�Z���~���kr41 S���0��V���t�����U�p7nuqQ%�A]��V�1\�Qn�BJ�2W�EM!5���)�#:�64��F�e50S�\��0�=� PV���e�������E�����m7shqQSH"U��)��9�!A��(���� ,�������TR1!��,�6�0e=�4F�����2��	 R-������ �����Ж��4���LSR�)"�!lO�A��Q�) %!� 16�
U/��2�"2�E��9p���2X� SA/Ai��'�
7F�H�@ !B�0��D���5V� �@2cVE��p��T��pt갖�1L~E�#�Fd�Q��9E�#De/��RT��59���	�A�E�iR������9\m20�20��+�-u�19r4�`�E1�=` O9`�1"ae��O��2��_$W}am41��4�3�/d1c_std��1)�!�`�_T��r�_ 4\jdg�a�q�PJ%!~` -�r�+bgB��#c'300�Y�5j�QpQb1�bq��vB��v�25�U�����qm43� �Q<W�"Ps� �A��e����t� i�P�W.��c�F�X.�e�kE14�4y4�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf��`coWo!\�2a��K2A;_2��QW2�`bF�(�V11�23�`���X5�Ra21�J�*9�a:88J9X�l5�m1a첚��*���(85�&��������P6���R,52&A����,fA9IfI'50\u�z�OV
�v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&ŦP 1��vB)e�m�����ު1p� �1D��ʹ27�F�KAR�EL Use S���FCTN��� �J97�FA+�� �(�Q޵�p%�)?�Vj�9F?(�j�Rtk208 "Km�6Q�yB�j��iæPr�9�sx#��v�krcfp��RCFt3���Q��k�cctme�!ME�g����6�mainj�dV�� ��ru��kDº�c���o����&J�dt�F �»��.vrT�f�����E�%�!��5�FRj73�B�K���UER�HJn�O  J�� (ڳF���F�q�Y�&T��`p�F�z��19�tkvBr���V�h�9p�E�y�<�k������;�v���"CT��f���� )�
І��)�V	�6� ���!��qFF��1q� ��=�����O�?�$"����$��je���TC�P Aut�r�<5�20 H5�J5�3E193��9��96�!8��9��	 �B�574��52�J:e�(�� Se%!Y������u��ma�Pqtool�ԕ�����~�conrel�F�trol Rel�iable�RmvCU!��H51�����8 a551e"�CNRE¹I��c�&��it�l\s�futst "UaTա��"X�\u�� g@�i�6Q]V0�B,Eѝ6A� �Q�)C ���X��Yf�I�1|�6s@6i��T6I U��vR�d�
$e%1���2�C58�E6��8`�Pv�iV4OFH58SOteJ� mvBM6E~O58�I�0�E�#+@� &�F�0���F�P6a����)/++�</N)0\�tr1�����P ,��ɶ�rmask�i�msk�aA���k�y'd�h	A	�P�sD�isplayIm��`v����J887# ("A��+Heůצprds��Iϩǅ�Uh�0pl�2�R2���:�Gt�@��PRD �TɈ�r�C�@Fm��D��Q�AscaҦ� �V<Q&��bVvbrl �eې@��^S��&5U�f�j8710�yl 	��Uq���7�&�p��p��P^@�P�firmQ����Pp�2�=b�k�6�r�3��6��t7ppl��PL���O�p<b�ac�q	��g1�J�U�d�J��gait_9e��Y�&��Q����	�Shap��e?ration�0��R67451j9(`sGen�ms�42-f��r�p�5����2�rsgl�E��p�G����qF�205p�5pS���Ձ�retsap��BP�O�\s� O"GCR�ö? �q/ngda�G���V��st2axU��Aa]��bad�_�btputl/�&�e�>��tplibB_���=�2.����5���c3ird�v�slp���x�hex��v�re8?�Ɵx�key�v�cpm��x�us$�6�gcr��F�����8�[�q27j92�v��ollismqSk��9O�ݝ� (pl�.���t��p!o��2 9$Fo8��cg7no@ƿtptcls` C�LS�o�b�\�km�ai_
�s>�v�o	��t�b���ӿ�E�H��6�1enu5�01�[m��uti|a|$calmaUR���CalMateNT;R51%�i=1]@ -��/V� ��Z�� �tfq1�9 "K9E��L����2m�CLcMTq�S#��et ��LM3!} �F�c��nspQ�c���c�_moq��� ��c1_e�����su��ޏ� �_ �@�5�G�join�i�j��oX��ł&cWv	 ���N�v9e��C�clm�&A�o# �|$finde��0STD �ter FiOLANG���R���
��n3��z0Cen���r,������ J����� ���K�〪Ú�=���_Ӛ��r~� "FNDR��� 3��f��tguid�䙃N�."��J�tq�� ��������� ����J����_������c��	m�Z��?\fndr.��n#�>
B2p��Z�CP� Ma�����38PA��� c��6� (�� �N�B�������H 2�$�81��m_���"ex�z5� .Ӛ��c��bSа�efQ��	���RBT;�OPTN �+#Q�*$�r*$ ��*$r*$%/s#C�d/�.,P�/0*ʲD�PN��$���$*�G}r�$k Exc�'{IF�$MASK�%�93 H5�%H5�58�$548 H��$4-1�$��#1(�$�0 E�$��$-b��$���!UPDT ��B�4�b�4�2�49�0`�4a�3�9j0"M�4<9�4  ��4��4tpsh���4�P�4- DQ� �3�Q�4�R�4�pR%0�2�r�4.b
E\���5�A�4���3adq\�5K�979":E�ajO l "DQ^E^�3�i�Dq ��4ҲO ?R�? ��q�5��T���3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F��t�4��.�5y N� >�2il(in�4��31 JH1�2Q4�2�51ݠ�4rmal� �3)�REo�Z_�� �Ox����4��^F�?onorTf��7_ja�UpZҒ4l�5rmsAU��Kkg���4�$HCd\��fͲ�eڱ�4�REM����4yݱ"u@�RERG5932fO��47Z�>�5lity,�U��8e"Dil\�5�r�o ��7987�?8�25 �3hk910�3 ��FE�0=0P_�Hl\mhm�5� �qe�=$�^�
E��u<�IAymptm�U��BU��vste�y\� 3��me�b�DvI�[�Qu �:F�Ub�*_�
E&,�su��_ E�r��ox���4hu#se�E-�?�sn��������FE��,�box�����c݌,"��� ����z��M��g��pdspw)�	�� 9���b���(��1���c��Y�R��  �>�P���W��������'�0ɵ�[���͂���  �w ,�@� �zA�bumpšuf��B*�Box%��7Aǰ60�BBw���MC� (6�,f�t{ I�s� ST���*��}B�����w��"BBF
�>�`����)��\bbk968 "�4��։�bb�9va69�����etbŠ��X�����ed	�F��1u�f� �sea"������'�\��,���b�ѽ�o6�H�
�	x�$�f���!y����Q[�! tpermr�fd� TPl0~o� Recov,���3D��R642� � 0��C@}s� tN@��(U�rro����yu2r��  ?�
  �����$$CLe� O�������������$z�_DIGsIT��������.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$j����+c:PRODU�CTM�0\PGSTKD��V&ohozf�99��D����$FEAT_I�NDEX��xd���  
��`ILECOMPW ;���#��`��cSETUP2� <�e�b��  N �a�c_�AP2BCK 1�=�i  �)�wh0?{%&c�� ��Q�xe%�I� m���8��\�n� ���!���ȏW��{� �"���F�Տj���w� ��/�ğS������� ��B�T��x������ =�үa������,��� P�߯t������9�ο �o�ϓ�(�:�ɿ^� ��Ϗϸ�G���k�  �ߡ�6���Z�l��� ��ߴ���U���y�� ���D���h��ߌ�� -���Q��������� @�R���v����)��� ��_�����*��N ��r��7�� m�&�3\�i�
pP 2#p�*.VRc�*��� /���PC/1/FR6:/].��/+T�`�/�/F%�/�,�`xr/?�*.F�D8?	H#&?e<�/<�?;STM �2�?н.K �?�=i�Pendant �Panel�?;H �?@O�7.O�?y?�O:GIF�O�O�5�OoO8�O_:JPG _J_��56_�O_�_�	P�ANEL1.DT�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�WI���
TPEINS.XML���0\���qC�ustom To�olbar	���PASSWORD�yFRS:\�L�� %Pas�sword Config���֏e� Ϗ�B0���T�f��� �������O��s�� ����>�͟b��[��� '���K��򯁯��� :�L�ۯp�����#�5� ʿY��}��$ϳ�H� ׿l�~�Ϣ�1����� g��ϋ� ߯���V��� z�	�s߰�?���c��� 
��.��R�d��߈� ��;�M���q���� ��<���`������%� ��I��������8 ����n���!�� W�{"�F� j|�/�Se ��/�/T/�x/ /�/�/=/�/a/�/? �/,?�/P?�/�/�?? �?9?�?�?o?O�?(O :O�?^O�?�O�O#O�O GO�OkO}O_�O6_�O /_l_�O�__�_�_U_ �_y_o o�_Do�_ho �_	o�o-o�oQo�o�o �o�o@R�ov ��;�_��� *��N��G������ 7�̏ޏm����&�8� Ǐ\�돀��!���E� ڟi�ӟ���4�ßX� j��������įS���w������B�#��$�FILE_DGB�CK 1=���/���� ( �)
SU�MMARY.DG<L���MD:������Diag Summary���Ϊ
CONSLO�G�������D�ӱ�Console �logE�ͫ��MEMCHECK:��!ϯ���X�Mem�ory Data|��ѧ�{)��HADOW�ϣϵ��J���Shado�w Change�sM�'�-��)	FTP7Ϥ�3ߨ����Z�mment� TBD��ѧ0=�4)ETHERNET�������T��ӱEthern�et \�figu?rationU�ؠ~��DCSVRF��p�߽�����%��� verify �all��'�1PY=���DIFF�����[���%��d�iff]������1pR�9�K��� ����X��CHGAD������c��r����2ZAS�� ��GD ���k��z��FY3bI[�� �/"GD ���s/����/�*&UPDATE�S.� �/��FR�S:\�/�-ԱU�pdates L�ist�/��PSRBWLD.CM(?����"<?�/Y�PS�_ROBOWEL ��̯�?�?��?&�O -O�?QO�?uOOnO�O :O�O^O�O_�O)_�O M___�O�__�_�_H_ �_l_o�_�_7o�_[o �_lo�o o�oDo�o�o zo�o3E�oi�o ���R�v� ��A��e�w���� *���я`�������� �O�ޏs������8� ͟\�����'���K� ]�쟁����4���ۯ j������5�įY�� }������B�׿�x� Ϝ�1���*�g����� Ϝ���P���t�	�� ��?���c�u�ߙ�(� ��L߶��߂���(� M���q� ���6��� Z������%���I��� B�����2�����h�����$FILE�_� PR� ���������MDONLY� 1=.�� 
 ���q����� �����~%� I�m�2� �h��!/�./W/ �{/
/�/�/@/�/d/ �/?�//?�/S?e?�/ �??�?<?�?�?r?O �?+O=O�?aO�?�O�O &O�OJO�O�O�O_�O�9_�OF_o_
VIS�BCKL6[*�.VDv_�_.PF�R:\�_�^.P�Vision V?D file�_�O 4oFo\_joT_�oo�o �oSo�owo�oB �of�o�+�� �����+�P�� t������9�Ώ]�� ����(���L�^���� ���5���ܟk� ��� $�6�şZ��~������
MR_GRPw 1>.L���C4  B���	� W������*u���R�HB ��2 ���� ��� ���B�����Z�l��� C���D�������Ŀ���K��L5��PJ��tF�5�UT��Q�`񗲿�ֿ G,��FI�/E����.��9:��]�@�'�A&�#A~�kf��?�f�A~���r��E�� F�@ �������J���NJk�H9��Hu��F!���IP�s�?�����(�9�<9��896�C'6<,6\b��+�&�(�a�0L߅�XȞ�A��߲� v���r������
�C� .�@�y�d������ ��������?�Z�l�v��BH�� ��Ж�������
0�P=?��P�K|��ܿ�� �B���/ ��@'�33:��.�g^&�@UUU�U���q	>u.�?!rX��	�-�=[z�=����=V6<�=��=�=$q������@8�i�7G��8�D��8@9!��7�:����D��@ D�� CYϥ��C������ Q�,/������/M� �/q��/�/�/�?? :?%?^?p?[?�??�? �?�?�? O�?�?6O!O ZOEO~OiO�O�O�O�O W�ߵ��O$_�OH_3_ l_W_�_{_�_�_�_�_ �_o�_2ooVohoSo �owo�o�i��o�o�o ��);�o_J� j������� %��5�[�F��j��� ��Ǐ���֏�!�� E�0�i�{�B/��f/�/ �/�/���/��/A�\� e�P���t�������� ί��+��O�:�s� ^�p�����Ϳ���ܿ � ��OH��o�
ϓ� ~ϷϢ���������� 5� �Y�D�}�hߍ߳� ���������o�1�C� U�y��߉����� ��������-��Q�<� u�`������������� ��;&_J\ ���������� ڟ�F�j4��� ������!// 1/W/B/{/f/�/�/�/ �/�/�/�/??A?,? e?,φ?P�q?�?�?�? �?O�?+OOOO:OLO �OpO�O�O�O�O�O�O _'__K_�o_�_�_ �_l��_0_�_�_�_#o 
oGo.okoVoho�o�o �o�o�o�o�oC .gR�v��� ��	���<�`� *<��`����� ޏ��)��M�8�q�\� ������˟���ڟ� ��7�"�[�F�X���|� ��|?֯�?�����3� �W�B�{�f�����ÿ ���������A�,� e�P�uϛ�b_������ �_��߀�=�(�a�s� Zߗ�~߻ߦ������� � �9�$�]�H��l� ������������#� �G�Y� �B������� z�������
ԏ:�C .gRd���� ��	�?*c N�r����� /̯&/�M/�q/\/ �/�/�/�/�/�/�/? �/7?"?4?m?X?�?|? �?�?�?�?��O!O3O ��WOiO�?�OxO�O�O �O�O�O_�O/__S_ >_P_�_t_�_�_�_�_ �_�_o+ooOo:oso ^o�o�op��o��  ��$��o�o� ~������� 5� �Y�D�}�h����� ��׏����
�C� .�/v�<���8����� �П����?�*�c� N���r��������̯ ��)��?9�_�q��� JO�����ݿȿ�� %�7��[�F��jϣ� ���ϲ�������!�� E�0�i�T�yߟߊ��� ���߮o�o��o>� t�>��b������ �����+��O�:�L� ��p������������� 'K6oZ� Z�|�~����� 5 YDi�z� �����/
// U/@/y/@��/�/�/�/ ���/^/???Q?8? u?\?�?�?�?�?�?�? �?OO;O&O8OqO\O �O�O�O�O�O�O�O_��O7_��$FNO ���VQ��
F�0fQ kP FLA�G8�(LRRM_�CHKTYP  �WP��^P��WP�{QOM�P_MsIN�P����P��  XNPSS�B_CFG ?�VU ���_���S ooIUT�P_DEF_OW�  ��R&hI�RCOM�P8o�$�GENOVRD_�DO�V�6�flT[HR�V d�edkdo_ENBWo k`�RAVC_GRP� 1@�WCa X "_�o_1U< y�r����� 	��-��=�c�J��� n��������ȏ�� ��;�"�_�F�X���ib�ROU�`FVX�P��&�<b&�8�?��埘��������  D�?�јs���@@g�B��7�p�)�ԙ���`S+MT�cG�mM����� �LQHOSTC��R1H���P�\�at�SM��f��\���	12�7.0��1��  e��ٿ����� ǿ@�R�d�vϙ�0�*��	anonymous����������֣0�[�� � � ����r����ߨߺ��� ��-���&�8�[�I� �π������ 1�C��W�y���`�r� �����ߺ������� %�c�u�J\n�� �������M�" 4FX��i��� ���7//0/B/ T/���m/��/ �/�/??,?�/P?b? t?�?�/�?��?�?�? OOe/w/�/�/�?�O �/�O�O�O�O�O=?_ $_6_H_kOY_�?�_�_ �_�_�_'O9OKO]O__ Do�Ohozo�o�o�o�O �o�o�o
?o}_R dv���_�_oo !�Uo*�<�N�`�r� �o������̏ޏ�?�Q&�8�J�\���>�E�NT 1I�� sP!􏪟  ����՟ğ������� A��M�(�v���^��� ��㯦��ʯ+�� � a�$���H���l�Ϳ�� ���ƿ'��K��o� 2�hϥϔ��ό��ϰ� ������F�k�.ߏ� R߳�v��ߚ��߾����1���U��y�<�QUICC0��b�t����1�����%����2&���u�!ROUTERv�R�d����!PCJOG�����!192�.168.0.1�0��w�NAME �!��!ROB�OTp�S_CF�G 1H�� ��Auto�-started^�tFTP�� ����� 2 D��hz���� U��
//./�v� ��/���/�/�/ �/�/�!?3?E?W?i? �/?�?�?�?�?�?�? ���AO�?eO�/�O �O�O�O�?�O�O__ +_NO�OJ_s_�_�_�_ �_
OO.OoB_'ovO Ko]ooo�oP_>o�o�o �o�oo�o5GY k}�_�_�_�� 8o��1�C�U�$y� �������ӏf���	� �-�?�����Ə ���ϟ����� ;�M�_�q���.�(��� ˯ݯ��P�b�t��� ��m���������ǿٿ �����!�3�E�h�� {ύϟϱ����$�6� H�J�/�~�S�e�w߉� ��jϿ��������*߀��=�O�a�s��YT_ERR J5
����PDUSIZW  ��^J�����>��WRD ?�t��  guest}���%�7�I�[�m�$S�CDMNGRP �2Kt��C����V$�K��� 	P01.1�4 8��   �y����B  �  ;������ ���������
 �������������~����C.gR�|���  i  �  
��������� +��������
��k�l .r����"�l��� m
d�������_GR�OU��L�� ��	����07EQ?UPD  	պ�YJ�TYa �����TTP_AU�TH 1M�� �<!iPend�any��6�Y�!KAREL:q*��
-KC/�//A/ VISI?ON SETT�/v/�"�/�/�/# �/�/
??Q?(?:?�?�^?p>�CTRL CN����5�
��.FFF9E�3�?�FRS:DEFAULT�<�FANUC �Web Server�:
�����<�kO}O�O�O�O�O��W�R_CONFIGw O�� �?���IDL_CPU�_PC@�B���7P�BHUMI�N(\��<TGNR_�IO������PN�PT_SIM_D�OmVw[TPMO_DNTOLmV �]_PRTY�X7RTOLNK 1P����_o!o3oEoWo|io�RMASTElP���R�O_CFG��o�iUO��o�bC�YCLE�o�d@_?ASG 1Q����
 ko,>Pb t�������p��sk�bNUM�����K@�`IPCH��o��`RTRY_�CN@oR��bSC�RN����Q��� �b�`�bR���Տ���$J23_D_SP_EN	�����OBPROC��U�iJOGP1�SY@��8��?�!�T�!�?*�P�OSRE�zVKANJI_�`��o_��$ ��T�L�6͕����CL_LGP<�_����EYLOGGI�N�`��L�ANGUAGE YYF7RD w����LG��U�?⧕��x� �����Z=P��'0��$� NMC:\RSCH\00\���LN_DISP V��
���������OC�R.RDzVTA�{�OGBOOK W
{��i��ii��X�����ǿٿ������"��6	�h�����e�?�G�_BUFF 1X�]��2	աϸ� ����������!� N�E�W߄�{ߍߺ߱� ���������J�~��DCS Zr� =����^�+��ZE��������a�IOw 1[
{ ُ!� �!�1�C�U�i� y��������������� 	-AQcu��������EfPTM  �d�2/ ASew���� ���//+/=/O/�a/s/�/�/��SE�V����TYP�/??y͒��RS@"��×�FLg 1\
������ �?�?�?�?�?�?�?/?STP6��">�NGNAM�ե�Un`�UPS��GI}��𑪅mA_LOA�D�G %�%�DF_MOTN����O�@MAXUALRM<��J��@sA��Q����WS ��@C �]m�-_���MP2��7�^
{ ر�	V�!P�+ʠ�;_�/��Rr�W�_�WU�W�_��R	o�_o ?o"ocoNoso�o�o�o �o�o�o�o�o;& Kq\�x��� ����#�I�4�m� P���|���Ǐ���֏ ��!��E�(�i�T�f� ����ß��ӟ����  �A�,�>�w�Z����� ��ѯ����د��� O�2�s�^�������Ϳ����ܿ�'��BD_LDXDISAX@�	��MEMO_A�PR@E ?�+
 � *�~ϐϢ�������������@IS�C 1_�+ � �IߨT��Q�c�Ϝ� ���ߧ�����w���� >�)�b�t�[���� {����������:��� I�[�/���������� ��o�����6!Zl S��s��� �2�AS'� w����g���.//R/d/�_MS�TR `�-w%S_CD 1am͠L/ �/H/�/�/?�/2?? /?h?S?�?w?�?�?�? �?�?
O�?.OORO=O vOaO�O�O�O�O�O�O �O__<_'_L_r_]_ �_�_�_�_�_�_o�_ �_8o#o\oGo�oko�o �o�o�o�o�o�o" F1jUg��� ������B�-� f�Q���u�����ҏh/�MKCFG b�-㏕"LTAR�M_��cL�� σQ�N�<��METPUI�ǂ����)NDSP_CMNTh���|�N  d�.��ς��ҟܔ|�POSC�F����PSTOoL 1e'�4@�<#�
5�́5�E� S�1�S�U�g������� ߯��ӯ���	�K�-��?���c�u�����|�S�ING_CHK � ��;�ODAQ�,�f��Ç��DE�V 	L�	M�C:!�HSIZE�h��-��TASK� %6�%$12�3456789 ��Ϡ��TRIG �1g�+ l6�% ���ǃ�����8�p��YP[� ��EM_�INF 1h3�� `)�AT&FV0E0�"ߙ�)��E0V�1&A3&B1&�D2&S0&C1�S0=��)ATZ������H�����A���AI�q�,��|���� ���ߵ� ����J���n������ W�����������"�� ��X��/����e� �����0�T ;x�=�as� �/�,/c=/b/ �/A/�/�/�/�/�� ?���^?p?#/�? �/�?s?}/�?�?O�? 6OHO�/lO?1?C?U? �Oy?�O�O3O _�?D_��OU_z_a_�_�ON�ITOR��G ?�5�   	EOXEC1Ƀ�R2�X3�X4�X5�X���VU7�X8�X9Ƀ�R hBLd�RLd�RLd�RLd 
bLdbLd"bLd.bLdP:bLdFbLc2Sh2_hU2kh2wh2�h2�hU2�h2�h2�h2�h�3Sh3_h3�R�R�_GRP_SV �1in���(ͅ��
�3�8��r��ۯ_MOx�_D�=R^��PL_NA_ME !6��p��!Defau�lt Perso�nality (�from FD)� �RR2eq 1�j)TUX)TX9��q��X dϏ8� J�\�n���������ȏ ڏ����"�4�F�X� j�|������2'�П �����*�<�N�`�r��<��������ү �����,�>�P�b�: �Rdr 1o�y �{\�, �3����� @D� M ��?�����?�<���A'�6�����;�	lʲ	 ��x�J����� �< �"��� �(pK���K ��K=*��J���J���JV���Z��ƌ��rτ́p@j��@T;f����f��ұ]�l��Ik��p������������b��3���o�  �
`�>�����bϸ�z��;꜐r�Jm��
� B�H�˱]Ӂt��q�	� p� W P�pQ�p��p|  Ъ�g����c�	'� � ���I� � � ����:����
�È=����"�s��	�ВI  �n @B� cΤ�\��ۤ��tq��y߁rN���  '������@2�@�����/��C��C�C�@ �C������
S�A�W�@<�PΕR�
h�B�b�A��j�����:��Dz۩��߹������j��( �� -��C���0'�7�����q�Y������ �?�f�f ��gy �����q+qt��
>+�  PƱj�(����7	�x��|�?�����xZ�p<
6b<�߈;܍�<��ê<� <G�&Jσ�AI��ɳ+���?fff�?I�?&�k�@��.��J<?�`�q�.�˴f� ��/��5/����j/ U/�/y/�/�/�/�/�/`?�/0?q��F� ?l??�?/�?+)�?��?�E�� E�~I�G+� F� �?)O�?9O_OJO�OnO,�Of�BL޳B�?_ h�.��O�O��%_�OL_ �?m_�?�__�_�_�_<�_�
�h�Îg>��_Co�_go0Rodo�o�GA�ds��q�C�o�o�o|��Ƀ�$]Hq��6�D��pC���pCCHmZZ7t���6q��q��ܶN'�3A��A�AR1A�O�^?�$�?��K�0±
=�ç>����3�W
=�#�W���e��9������{����<���(�B��u��=B0�������	�L��H�F�G����G��H��U`E���C��+���I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3� l�W���{�������� ՟���2��V�A�z� ��w�����ԯ����� ���R�=�v�a��� ���������߿�� <�'�`�Kτ�oρϺ� ���������&��J� \�G߀�kߤߏ��߳� ������"��F�1�j� U��y��������� ���0��T�?�Q���:�(�1��3/E������5��x����q3�8���<��q4Mgs�&IB+2D�a?���{�^^	�������uP2P7Q4_A��`M0bt��R�������/   �/�b/P/�/t/ �/ *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?�?�?O 2 wF�$�vGb�/��A��@�a�`�qC���C@�o�O2���OF�� DzH@��� F�P D���O�O�ys<O!_3_�E_W_i_s?��ͫ@@pZ.t2�2!2~
 p_�_�_�_	oo-o ?oQocouo�o�o�o�o���Q ��+���1��$MSKCFMAP  �5� �6�Q�Q"~�cONREoL  
q�3�bEXCFEN�B?w
s1uXqFN�C_QtJOGOV�LIM?wdIpMrd��bKEY?w�u��bRUN�|�u��bSFSPDTY��avJu3sSIGN|?QtT1MOT��Nq�b_CE_G�RP 1p�5s\r���j�����T ��⏙������<�� `��U���M���̟�� 🧟�&�ݟJ��C� ��7�������گ��������4�V�`TCO�M_CFG 1qB}�Vp�����
P�__ARC_\r
�jyUAP_CPL���ntNOCHEC�K ?{ 	r��1�C�U� g�yϋϝϯ����������	��({NO_WAIT_L�	uM��NTX�r{�[�m�_ERRY�2sy3� &����߄��r�c� ��T�_MO��t��, �#�$�k�3�PA�RAM��u{���V[��!�u?�� �=9@345678901��&���E� W�3�c�����{������� ����=��UM_RSPA�CE �Vv��$?ODRDSP����jxOFFSET_�CARTܿ�DI�S��PEN_FILE� �q��c֮��OPTION_I�O��PWORK� v_�ms  �P(�R�Q
�j.j	 ��Hj&6$�� RG_DSBOL  �5Js�\���RIENTT5O>p9!C��Pq�fA� UT_SIM�_D
r�b� V~� LCT ww��bc��U)+$_PEsXE�d&RATp Тvju�p��2X�j)TUX)TX�##X d-�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	OO-O?O�H2�/oO�O �O�O�O�O�O�O�O_]�<^O;_M___q_�_ �_�_�_�_�_�_o���X�OU[�o(ҿ�(���$>o�, ��Ip~B` @D�  Ua?�[cAa?��]a]��DWcUa쪋l;��	lmb�`�xoJ�`�������a�< ���`� ��b, H�(��H3k7H�SM5G�22G���Gp
��
�!��'|, C%R�>�>q�Gsua|T�3���  �4spBpyr  ]o��*SB_���{�j]��t�q� ��rna �,����6  ���PQ�|�N�M�,k�!�	'�� � ��I�� �  �=�%�=��ͭ����ba	���I  ?�n @��~���p����� �9N	 W�  '!o�t:q�pC	 C�@@s�Bq�|��� m�
��!�h@ߐ�nH����Z�B	 �A���p� �-�qbz�P��t�_�������( �� -��恊�n��ڥ[A]Ѻ�b4�'!���(p �?�ff � ��
����OZ�DR��8��z���>΁'  Pia��(�ವ�@���ک�a�c�dF#?�����x����<�
6b<߈;�܍�<�ê<� <�&�o&�)�A�lcΐI�*��?fff?�?&�c���@�.u?J<?�`��Y ђ^�nd��]e��[g�� Gǡd<����1��U� @�y�dߝ߯ߚ����� ��	���-������&����"�E�� E�~�G+� Fþ� ����������&��PJ�5��bB��AT� 8�ђ��0�6���>��� J�n�7��[m<�0��h��1��>�M�I
0�@��A�[���C-�)��?���� /�Y�Ē��Jp��vav`CH/������}!�@I�Y�'�3�A�A�AR1�AO�^?�$��?����±
�=ç>�����3�W
=�#�\���+e��ܒ������{����<���.(�B��u��=B�0�������	�*H�F�G����G��H��U`E���C��+�-I#��I��HD��F��E��R�C�j=U>
�I��@H�!�H�( E<YD0/�?�?�?�? �?O�?3OOWOBOTO �OxO�O�O�O�O�O�O _/__S_>_w_b_�_ �_�_�_�_�_�_oo =o(oaoLo�o�o�o�o �o�o�o�o'$ ]H�l���� ���#��G�2�k� V���z���ŏ���ԏ ���1��U�g�R��� v�����ӟ�������t-��(���������a�����Q�c�,!3�8�x}���,!4Mgs�����ɢIB+կ篴a���{�� �A�/�e�S���w��%P!�P��������7��ӯ�ϑ�R�9�Kτ�oχϓϥ�  ���χ����)� �M����������{��ߛ���ߒߤ���8����  )�G��q�_���2 �F�$�&Gb����n�[ZjM!C�s�@j/�A�S���F� Dz���� F�P D�!�W����)������������x?��W�@@
9�E�E��E��
 v���� ���*<N�`�*P ���˨��1��$PAR�AM_MENU �?-���  DE�FPULSEl�	WAITTMO{UT�RCV�� SHELL�_WRK.$CU�R_STYL��,OPT�/P�TB./("C�R_DECSN���, y/�/�/�/�/�/�/? 	??-?V?Q?c?u?�?��USE_PRO/G %�%�?�?.�3CCR������7_HOST �!�!�44O�:T ̰�?PCO)ARC�O>�;_TIME�XB�  �GDE�BUGV@��3GI�NP_FLMSKĵO�IT`��O�EPG�AP �L��#[CyH�O�HTYPE����?�?�_�_�_ �_�_oo'o9obo]o oo�o�o�o�o�o�o�o �o:5GY�} ����������1�Z��EWORD� ?	7]	R}S`�	PNS��$��JOE!>��TEs@WVTRACECTL 1x-�� ���Ӱ��ɆDT �Qy-���Do � ��,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�T� (�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_j��_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�� �&�8�J�\�n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�_����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv��������//"#�$PG�TRACELEN�  #!  �_�" �8&�_UP z����g!o S!�h 8!_CFG �{g%Q#"!x!��$J �" |"DEF�SPD |�,l!!J �8 IN �TRL }�-�" 8�(IPE_C�ONFI� ~g%O�g!�$�$\�"8 LID�#�-�74GRP 1��7Q!�#!A ����&ff"!A�+33D�� D�]� CÀ A)@+6�!�" d�$�9��9*1*0� 	 �+9�-+6�? ´	C�?�;B@3AO�?�OIO3OmO"!>�T?�
5�O�O�N��O =��=#�
�O_�O_J_5_ n_Y_�O}_�_y_�_�_�_  Dzco" 
oBo�_Roxoco�o �o�o�o�o�o�o�>)bM��;
�V7.10bet�a1�$  �A�E�rӻ��A " �p?!G�^�q>���r��0��q�ͻqBQ��qA\�p�q�4�q*�p�"�BȔ2�D�V�h�w��p�?�?)2{ȏw�׏� ��4��1�j�U���y� ����֟������0� �T�?�x�c������� ү����!o�,�ۯP� ;�M���q�����ο�� �ݿ�(��L�7�p�x+9��sF@ �� �ͷϥ�g%������ +�!6I�[߆������� �ߠ���������!�� E�0�B�{�f����� ���������A�,� e�P���t��������� ���=(aL ^������ �'9$]�Ϛ��� ��������/<� 5/`�r߄ߖߏ/>�/ �/�/�/�/?�/1?? U?@?R?�?v?�?�?�? �?�?�?O-OOQO<O uO`O�O�O�O�O���O _�O)__M_8_q_\_ n_�_�_�_�_�_�_o �_7oIot���o�o ���o�o�o(/!L/ ^/p/�/{*o��� ������A�,� e�P�b���������� Ώ��+�=�(�a�L� ��p������Oߟ񟠟 � �9�$�]�H���l� ~�����ۯƯ���#� No`oro�on��o�o�o �oԿ���8J\ ng����vϯϚ��� ����	���-��Q�<� u�`�r߫ߖ��ߺ��� ����;�M�8�q�\� ��������z������ %��I�4�m�X���|� ����������:�L� ^���Z�������� ���$�6�H�S wb����� ��//=/(/a/L/ �/p/�/�/�/�/�/? �/'??K?]?H?�?�� �?�?f?�?�?�?O�? 5O OYODO}OhO�O�O �O�O�O�O&8J4_ F_����_�_��_ �_"4-o�O*oco No�oro�o�o�o�o�o �o)M8q\ �������� �7�"�[�m��?���� R�Ǐ���֏�!�� E�0�i�T���x����� ���_$_V_ �2�l_�~_�_�����R�$P�LID_KNOW�_M  �T������SV� ��U͠�U��
��.� ǟR�=�O�����mӣ�M_GRP 1�T�!`0u��T@ٰ)o�ҵ�
���P зj��`���!�J� _�W�i�{ύϟϱ���`������߱�MR��Ņ��T��s�w�  s��ߠ޴߯߅��ߩ� ������A���'�� ����������� ��=���#����������}������S��ST^��1 1��U# ����0�_ A  .��,>Pb�� ������3 (iL^p���(��2*��'�<-/3/)/;/M/4f/x/�/�/�5�/�/�/�/6 ??(?:?7S?e?w?�?8�?�?�?�?~MAD  d�#`PARN_UM  w�\%OSCH?J ME�
�G`A�Iͣ�EUP�D`OrE
a�OT_CMP_��B@�P@�'˥TER_C;HK'U��˪?R�$_6[RSl�¯��_#MOA@�_�U_�_RE�_RES_G � �>�oo8o+o\o Oo�oso�o�o�o�o�o@�o�o�W �\�_ %�Ue Baf�S�  ����S0��� �SR0��#��S�0>� ]�b��S�0}������R�V 1�����rB@�c]��t�(@�c\����D@�c[�$���RTHR_INRl�DA��z˥d,�MASS9�� ZM�MN8�k�M�ON_QUEUE� ���˦��x� URDNPUbQN{�P[��END���_ڙ�EXE�ڕ�@BE��ʟ��OPTIO�Ǘ�[��PROGR�AM %��%�ۏ�O��TASK�_IAD0�OCFG� ���tO��ŠD�ATA���Ϋ@��27�>�P�b�t� ��,�����ɿۿ������#�5�G���INFOUӌ�������� �Ͽ���������+� =�O�a�s߅ߗߩ߻�@�������^�jč�� yġ?PDIT� �ίc���WE�RFL
��
RG�ADJ �n�A	����?����@���?IORITY{�QV}���MPDSPH������Uz����O�TOEy�1�R�� (!AF4�E��P]���!tc�ph���!ud|��!icm���ݏ6�XY_ȡ��R��ۡ)� *0+/ ۠�W :F�j���� ��%7[B��*��PORTT#�BC۠�����_CARTREP�
�R� SKSTA�z��ZSSAV����n�	2500H863���r�$!�U�R����q��n�}/�/�'� URGeE�B��rYWF� #DO{�rUVWV��$��A�WRUP_DELAY �R�>�$R_HOTk���%O]?�$R_NORMALk�L?�?p6SEMI?�?�?3A_QSKIP!�n�;l#x 	1/+O + OROdOvO9Hn��O �G�O�O�O�O�O_�O _D_V_h_._�_z_�_ �_�_�_�_
o�_.o@o Roovodo�o�o�o�o �o�o�o*<L�r`���n��$�RCVTM���]��pDCR!�L�ЈqCl�fC���C��>?��A�>:��<�l��4M�b�����O
��n��������{�4Oi��O �<
6b<���;܍�>u.��?!<�&{�b�ˏݏ��8��� ��,�>�P�b�t��� ������Ο���ݟ� �:�%�7�p�S����� �ʯܯ� ��$�6� H�Z�l�~�������ƿ ���տ���2�D�'� h�zϽ��ϰ������� ��
��.�@�R�d�O� �ߚ߅߾ߩ������ ���<�N��r��� �����������&� 8�#�\�G�����}��� ��������S�4F Xj|����� ����0T? x�u����' //,/>/P/b/t/�/ �/�/�/�/�/�?�/ (??L?7?p?�?e?�? �?��?�? OO$O6O HOZOlO~O�O�O�?�? �O�O�O�O __D_V_ 9_z_�_�?�_�_�_�_ �_
oo.o@oRodovo��X�qGN_ATC� 1�� �AT&FV0E�0�kATDP�/6/9/2/9��hATA�n,�AT%G1%�B960�i+�++�o,�aH,��qIO_TYPE'  �u�sn_�o�REFPOS1 �1�P{ x�o�Xh_�d_�� ���K�6�o�
����.���R����{{2 1�P{���؏V��ԏz����q3 1� �$�6�p��ٟ���S4 1�����˟����n���%�S5 1�<�N�`�����|<���S6 1�ѯ����/�����ѿO�S7 1�f�x���Ŀ�B�-�f��S8 1�����Y��������y�SMASK 1�P  
9�G��'XNOM���a~���ӁqMOTE  �h�~t��_CFG �������рrPL_RANG�ћQ���POWER ��e��SM_D�RYPRG %�i�%��J��TAR�T �
�X�UME_PRO'�9���~t_EXEC_E�NB  �e��GSPD������c��gTDB���RM�.�MT_!�T����`OBOT_N�AME i����iOB_ORD_NUM ?
��\qH863  �T���������bPC_TI�MEOUT�� xޔ`S232��1���k LTE�ACH PENDcAN �ǅ�}����`Maint�enance CGons�R}�m
"{~�dKCL/Cg�ȔZ ��n� No Use}p�	��*NPO�\�х���(oCH_L��������	�mMAVGAIL��{������SPACE1 ;2��| d�� (>��&���p��~M,8�?�e p/eT/�/�/�/�/�W //,/>/�/b/�/v? �?Z?�/�?�9�e�a�= ??,?>?�?b?�?vO �OZO�?�O�O�Os�2�/O*O<O�O `O�O�_�_u_�_�_�_�_[3_#_5_G_Y_ o}_�_�o�o�o�o�o[4.o@oRodo vo$�o�o����"�	�7�[5K]o ��A����	�̏ �?�&�T�[6h�z� ������^�ԏ���&�@�;�\�C�q�[7�� ������͟{���"��C��X�y�`���[8 ����Ưدꯘ��0� ?�`�#�uϖ�}ϫ�[�G �i� t�ϋ
G� �� ��$�6�H�Z�l�~ߐ� �8 ǳ�����߈���d(���M�_�q� �����������? ���2�%�7�e�w��� ���������������� �!�RE�W���� �������?Q `�� @0��ߖrz	�V_����� 
/L/^/|/2/d/�/�/ �/�/�/�/?�/�/�/ *?l?~?�?R?�?�?�?��?�?�?�?2O�?
���O[_MODE�  �˝IS E���vO,*���O-_��	M_v_#d�CWORK_ADޭM�P%aR  ��ϰ�P{_�P_INTVAL�@�����JR_OPT�ION�V �E�BpVAT_GRPw 2����G(y_Ho �e_ vo�o�oYo�o�o�o�o �o*<�bOoND pw������ 	���?�Q�c�u��� ��/���ϏᏣ���� )�;���_�q������� ��O�ɟ���՟7� I�[�m�/�������ǯ ٯ믁��!�3���C� i�{���O���ÿտ� ��ϡ�/�A�S�e�'� �ϛϭ�oρ������ �+�=���a�s߅�G� �߻����ߡ���'� 9�K�]��߁���� y����������5�G��Y��E�$SCAN�_TIM�AYue�w�R �(�#�((�<0.aWaPaP
T�q>��Q��o������OO"2/��:	d/JaR��WY��^����^R^	r  P~��� �  8�P�	�D��GYk }�������8�Qp/@/�R//)P;�o�\T��Qpg-�t�_DiKT��[  � lv%�� �����/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O WW�#�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ olO~Od+No`oro�o �o�o�o�o�o�o &8J\n���p���u�  0�" 0g�/�-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q����� $o��˟ݟ���%� 7�I�[�m�������� ǯٯ����!�3�E� ����Do��������ҿ �����,�>�P�b� tφϘϪϼ���������w
�  58�J� \�n߀ߒߜկ����� ����	��-�?�Q�c��u����� � ��-����� �2�D��V�h�z�������������������&� ��%	12�345678�"W 	��/� @`r������ ��(:L^ p�������  //$/6/H/Z/l/~/ ��/�/�/�/�/�/?  ?2?D?V?h?�/�?�? �?�?�?�?�?
OO.O @Oo?dOvO�O�O�O�O �O�O�O__*_YON_ `_r_�_�_�_�_�_�_ �_ooC_8oJo\ono �o�o�o�o�o�o�oo "4FXj|� ���������	��s3�E�W�{��Cz  Bp�� /  ��2���z��$SCR_GR�P 1�(�U8�(�\x�^ @  �	!�	 ?׃� ��"�$� ��-��p+��R�w����CD~�����#�����O���M-10�iA 89099�05 Ŗ5 M61�C >4��Jׁ

� ���0� ����#�1�	"�z��������¯Ҭ ���c���O�8� J�������!������ֿ��B�y�Ɛ�������A��$� C @��<� �R�?�Єd���Hy�u�O���F?@ F�`�§� ʿ�϶�������%�� I�4�m��<�l߃��ߧ߹�B���\�� ��1��U�@�R��v� ����������� ;���*<=�
F���x?�d�<�>m����@�:��� BȆ��ЗЙ���E�L_DEFAUL�T  �����B�MI�POWERFL � �$1 WF�DO $��E�RVENT 1������"�pL�!DUM_EI�P��8��j!AF_INE �=�O!FT���r!��4 ���[!RPC_M'AIN\>�J�NnVISw=����!TP�PU���	d�?/!
P�MON_PROX	Y@/�e./�/"Y/�fz/�/!RD�M_SRV�/�	g�/#?!R C?�Yh?o?!
pM�/�i^?�?!RL�SYNC�?8�8|�?O!ROS�.L�4�?SO"wO�# DOVO�O�O�O�O�O_ �O1_�OU__._@_�_ d_v_�_�_�_�_o�_�?oocoiICE_�KL ?%y �(%SVCPRG1ho8��e���o�m3�o�o�`4 �`5(-�`6PU�`�7x}�`���l9��{�d:?��a�o ��a�oE��a�om��a ���aB���aj� �a���a�5��a� ]��a����a3����a [�՟�a�����a��%� �aӏM��a��u��a#� ���aK�ů�as���a ��mob�`�o�`8�}� w�������ɿ���ؿ ���5�G�2�k�VϏ� zϳϞ���������� 1��U�@�y�dߝ߯� ���߾�������?� *�Q�u�`����� �������;�&�_� J���n������������sj_DEV �y	�MC:�P�_OU�T",RE�C 1�Z� d {  	 	�������
 �PJ��%6 (�&��[w�,�n*  T - %�- �A�- c|� P�����// B/0/f/x/Z/�/�/�/ �/�/�/�/?�/?P? >?t?b?�?�?�?�?�? �?�?OOOLO:OpO �OdO�O�O�O�O�O�O �O$__H_6_X_~_l_ �_�_�_�_�_�_�_ o oDo2oTozo\o�o�o �o�o�o�o�o. R@vd���� },����4�"� X�F�|���p�����֏ ď����0��@�f� T���x�����ҟ�Ɵ ���,��<�b�P��� h�z������ί�� (�:��^�L�n�p��� ����ܿ�п� �6� $�Z�H�jϐ�rϴϢ� ���������2�D�&� h�Vߌ�z߰ߞ����� ������
�@�.�d�R�x��ZjV 1�w� P�m��	>�   <��
TYPEV�FZN_CFG ;��d�7�GRP 1y�A�c ,B� �A� D;� B}���  B4�RB21H�ELL:�(
ƶ X����%RSR����E0 iT�x���� ��/Sew��  ��%@w�����#�1�������2#�d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he��_ &_8_J_\_��_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}6copy f�rs:order�fil.dat �virt:\te�mp\=>192�.168.4�P4?6:3020>_�_��_o}.�V*.d��_�^�_`oro�oe
�xyzrate 61 +o=oOo�o�oe�g�o�a�o�o�cu�b4�Rmd�:prgst�`.dg�o�]U��
�� }3�ucons'log�� �e�w����io�<�N��ߏ��f2�uerrall.ls����_Տf�x��� }9��_�Xmpback�<�R���
� }0J�tb(`*��ǟ џ�b�t���c�_�_=�8144 W������ o��˩ϯ`�r����o �o;�M�޿��' д��ҿc�uχϚ��� 5�ͧ�������"���@̨��b�t߆ߙtx��:\)ߪ�;�S�U���\��
� }5��a�� ��H���i�{�Ϡϲ� @�V������߹�B� ��e�w�����/�<��� ��������P�a s����3����� �(��L�]o� ����9����� $�HY/k/}/���� +/=/O/�/�/?�)�6788 �/�/c? u?�?��567�?�? �?"�?58�?bOtO��O���?��81976 WO�O�O�O��O�I �O`_r_�_�/��;_M_ �_�_o?'?�T�_�_ couo�o�?�?5O�G�o �o�oO"O�o�H�ob t���/�/:dV�`��/��6 � g�y����o�o9T� ��	���@ҏc�u�������$SNPX�_ASG 1��������� P 0 '�%R[1]@g1.1����?���%֟��&�	��\� ?�f���u�������� ϯ��"��F�)�;�|� _�������ֿ��˿� ��B�%�f�I�[Ϝ� Ϧ��ϵ�������,� �6�b�E߆�i�{߼� ������������L� /�V��e������ �������6��+�l� O�v������������� ��2V9K� o������ �&R5vYk� ����/��</ /F/r/U/�/y/�/�/ �/�/?�/&?	??\? ??f?�?u?�?�?�?�? �?�?"OOFO)O;O|O _O�O�O�O�O�O�O_ �O_B_%_f_I_[_�_ _�_�_�_�_�_�_,o o6oboEo�oio{o�o �o�o�o�o�oL /V�e���� ����6��+�l��O�v�������PAR�AM ������ �	��P�����OFT�_KB_CFG � ヱ���PIN_SIM  ����C�U�g�����R�VQSTP_DS�B,�򂣟����S�R �/�� &�  ULTIR�OBOTTASK������TOP_�ON_ERR  ����PTN� /�@��A	�RING_�PRM� ��V�DT_GRP 1y�ˉ�  	�� ����������Я��� ��*�Q�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߣߠ߲��� ��������0�B�i� f�x���������� ���/�,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZ�~��� ����/ /G/D/ V/h/z/�/�/�/�/�/ �/?
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8___\_��VPRG_COUNT���@���RENB�U��UM�S��__U�PD 1�/�8  
s_�oo*o SoNo`oro�o�o�o�o �o�o�o+&8J sn������ ���"�K�F�X�j� ��������ۏ֏��� #��0�B�k�f�x��� ������ҟ������ C�>�P�b����������ӯί�����UY?SDEBUG�P�P��)�d�YH�SP_�PASS�UB?~Z�LOG ��U+�S)�#�0��  ��Q)�
M�C:\��6���_M�PC���U���Q�ñ8� �Q�SAV �����ǲ&��ηSV;�TE�M_TIME 1]��[ (m�4&��1:�}YT1SV�GUNS�P�U'��U���ASK_OPTION�P�U�Q��Q��BCCFGg ��[u� n�A�a�`a�gZo� �߃ߕ��߹������ �:�%�^�p�[��� ������� �����6� !�Z�E�~�i���������&�������&8 ��nY�}�?� �ԫ ��( L:p^���� ���/ /6/$/F/ l/Z/�/~/�/�/�/�/ �/�/�/2?8 F?X? v?�?�??�?�?�?�? �?O*O<O
O`ONO�O rO�O�O�O�O�O_�O &__J_8_n_\_~_�_ �_�_�_�_�_o�_ o "o4ojoXo�oD?�o�o �o�o�oxo.T Bx��j��� �����,�b�P� ��t�����Ώ��ޏ� �(��L�:�p�^��� ����ʟ��o�� 6�H�Z�؟~�l����� ��د���ʯ ��D� 2�h�V�x�z���¿�� �Կ
���.��>�d� Rψ�vϬϚ��Ͼ��� ����*��N��f�x� �ߨߺ�8�������� �8�J�\�*��n�� �����������"�� F�4�j�X���|����� ��������0@ BT�x�d��� ��>,Nt b������/ �(//8/:/L/�/p/ �/�/�/�/�/�/�/$? ?H?6?l?Z?�?~?�? �?�?�?�?O�&O8O VOhOzO�?�O�O�O�O �O�O
__�O@_._d_ R_�_v_�_�_�_�_�_ o�_*ooNo<o^o�o ro�o�o�o�o�o�o  J8n$O�� ���X���4��"�X�B�v��$TB�CSG_GRP �2�B���  �v� 
 ?�  ������ ׏�������1��U��g�z���ƈ�d�, ���?v�	 �HC��d�>�����e�CL  Bጙ�Пܘ������\)��Y  3A�ܟ$�B�g�B�#Bl�i�X�ɼ���>X��  D	J���r�����C����үܬ���D�@v�=�W� j�}�H�Z���ſ���������v�	�V3.00��	�m61c�	�*X�P�u�g�p�>�d��v�(:�� ���p͟�  O�����p�����z�JCFoG �B���Y ��������9��=��=�c� q�K�qߗ߂߻ߦ��� �����'��$�]�H� ��l���������� ��#��G�2�k�V��� z����������� ���p*<N���l �������# 5GY}h�� ��v�b��>�//  /V/D/z/h/�/�/�/ �/�/�/�/?
?@?.? d?R?t?v?�?�?�?�? �?O�?*OO:O`ONO �OrO�O�O��O�O�O _&__J_8_n_\_�_ �_�_�_�_�_�_�_�_ oFo4ojo|o�o�oZo �o�o�o�o�o�oB 0fT�x��� ����,��P�>� `�b�t�����Ώ��� ����&�L��Od�v� ��2�����ȟʟܟ�  �6�$�Z�l�~���N� ����دƯ�� �2� �B�h�V���z����� Կ¿����.��R� @�v�dϚψϪ��Ͼ� ������<�*�L�N� `ߖ߄ߺߨ����ߚ� ������\�J��n� ����������"� ��2�X�F�|�j����� ����������. TBxf���� ���>,b P�t����� /�(//8/:/L/�/ �ߚ/�/�/h/�/�/�/ $??H?6?l?Z?�?�? �?�?�?�?�?O�?O DOVOhO"O4O�O�O�O �O�O�O
_�O_@_._ d_R_�_v_�_�_�_�_ �_o�_*ooNo<oro `o�o�o�o�o�o�o�o &�/>P�/� �������� 4�F�X��(���|��� ��֏����Ə0�� @�B�T���x�����ҟ ������,��P�>� t�b������������ ���:�(�^�L�n� ������2d����� ̿�$�Z�H�~�lϢ� ���������Ϻ� �� 0�2�D�zߌߞ߰�j� ���������
�,�.� @�v�d������� ������<�*�`�N� ��r����������� ��&J\�t� �B������ F4j|��^�����/�  92 6# 6&J/�6"�$TBJOP_GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� =�6$ @2 �"	 �C�� �&b  Cق'�!�!�>���
559>��0+1�33=�CL� fff}?+0?�ffB� �J1�%Y?d7�.��/>w��2\)?�0�5���;���hCY� �  @�� �!B�  A��P?�?�3EC�  �D�!�,�0*BO�ߦ?�3JB��
:_���Bl�0��0��$�1�?O6!Aəg�AДC�1D�G�6�=q�E6O0��p��B�Q�;��A�� ٙ�@L3D	�@�@_x_�O�O>B�\JU��OHH�1ts�A@�33@?1� C��� �@�_�_&_8_>�#�D�UV_0�LP�Q�30<{�zR� @ �0�V�P!o3o�_<oRi foPo^o�o�o�oRo�o �o�o�oM(�ol@�p~��p4�6&��q5	V3.�00�#m61c�$*(��$1!6�A�� Eo�E���E��E��F��F�!�F8��F�T�Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G�,IR�CH`��C�dTDU�?�D��D��D�E(!/E\��E��E�h��E�ME��s�F`F+'\�FD��F`=�F}'�F���F�[
F����F��M;S@;Q���|8�`rz(@/&�8�6&<��1��w�^$ESTPARS  *({ _#�HR��ABLE K1�p+Z�6#|��Q� � 1�|�|�P|�5'=!|�	|�
|�Q|�˕6!|�|�u|���RDI��z!ʟܟ� ��$���O������¯ԯ�$����S��x# V��� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����U-����ĜP� 9�K�]�o��-�?�Q��c�u���6�NUM [ �z!� �>  Ȑ����_CFG �����!�@b IMEBF_�TT����x#��a�V�ER��b�w�a�R� 1�p+
 ($3�6"1 ��  6! ���������� �9�$� :�H�Z�l�~����������������^$��_���@x�
b MI__CHANm� x�} kDBGLV;0�o�x�a!n ETHERAD ?�� �y�$"��\&n ROUT���!p*!*�SNMASK�x#�255.h�f�x^$OOLOFS�_DI��[ՠ	O�RQCTRL �p+;/���/+/ =/O/a/s/�/�/�/�/��/��/�/�/!?��PE_DETAI���PON_SVO�FF�33P_MOON �H�v�2-9�STRTCHK ����42VT?COMPATa8��24:0FPROG �%�%MUL�TIROBOTT�O!O06�PLAY���L:_INST_�MP GL7YDUqS���?�2LCK�L�PKQUICKMExt �O�2SCRE�@��
tps���2�A�@�I��@_�Y���9�	SR_G�RP 1�� ���\�l_zZ�g_�_�_�_�_�_�^� ^�oj�Q'ODo/oho Se��oo�o�o�o�o �o�o!WE{�i������	�1234567���!���X�E1��V[
 �}ip�nl/a�gen.htmno���������ȏ~�Panel setup̌}�?��0�B�T�f� ��񏞟��ԟ ���o����@�R�d� v������#�Я��� ��*���ϯůr��� ������̿C��g�� &�8�J�\�n������ ����������uϣϙ� F�X�j�|ߎߠ���� ;�������0�B�߾*NUALRMb@G7 ?�� [�� ����������� �� %�C�I�z�m�������~v�SEV  �����t�ECFG� Ձ=]/BaA�$   B�/D
 ��/C�Wi{ �������h PRց; �(To\o�I�6?K0(%����0��� ��//;/&/L/q/�\/�/�/�/l�D ؅Q�/I_�@HI�ST 1ׁ9  �(  ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,1 Ec0p?�?�?�?�/C�� >?P=962n?�?
OO.O�?�?�136c?|O�O�O�O AOSO�?�O__0_�O �O_Lu_�_�_�_:_�/ �_�_oo)o;o�__o qo�o�o�o�oHo�o�o %7I~��a81 �ou������o ���)�;�M��q� ��������ˏZ�l�� �%�7�I�[����� ����ǟٟh����!� 3�E�W���������� ïկ�v���/�A� S�e�Pb������ѿ ������+�=�O�a� s�ϗϩϻ������� ߒ�'�9�K�]�o߁� ߥ߷��������ߎ� #�5�G�Y�k�}��� �������������1� C�U�g�y���v����� ������	�?Q cu��(��� �)�M_q ���6���/ /%/�I/[/m//�/ �/�/D/�/�/�/?!? 3?�/W?i?{?�?�?�? �����?�?OO/OAO D?eOwO�O�O�O�ONO `O�O__+_=_O_�O s_�_�_�_�_�_\_�_ oo'o9oKo�_�_�o �o�o�o�o�ojo�o #5GY�o}������?��$U�I_PANEDA�TA 1������  	�}�0�B�T�f�x��� )����mt �ۏ����#�5��� Y�@�}���v�����ן �������1��U�g��N������ �1 ��Ïȯگ����"� u�F���X�|������� Ŀֿ=������0� T�;�x�_ϜϮϕ���@�������,ߟ�M� �j�o߁ߓߥ߷��� ���`��#�5�G�Y� k��ߏ�������� ������C�*�g�y� `���������F�X�	 -?Qc����� �����~ ;"_F��|� ����/�7/I/ 0/m/�����/�/�/�/ �/�/P/!?3?�W?i? {?�?�?�??�?�?�? O�?/OOSOeOLO�O pO�O�O�O�O�O_z/ �/J?O_a_s_�_�_�_ �O�_@?�_oo'o9o Ko�_oo�oho�o�o�o �o�o�o�o#
GY @}d��&_8_� ���1�C��g��_ ��������ӏ���^� ��?�&�c�u�\��� ����ϟ���ڟ�)� �M����������� ˯ݯ0�����7�I� [�m����������ٿ �ҿ���3�E�,�i� Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#����� �� ��$�6��Z�A� ~�e�w�������� ���2��V�h�O������v�p��$UI_�PANELINK� 1�v��  �  ���}1234567890����	 -?G ���o� ����a�� #5G�	����p&���  R�� ���Z��$/6/ H/Z/l/~//�/�/�/ �/�/�/�/
?2?D?V? h?z??$?�?�?�?�? �?
O�?.O@OROdOvO �O O�O�O�O�O�O_ �O�O<_N_`_r_�_�_�0,���_�X�_�_ �_ o2ooVohoKo�o oo�o�o�o�o�o�o ��,>r}���� �������� /�A�S�e�w������ ��я���tv�z�� ��=�O�a�s����� ��0S��ӟ���	�� -���Q�c�u������� :�ϯ����)��� M�_�q���������H� ݿ���%�7�ƿ[� m�ϑϣϵ�D����� ���!�3�Eߴ_i�{� 
�߂����߸���� ��/��S�e�H��� ~��R~'�'�a�� :�L�^�p��������� ������ ��6H Zl~���#�5� �� 2D��h z�����c� 
//./@/R/�v/�/ �/�/�/�/_/�/?? *?<?N?`?�/�?�?�? �?�?�?m?OO&O8O JO\O�?�O�O�O�O�O �O�O[�_��4_F_)_ j_|___�_�_�_�_�_ �_o�_0ooTofo�� �o��o��o�o�o ,>1bt�� ��K����(� :����{O������ ʏ܏�uO�$�6�H� Z�l���������Ɵ؟ ����� �2�D�V�h� z�	�����¯ԯ��� ���.�@�R�d�v��� �����п���ϕ� *�<�N�`�rτ��O�� ��Io���������8� J�-�n߀�cߤ߇��� �߽����o1�oX� �o|��������� ����0�B�T�f��� ������������S�e� w�,>Pbt�� '����� :L^p��#� ��� //$/�H/ Z/l/~/�/�/1/�/�/ �/�/? ?�/D?V?h? z?�?�?�???�?�?�? 
OO.O��ROdO�߈O kO�O�O�O�O�O�O_ �O<_N_1_r_�_g_�_�7OM�m�$U�I_QUICKM�EN  ���_AobRE�STORE 1��  �|��Rto�o�im�o�o�o�o�o :L^p�%�� ����o���� Z�l�~�����E�Ə؏ ���� �ÏD�V�h� z���7�������/��� 
��.�@��d�v��� ����O�Я����� ßͯ7�I���m����� ��̿޿����&�8� J��nπϒϤ϶�a� ������Y�"�4�F�X� j�ߎߠ߲������߀����0�B�T�gS�CRE`?#m�u1sco`�u2��3��4��5*��6��7��8��b�USERq�v��TLp���ks����4��U5��6��7��8���`NDO_CFG� �#k  n` �`PDATE ����No�nebSEUFR�AME  �T�A�n�RTOL_A�BRTy�l��EN�B����GRP 1��ci/aCz  A�����Q�� $6HRd��`�U�����MSK � �����Nv��%�U�%���bV�ISCAND_M;AX�I���FAIL_IMG�� �PݗP#��IMREGNUM�9
,[SIZ�n`��A�,VONOTMOU��@����2��a���a�����FR:\ � MC:\��\LOG�B@F� !�'/!+/O/��Uz MCyV�8#UD1r&�EX{+�S�PPOO64_��0'f�n6PO��L!Ib�*�#V���,�f@�'�/� =�	�(SZV�.�����'WAI�/S?TAT ����P!@/�?�?�:$�?�?���2DWP  ?��P G@+b=��� H�O�_JMPERR �1�#k
  �2�345678901dF�ψO{O�O�O�O �O�O_�O*__N_A_�S_�_
� MLOWpc>
 �_TI��=�'MPHA�SE  ��F�|�PSHIFT�k1 9�]@<�\ �Do�U#oIo�oYoko �o�o�o�o�o�o�o6 lCU�y� ���� ��	�V��-�e2����	V�SFT1�2	V:M�� �5�1G�� ���%A�  �B8̀̀�@ p�كӁ˂�у��z�ME@�?�{��!c>W&%�aM1��k��0�{ �$`0TDINEND��\�AO� �z����S���w��P���ϜRELE�Q��Y���~\�_ACTIV�x�:�R�A ��0e���e�:�RD� ����YBOX �X9�د�6��02����190.�0.�83�N�254��QF�	 �X�j��1��robot����   �p�૿�5pc ��̿�����7������-�f�ZABC�����,]@U��2ʿ�e� �ωϛϭϿ����� � ��V�=�z�a�s߰�E�Z��1�Ѧ