��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �P  �ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  �1�GPCU�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|GRG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"GSBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�H UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�H W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2FX�D�#
 d �$CARD_E�XIST4$FSSB_TYP~uAHKBD_S�B֒1AGN Gn �$SLOT_N�UMJQPREV�,DBU� g1G ;1_�EDIT1 �� 1G=� S<�0%$EP�O$OP�A�ETE_OKRU�S�P_CRQ�$;4�V� 0LACIw1�RAPk �1�x@ME@$D�V�Q�Pv�A{�oQL� OUzR A,mA�0�!� B� OLM_O�^eR�"�CAM_;1 �xr$ATTqR4NP� ANN�@�5IMG_HEI�GHQ�cWIDTMH4VT� �UU0F_ASPECQw$M�0EXP�v�@AX�f�CFT� X $GR�� � S�!�@B@N�FLI�`t� UI�RE 3dTuGITC�HC�`N� S�d_�L�`�C�"�`ED(lpE� J�4S�0� ��zsa�!ip;G0� � 
$WARNM�0f�!,P� �s��pNST� CORyN�"a1FLTR�u�TRAT� T�p H0ACCa1��8�{�ORI
`"S6={RT0_S�B�q�HG,I1 �[ Tp�"3I9�T�Y�D,P*2 �``w@� �!R*HD�cQJ* C��2��3��U4��5��6��7��U8��94�qO�$ <� $6xK3� 1w`O_M�@�C/ t � E#63NGP�ABA� �c���ZQ���`���@nr��� ��P�0����x�p�PzPb2�6����"J�_R��BC�J��3�JVP��tBS��}Aw؅�"�tP_*0OF�SzR @� RO1_K8���aIT�3��ONOM_�0�1ĥp34 ��T �� �$���AxP��K}EX �� �0g0I01��p��
$TFa��C$M�D3��TO�3�0U�� �� �H�w2�C1|�EΡg0�wE{vF�vF�40C�Pp@�a2 
P$�A`PU�3N1)#�dR*�AX�!sD�ETAI�3BUFpV��p@1 |�p�۶�pPIdT� PP[�MZ�Mg�Ͱj�}F[�SIMQSI �"0��A.�����lw' Tp|zM��P��B�FACTrbHPEW7�P1Ӡ��vv��MCd� ��$*1JB�p<�*1DECHښ�H��(�c�� � +PNS�_EMP��$GP���,P_��3�p�@Pܤ��TC��|r�� 0�s��b�0�� �B����!
���JR� ��S/EGFR��Iv �a�R�TkpN&S,�P�VF4��� &k�Bv�u�cu��a E�� !2��+�MQ��EчSIZ�3����T��P�����aRSINF�����kq��������LX������F�CRCMu�3CC lpG��p���O}���b��1�������2�V�D
xIC��C���r����0P��{� EV �zUF_��F�pNB
0�?������A�! �r�Rx���� V�lp�2��aR�t�,��g���]�Sx #�5�5"2��uA�R���`CX�$LG�p��B�1 `s�P�tB�aA�0{�У+0R���tME�`!BupCfrRA 3tAZ��h��pc�OT�FC�b�`�`FNp���1��ADI+�a%��b �{��p$�pSp�c�`aS�P��a,QMP6䒁`Y�3��M'�pUt��aU  $>�TITO1�S�S�!���$�"0�DBPX�WO��!��$cSK��2�DB��"�"@�PR8�� 
� ���# �>�q1$��$��+�L9$?(�V�R%@?R4C&_?�R4ENE��'�~?(�� RE�pY2(oH �OS��7#$L�3$$3RЯ�;3�MVOk_D@!V�ROScrr�w��S���CRIGGE�R2FPA�S��7�E�TURN0B�cMR-_��TUː[��0�EWM%���GN>`��RLA���Eݡy�P�&$P�"t�'�@4a��C�DϣV�DXQ��4�1��MVGO_AWAYR�MO#�aw!� C{S_)  `IS#� �� �s3S�AQ汯 4Rx�ZS W�AQ�p�@1UW��cT'NTV)�5RV
a�@��|c�éWƃ��JBx��x0��SAFEۥ��V_SV�bEXC�LUU�;��ON�L��cYg�~az�OyT�a{�HI_V? ���R, M�_ *Ȥ0� ��_z�2� ��"PSGO  +�rƐm@�A�c~b����w@��V�i�b�fA�NNUNx0�$�dI%DY�UABc�@Sp �i�a+ �j�f�!�p�OGIx2,��$1F�b�$ѐOT�@A� $DUMMAY��Ft��Ft±� |6U- ` !�HE�|s��~bc�B�@ SUFFI���4PCA�Gs5rCw6CqrMSWU�. 8!�KEYI��5�TM�1�s�qoA&�vINޱw��!, �/ D��HOST�P!4���<���`<�°<��p<�EM'����Z�� SBL� U}L��0  �	���E�� T�01� � $��9USAMPLо�/���決�$ I@갯 $SUBӄ��w0QSp�����#��SAV� ����c�S< 9�`�f�P$�0E!� YN�_B�#2 0�`D�I�d�pO|�m��#�$F�R_IC� �ENC2_Sd3  ��< 3�9���� cgp����!4�"��2�A��ޖ5���`ǻ�@�Q@K&D-!�a�AV�ER�q����DSP
���PC_�q��"��|�ܣ�VALU�3�HE�(�M�I�P)���OPPm ��TH�*��SH" T�/�Fb�;�d�����d ��q�16� H(rLL_DU ǀ�a�@��k���֠OT�"U�/����@@�NOAUTO7�0�$}�x�~�@sT��|�C͠��C� �2v�L�� 8/H *��L� � ��Բ@sv��`� �� � ����Xq��cq���q��T�q��7��8��9���0���1�1 �1�-�1:�1G�1T�1*a�1n�2|�2��U2 �2-�2:�2G�U2T�2a�2n�3|ʥ3�3� �3-�3�:�3G�3T�3a�3zn�4|­'�����9 <���z�ΓKI����H硵Ba�FEq@{@: ,<��&a? P_P�?��>�����E��@��r�RP��;�fp$TP�$�VARI����,�U�P2Q`< W�߃TD��g���`�������͠��BAC�"= T2����$)�,+r³�p IFI��p��H� q M�P"u�Fl@|``>t ;��46����ST����T��M ����0	 ��i���F����������kRt ����FORC�EUP�b܂FLUS
pH(N��� ��^6bD_CM�@E��7N� (�v�P��REM� Fa��@Pj���
K�	N����EFF/���@I�N�QOV��O{VA�	TROV� DT)��DTMX:e �P:/��P`q�vXpCLN A_�p��@ ��	_|�F�_T: �|�&P%A�QDI���`1��0�Y0RQ"m�_+qH���M���sCL�d#�RIV{��ϓN"EAR/�IOF�PCP��BR���CM�@N 1b �3GCLF��!DaY�(��a�#5T��DG���� �%%�FsSS� )�? P(q(1�1�`_1"8J11�EC13D;=5D6�GRA����@�����PW�OyN2EBUG�S��2�C`gϐ_E �A �?����/TERM�5B�5��O�ORIw�0C�5��SM_-`���0}D�6 �TA�9�E�5"��UP>��F� -Qϒ�A�P�3�@B$S�EGGJ� EL�UU�SEPNFI���pBx��1@��4>DC$sUF�P��$����Q�@C���G�0T������SNSTj�P�ATۡg��APTH	Jq�A�E*�Z%qB\`@F�{E��F�q�pARxP<Y�aSHFT͢qA|�AX_SHOR$��>��6 @$GqPE���OVR���aZP�I@P@$U?r *aAGYLO���j�I�"���Aؠ��ؠERV ��Qi�[Y)��G�@R���i�e��i�R�!P�uASYM���uqA#WJ�G)��E��Q7i�RD�U[d�@i�U��C�%UP���P���WkOR�@M��k0�SMT��G��GR��3�aPA�@��p|5�'�H � j��A�TOCjA7pP<]Pp$OPd�O�P�C�%�p�O!���RE.pR�C�AOX�?��Be5pR�E�ruIx'QG�e$PW�R) IMdu�RR_p$s��5��B Iz2�H8�=�_ADDR~H�H_LENG�BP�q�q:�x�R��So�mJ.�SS��SK������� ��-�SEh*���rSN�MN1K	�j�5�@r�֣OL��\�WpW�Q�>pACRO�p���@�H ����Q� ��OSUPW3�b_>�I��!q�a1�������� |��������-���X:���iIOX2S=��D�e��]���L� $��p�!_OFyF[r_�PRM_炽�rTTP_�H��M (�pOBJر"�pG�$H�LE��C��ٰN � �9�*�AB_�T���
�S�`�S��LV漣KRW"duHIT�COU?BGi�LO�q����d� �Fpk�GpSS� ����HWh�wA��O.���`INCPUX2VISIO��!��¢�.�á<�á-� �IwOLN)�P 87�yR'�[p$SL�b�d PUT_��	$dp�Pz �� �F_AS2Q/��$LD���D�aQT U�0]P�A������P�HYG灱Z�̱5�U9O� 3R `F����H�Yq�Yx�ɱvpP �Sdp���x��ٶ���UJ��S����NEΊWJOG�G �DI�S��r�KĠ��3T� |��AV��`_�C�TR!S^�FLAG�f2r�LG�dU ��n�:��3LG_SIZ��ň��=���FD��I����Z  �ǳ��0�Ʋ�@s��-� ��-�=�-���-��0-�ISCH_��Dq���N?���V��EE !2�C��n�U����r�`L�Ӕ�DAU�ՃEA��Ġt����G�Hr��OGBOO>)�WL ?`�� �ITV���0\�REC�SCRf 0�a��D^�����MARG ��`!P�)�T�/ty�?I�S�H�WW�I����T�JGM��MNC�H��I�FNKEY���K��PRG��UqF��P��FWD��HL�STP��V`��@�����RSS�H�` �Q�C�T1�ZbT�R ���U����� |R��t�i���G��8PCPO��6�F�1�M���FOCU��RGE]XP�TUI��I���c��n��n�� ��ePf���!p6�eP7�9N���CANAI�jB޾�VAIL��CL�t!;eDCS_HI�4�.��O�|!�S Sn�1^I�BUFF1XY�5�PT�$�� ��v��fīPN6q1Y�Y��P �����pO+S1�2�3����� 0Z � � ��aiE�*��ID%X�dP�RhrO�+��A&ST��R��Y�z�<! Y$EK&CK+���Z&m&�5�0[ L��o�0 ��]PL�6pwq�t^�����w��7�_ \ �`��瀰�7��#�0�C��] ��CL�DP��;eTRQL�I�jd.�094FLAGz�0r1R3�DM��R7��LDR5<4R5ORG.���e2(`���V��8.��T<�4�d^ A�q�<4��-4R5S�`�T00m��0DFRCLMC!D�?�?3I�@��MIC��d_ Yd���RQm�q��DSTB	�  ؏Fg�HAX;b |�H�LEXCESZrRnFMup�a`��B�;d�rB`��`a��F_A�J��$[�O�H:0K�db \��ӂnS�$MB��LIБ~}SREQUIR�R�>q�\Á�XDEBUT��oAL� MP�c�b�a��P؃ӂ!BoAND���`�`d�҆�c�fcDC1��IN�� ���`@�(h?Nz�@qܮ�o�NV�SPS�T8� e�rLO�C�RI�p�EXfA�p��AoAOD�AQP�f X��ON��[rMF�����f )�"I��%�e��T��!�FX�@IGG� g �q��"E�0�h�#���$R�a%;#�7y��Gx��VvCPi�D'ATAw�pE:�y���RFЭ�NVh t_ $MD�qIёA)�v+�tń�tH�`��P�u�|��sANSAW}��t�?�uD��)�b�	@Ði �@CU��V�T0�ewRR2�j Dɐ��Qނ�Bd$CALII�@F�G�s�2⠧RIN��v�<��NTE���kE���,�X�b����_Nl���ڂ��kDׄRm�DIViFDH�@ـn�$V��'c!;$��$Z������~�[��o�H �$BELT|b��!ACCEL+q��ҡ��IRC��t����T/!��$SPS�@#2LPqЀƔ83������� ��P�ATH��������3̒Vp�A_�Q�.�4��B�Cᐈ�_MGh�$DDQ���G�$FWh��p��m�؝���b�DE��PP�ABNԗROTS�PEED����00J��Я8��@��P$OUSE_��P��Fs�SY��c�A >q�YNu@Ag��OF�F�q�MOUN�N�Gg�K�OL�H�INC*��a��q��Bj�<L@�BENCS��q`�Bđ���D��IN#"�I̒��4�\BݠVE�O�w�Ͳ23_UP�E�߳LOWL ���00����D���B wP��� �1RCʀƶ�MOSIV�JRMO����@GPERCH  �OV��^� �i�<!�ZD<!�c�� d@�P��V1�#P͑��L���EW��ĸ�UP������TR�Kr�"AYLOA 'a�� Q-�̒<�1Ӣ`0 ��RTI$Qx�0 MO���МB R�0J��D��s�H����b��DUM2(�S_BCKLSH_C̒ ��>�=�q�#�U��ԑ����2�t�]ACLAL�vŲ�1n�P�CH�K00'%SD�RTY@4�k��y�1�q_6#N2�_UM$Pj�Cw��_�SCL��ƠLM?T_J1_LO��@���q��E�����p�๕�幘SPC��07������PCo���!H� �PU�m�C/@�"sXT_�c�CN_��1N��e���SFu���V�&#����9�̒��2=�C�u�SH6#�� c����1�Ѩ�o�0�͑�
��_�PAt�h�_	Ps�W�_10��4�R�P01D�VG�J� L�@�J�OGW���TO7RQU��ON*�M����sRHљ��_W��-�_=��C��I���I�I�II�F��`�JLA.�1[�VEC��0�D�BO1Up�@i�B\JRKU���	@DBL_S�Md�BM%`_DLC�BGRV��C��I��H_� ��*COS+\�(LN�7+X>$C�9)I�@9)u*c,)�Z2 �HƺMY@!�( "T�H&-�)THET0�NK23I��"=��A CB6CB=�C �A�B(261C�616�SBC�T25GTS QơC��aS$" ��4c#�7r#$DU D�EX�1s�t��B�6��r�AQ|r�f$NE�D�pIB U�\B5��$!��!A�%E(G%(!LPH$U�2׵�2SXpCc%pCr%�2�&P�C�J�&!�VAHV6HT3�YLVhJVuKV�KUV�KV�KV�KV�IHAHZF`RXM��wXuKUH�KH�KH�KH�KUH�IO2LOAHO�Y�WNOhJOuKO�KO��KO�KO�KO�&F��2#1ic%�d4GSP�BALANCE_l�!�cLEk0H_�%SP��T&�bc&�br&PFULC�hr�g�rr%Ċ1ky�UT�O_?�jT1T2Cy��2N&�v�ϰct�w�g�p�0Ӓ~���T���O���� INSsEGv�!�REV�v�!���DIF��1�l�w�1m�0OB0�q
����MIϰ1�~�LCHWAR��波AB&u�$MECH,1� :�@�U�AX:�P��Y�G$�8pn 
Z��|���7ROBR�CR���N�'�MSK�_�`f�p P 
Np_��R����΄ݡ�1��ҰТ΀ϳ���΀"�IN�q�M?TCOM_C@j�q  L��p��?$NORE³5�y��$�r 8� �GR�E�SD�0A�BF�$XYZ_�DA5A���DEBaU�qI��Q�s �`�$�COD�� ���k�F�f�$BUFINDXРw  ��MOR��/t $-�U��)��r�B��������G�ؒu � $SIMULT ��~��< ���OBJE�` ��ADJUS>�1�A'Y_Ik��D_�����C�_FIF�=�T� ��Ұ��{��p@� �����p�@��D��FRI��ӥT��RIO� ��E�{�͐�OPWO�ŀv}0��SYSBU�@ʐ$SOP�����#�U"��pPRUN,�I�PA�DH�D�\���_OU�=���qn�$}�IMA�G��ˀ�0P�qIM����IN�q���?RGOVRDȡ:����|�P~���Р�0L�_6p���i��RB����0��M���E�DѐF� ��N`Md*������˱SL�`�ŀw x $OwVSL�vSDI��DEXm�g�e�9w�$����V� ~�N���@w����Ûǖȳ�M��F͐�q<��� �x HˁE�F�AT+US���C�0à�ǒ��BTM����I
f���4����(�ŀy DˀEz�g���PE�r�����
���EXE��V��E�Y�8$Ժ ŀz @ˁ��3UP{�h�$�p��XN���9�H�� �PG"�{ h? $SUB��c��@_��01\�MPW�AI��P����LO��-�F�p�$R�CVFAIL_C�-�BWD"�F����DEFSPup | Lˀ`�D�� U�UNI��S�b��R`���_L�pAP��̐���ā}���� B�~���|��`ҲNN�`KET��y���P� $�~���0SIZE�ଠ{����S<�OR��FORMAT/p � F��ᖫrEMR��y�UqX�����PLI7�~ā  $�P_SWI�������_PL7�ALO_ �ސR�A���B�(0C��Df��$Eh����C_�=�U� � �c ���~�J3�0�����TIA4��5:��6��MOM������ �B�A�D��*��* PU70NRW��W �R����� A$PI�6���	�� )�4l�}69���Q���c�SPEED�PGq�7�D�>D� ���>tMt[��SAM�`痰8>��MOV���$���p�5��5�D�1�$2�������d{�Hip�IN?, {�F(b+=$�H*�(x_$�+�+GAMM�f|�1{�$GET���ĐH�D����
^pL�IBR�ѝI��$HI��_��Ȑ*B6�E��*8A$>G086LW=e6\<G9�686���R��ٰV��$PDCK�Q�H�_����;"��z�.%�7�4*�9� ��$IM_SRO�D�s"���H�"�LE�O�0\H���6@�� �ŀ�P~�qUR_SCR����AZ��S_SAV�E_D�E��NO��CgA�Ҷ��@�$�� ��I��	�I� %Z[ � ��RX" ��m�� �"�q�'"�8� Hӱt�W�UpS���
Q�M��O㵐.'}q ��Cg���@ʣ�����S�M�AÂ� � �$PY��$WH`'�NGp���H`���Fb��Fb��Fb��PLM���	� 0h�H�{�%X��O��z�Z�eT�M���� pS��C��O__0_B_�a:��_%�� |S��� �@	�v��v �@��ȯw�v��EM��% (�fr�B�ː��ft�P��PM��QU.� �U�Q��A�-�QTH=�HOLޛ�QHYS�ES��,�UE��B��O.#��  ��P0�|��gAQ���ʠu���O��ŀ�ɂv�-�A;ӎ�ROG��a2�D�E�Âv�_�ĀZ�INFO&��+�����bȜ�OI킍 =((@SLEQ/��#������o���DS`c0O�0�01�EZ0NUe�_�AUyT�Ab�COPY�P�Ѓ�{��@M��N������1�P�
� ��RiGI�����X_�P�l�$�����`�W��P��j@�G���EXT_CYCtb!���p����h�7_NA�!$�\��<�RO�`]�� � m��PORp�ㅣ���SRVt��)����DI �T_ l���Ѥ{�ۧ��ۧ Ъۧ5٩6٩7٩8�����S�B쐒���$�F6���PL8�A�A^�TAR��@ E `�Z�����<��d7� ,(@FLq`hѦ�@YNL���M�C���PWRЍ��=�e�DELAѰ��Y�pAD#qX� ��QSKIP�� iĕ�x�O�`NT!���P_x���� �@�b�p1�1�1� ��?� �?��>��>��&�>�3�>�9�Js2R;쐖 4��EX� TQ����ށ��Q���[�KFд�'��RDCIf� )�U`�X}�R�#%�M!*�0�)��$RGE7AR_0IO�TJB�FLG�igpER�a��TC݃������2�TH2N��� S1�b��Gq T�0' ����M���`qIb��v�REF��1�� l�h��E�NAB��lcTPE ?@���!(ᭀ��� �Q�#�~�+2 H�W�
��2�Қ���"�4�(F�X�j�3�қ{�������j�4�Ҝ���
��.�@�R�j�5�ҝu�����������
j�6�Ҟ��(L:L ���7���o�����j�8�Ҡ��"4�Fj�SMSK������a��E�A���MOTE�������@ "1��Q�IIO�5"%I��P���POWi@쐣 � �����X�gpi�쐤���Y"$DSB_S�IGN4A�Qi�̰C��ШP��RS232�%�Sb�iDEVI�CEUS#�R�RP�ARIT�!OP�BIT�Q��OWCONTR��Qⱬ��RCU� M�SU_XTASK�3NB���0�$TATU�P%�S@@쐦F�6��_�PC}�$FREEFROMS]p��ai�GETN@S�UKPDl�ARB73P%0����� !m$USA���az9ЎL�ERI�0f��pRIY�5~"_�@f�P�1��!�6WRK��D�9�F9ХFRIE3ND�Q4bUF��&��A@TOOLHFMY�5�$LENGT�H_VT��FIR��pqC�@�E� IU�FIN�R���R�GI�1�AITI�:�xGX��I�FG2�7G1a����3�B�GcPRR�DA��O_� o0e�I1RER�đ�3&���TC���AQJVG �G|�.2���F��1�!d�9Z�8+5K��+5��E�y�L0�4��X �0m�LN�T�3Hz��89��%�4�3%G��W�0�W�RdD�Z��Tܳ��K�a�3d��$cV 2!���1��I1H�0U2K2sk3K3J ci�aI�i�a�L��SLL��R$Vؠ�BV�E�Vk�]V*R��� � ,6Lc���9V2F{/P�:B��PS_�E���$rr�C�ѳ$A0��wPR���v�U�c1Sk�� {��6��G� 0���VX`�!�tX`��0P�Ё��
�5SK!� �"-qR��!0���z�MNJ AX�!h�A�@�LlA��A�THIC��1�������1TF�E���q>�IF_C	H�3A�I0�����G1�x������9��Ɇ_JF҇PR|(���RVAT�� �-p��7@�����DO�E��COU�(��AXIg��O�FFSE+�TRIG�SK��c���Ѽ�e��[�K�Hk���8�IG#MAo0�A-��ҙ��ORG_UNEV�����S�쐮�d �$�������GROU��ݓTqO2��!ݓDSP���JOG'��#	�_P'�2OR���>P67KEPl�IR�0�2PM�RQ�AP�Q���E�0q�e���SYS�G��"��PG��BRAK*Rd�r�3�-���0����ߒ<pAD�ݓ�J�BSOC� N��DUMMY14��p\@SV�PDE_�OP3SFSPD�_OVR��ٰC�O��"�OR-��Nı0.�Fr�.��OV��SFc�2�f��F���!4�S��RA�"L�CHDL�REC�OV��0�W�@M�յ�RO3��9_�0� @�ҹ@�VERE�$OF�S�@CV� 0BWD�G�ѴC��2j�
�T�R�!��E_F�DOj�MB_CM4��U�B �BL=r0�w�=q�tVfQ��x0spd��_�Gxǋ�AM��`k�J0������_M���2{�#�8$CA��{Й���8$HB�K|1c��IO��8.�:!aPPA"�N��3�^�F���:"�DVC_DB�C��d�w"����!��1���ç�y3����ATIO� �q0�UC�&CAB�BS�PⳐ�P�Ȗ��_0c�S�UBCPUq��S �Pa aá�}0�Sb��c���r"ơ$HW_AC���:c��IcA�A~-�l$UNIT��l��ATN�f�����CYCLųNEC�A��[�FLTR_2_FI���(��}&Ɩ�LP&�����_S[CT@SF_��F����G���FS|!�¹�CHAA/����2��RSD�x"ѡb��r�: _T��PROX��O�� EM�_�r��8u�q u��q��DI�0e�RAOILAC��}RMƐCLOԠdC��:anq���wq����PR��S�LQ�pfC�ѷ 	���FUNCŢ�rRINkP+a�0 ��!3RA� >R 
Я8�ԯWAR�#BLFQ��A�����DA�����LDm0�aB9�2�nqBTIvrb8ؑ���PRIAQ1�"AFS�P�!���𰠓�`%b���M�I1U�DF_j@��y1�°LME�FA�@H�RDY�4��Pn@R�S@Q�0"�MUL�SEj@f�b�q ��X��ȑ� lo .A$�1$c1� Ē���� x~�EG� ݓ��q!AR����09p>B�%��AXE���ROB��W�A4�_�-֣SY���!6��&MS�'WR���-1���STR��5�9�E�� 	5B��=QB90�@6������kOT�0o 	$�ARY8�w20����	%�FI��;�$�LINK�H��1��a_63�5�q�2XYZ"��;�q�3�@��1�2�8{0B�{D��� CFI��6G��
�{�_J��6��3a'OP_O4Y;5�Q#TBmA"�BC
�z��DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ ��@�5<:7�� +1�?0K�Mc�6�8Cb�vrb�4�ORQ��X�>8�#op�� ����wq�Uf�����T'OVE�Q��M;�@E#�UK#�UQ"�VW�Z Q�W���Tυ� ;� ���QH�!`�ҽ��U�Q��WkeK#kecXER��	GE	0��S�dAWaǢ:D���7!�!AX�rB! {q��1uy-!y �pz�@z�@z6Pz \Pz� z1v�y �y�+y�;y�Ky �[y�ky�{y��y��q�yDEBU��$����L�!º2WG`  AB!�,��S9V���� 
w��� m���w����1���1�� �A���A��6Q��\Q����!�m@��2CLAB3B�U�����So  V ER��>�� � $�@� mAؑ!p�PO���Z�q0w�^�_MR}Aȑ� d  9T�-�ERR��TYz�B�I�V83@�cΑTOQ�d:`�L� �d2�\�X�C�[! � p�`T8}0i��_V1�r�a('�4�2-�2<�����@P�����F�$QW��g��V_!�l�$�P����c��q�"�	V FZN_C;FG_!� 4��?� ��|�ų����@�ȲW8Z���\$� �n����Ѵ��9c�Q��(�FAp�He�,�XEDM� (�����!s�Q�g�yP{RV HELLĥ߷ 56�B_wBAS!�RSR��ԣo �#S��[��U1r�%��2ݺ3ݺU4ݺ5ݺ6ݺ7ݺ98ݷ��ROOI�̝0�0NLK!�CAB�� ��ACK��IN��T:�1�@�@ �z�m�_PU!�CO,� ��OU��P� Ҧ�) ��޶��TPF?WD_KARӑ�@&��RE~��P��(�QUE�����P
���CSTOPI_AL�����0&�������0SEMl�b�|��M��d�TY|�SOK�}�DI�����(����_TM\�MA'NRQ�ֿ0E+�|��$KEYSWI�TCH&	���H=E
�BEAT��c�E� LEҒ���U���FO�����O_�HOM�O�REF�PPRz��!&0ʉ�C+�OA�EC�O��B�rIOC�M�D8׵��'8��8�` � D�1����U��&�MH�»P��CFORC��� �]���OM�  �� @V��|�U�,3P� 1-�`� 3�-�4�p �SNP�X_ASǢ� 0�ȰADD����$�SIZ��$VA�Rݷ TIP]�\�2�A򻡐��Ȑ]�_� �"S꣩!C<ΐ��FRIF⢞�aS�"�c���NF�ҸV ��` � x�`S�I�TES�R6SSKGL(T�2P&���AU�� ) STMTdQZPm 6BW�P�*SHOWb���SV�\$�� ���A00P�a� 6�@�J�T�U5�	6�	7�	8�	9�	A�	� �!�'��C@�F�0u �	f0u�	�0u�	�@�u[Pu%121�?1L1Y1f1�s2�	2�	2�	2��	2�	2�	2�	2�22%222�?2L2Y2f2�s3P)3�	3�	3��	3�	3�	3�	3�33%323�?3L3Y3f3�s4P)4�	4�	4��	4�	4�	4�	4�44%424�?4L4Y4f4�s5P)5�	5�	5��	5�	5�	5�	5�55%525�?5L5Y5f5�s6P)6�	6�	6��	6�	6�	6�	6�66%626�?6L6Y6f6�s7P)7�	7�	7��	7�	7�	7�	7�77%727�?7,i7Y7Fi7�sA]�VP�UP}D��  ��x|�԰��YSLOǢ� � z��и� ��o�E��`>�^t��А�ALUץ����CU����wFOqID_L��ӿuHI�zI�$FILE_���t�ĳ$`�JvSA���� h���E_BL�CK�#�C,�D_CPU<�{�<�o�����tJr��R ���
PW O� -��LA��S��������RUNF�Ɂ�� Ɂ����F�ꁡ�ꁬ�_�TBCu�C� �X -$�LENi��v�����I��G�LOW_7AXI�F1��t2X�M����D�
 ���I�� ��}�TOR����Dh��� L=��⇒�s���#�_MA`�ޕ��ޑGTCV����T�� �&��ݡ����J������J����Mo���JH�Ǜ ��������2��� v�����F�JK��VKi�Ρv�Ρ�3��J0�ңJJvڣJJ�AALңP�ڣ��4�5z�&�N1-�9���␅�%L~�_Vj�9��ޠ�� ` �GR�OU�pD��B�N�FLIC��RE�QUIREa�EB�UA��p����2��������c��{ \��APPR��iC���
�EN��CLOe��S_M� v�,ɣ�
���7� ��MC�&����g�_MG�q�C�� �{�9���|�BRKz�NOL��|ĉ R��_LI|��Ǫ�k�J����P
���ڣ������&���/���6��6��8������� ��8�%��W�2�e�PATH a�z�p�z�=�vӥ�ϰm�x�CN=�CA������p�IN�UCh��bq��CO�UM��!YZ������qE%����2������PAYL�OA��J2L3pR'_AN��<�L��F��B�6�R�{�R_F2�LSHR��|�LO�G��р��ӎ���ACRL_u�������.�r��H�p�$H{�^��FLEX
��}J�� :� /����6�2�����;�M�_�F16����n�@��������ȟ��Eҟ �����,�>�P�b� ��d�{�������������5�T��X ��v���EťmF ѯ�������&��/�A�S�e�'	�x�� � ������j��4pAT����n�EL�  �%øJ���vʰJE��CTR�і��TN��F&��H�AND_VB[�
�pK�� $Fa2{�6� �rSWi���("U��� $$Mt�h�R��08�� @<b 35��^6A�p3�k��q{9t�A�̈p��A��A�ˆ0��U���UD��D��P��G���IST��$A��$AN��DYˀ�{�g4�5 D���v�6�v��5缧�^�@��P����@�#�,�5�>�D�J�� &0�_�ER!V<9�SQASYM��] 	�����x��ݑ���_SHl�������sT@�(����(�:�JA����S�cir��_V�I�#Oh9�``V_�UNI��td�~�J ���b�E�b��d��d �f��n���������u�N���5D��H̟�����"CqENL� a�DI��>�Obt8<rDpx�� ��2IxQA����q��-���s �� s����� ���OMME���rr�QTVpPT@�P ���qe�i�����P�x ��yT�Pj�� $DUMMY}9�$PS_��RFq�  ��:�� s���!~q� �X����K�STs��ʰSBR��M21�_Vt�8$SV_�ERt�O��z���C+LRx�A  O�r?p�? Oր � D $GLOB���#LO��Յ$�o���P�!SYSA�DR�!?p�pTCH>M0 � ,��ސ�W_NA���/�e���D�SR��l (:]8: m�K6�^2m�i7m�w9 m��9���ǳ��ǳ��� ŕߝ�9ŕ���i� L���m��_�_�_�T>D�XSCRE�ƀ5�� ��STF���#}�pТ6�<q] u_v AŁ� T����TYP�r�K��Pu�!u���O�@�IS�!��tC�UE{t� ����H�yS���!RSM_��XuUNEXCEPWv��CpS_��{ᦵ��ӕ���÷���CO�U ��� 1�O�UET�փr����PROGM� FL�n!$CU��POX*q��c�I_�pH;�� � 8��N�_�HE
p��Q��pRY ?���,�J�t*��;�OUS�� � @d���_$BUTT��R@�>��COLUM�íu��SERVc#=�P�ANEv Ł� �; �PGEU�!��F��9�)$HELyP��WRETER��)״���Q��� ���@� P�P �SIN��s�PNߠ�w v�1����� ����LN�ړ ����_��k�s$H��M TEX�#�����FLAn +RELV��D4p���j����M��?,��ӛ$����P=�U�SRVIEWŁ�S <d��pU�p0�NFIn i�FOC�U��i�PRILP�m+�q��TRIP>)�m�UNjp{t�� QP��XuWA�RNWud�SRTO�LS�ݕ�����O�|SORN��RAU�ư��T��%��VI�|�zu� $��PATHg��CwACHLOG6�O�LIMybM���'���"�HOST6��!�r1�R�OB�OT5���IMl� D�C� g!��E�L����i�VCPU_A�VAILB�O�EX
7�!BQNL�(���A0�� Q��Q ��.ƀ�  QpC���@$TOOL6��$�_JMP� ��I�u$SS��!$<qVSHIF��|s�P�p�6��s���R���OSU�RW�pRADIz��2�_�q�h�g!� �q)�LUza�$OUTPUT_3BM��IML�oRp6(`)�@TIL<'SCO�@Ce�; ��9��F��T��a ��o�>�3�����w�2u�b�V�zu✫�%�DJU��|#_�WAIT������%ONE���YBOư ��� $@p%�C�S�Bn)TPE��NE�C��x"�$t$���*B_T��R��%�qRH� ���sB�%�tM�+ ��t�.�F�R!݀���OPm�MAS�_�DOG�OaT	�D�����C3S�	�O2DE�LAY���e2JO ��n8E��Ss4'#J�aP`6%�����Y_��O2$��2���5��`?� r'�Z�ABCS��  �$�2��J�
b���$$CLAS�����AB�b�'@@VIRT��O.@gABS�$�1 <E�� < *AtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v�p����M@[�AXLրtK�*B�dC  ����IN��ā��PRE������LA�RMRECOV c<I䂥�NG��� \K	 A �  J�\�M@PPL�IC�?<E��E�Hand�lingTool� �� 
V7.�50P/28[� � �����
��_SW�� UPn*A� ��F0ڑ䢒��A@��� 20��*A����:���X�FB 7DA5��� '@���@��None엃���� ���T�*A4y�Wxl�_��V��t��g�UTOB��ค����HGAPCON8@��LA��U��oD 1<EfA���������� /Q 1שI Ԁ��Ԑ�:�i�n�����#B)B g���\�HE��Z�r�HTTHKY��$BI�[�m��� ��	�c�-�?�Q�o�u� �ϙϫϽ�������� _�)�;�M�k�q߃ߕ� �߹��������[�%� 7�I�g�m����� ��������W�!�3�E� c�i�{����������� ����S/A_e w������� O+=[as� ������K// '/9/W/]/o/�/�/�/ �/�/�/�/G??#?5? S?Y?k?}?�?�?�?�? �?�?COOO1OOOUO gOyO�O�O�O�O�O�O ?_	__-_K_Q_��(��TO4�s���DO_CLEAN��e��S�NM  9� �9oKo]ooo�o�DSPDRYR�_&%�HI��m@&o�o �o#5GYk} ����"���p�Ն# �ǣ�qXՄ���ߢ��g�PLUGGpҠ�Wߣ��PRC�`B`9��o�=��OB��oe�SEGF��K������o%o�����#�5�m���LAP�oݎ���������� џ�����+�=�O�|a���TOTAL�|.���USENUʀ�׫ �X���R(�R�G_STRING� 1��
�kM��Sc�
���_ITEM1 �  nc��.�@�R�d� v���������п������*�<�N�`�r��I/O SIG�NAL��Tr�yout Mod�e�Inp��S�imulated��Out���OVERR�` =� 100�In� cycl����Prog Abo�r�����Sta�tus�	Hea�rtbeat��MH FaulB�K�AlerUم�s� �ߗߩ߻��������� �S���Q� �f�x�������� ������,�>�P�b��t�������,�WOR ������V��
. @Rdv���� ���*<N`PO��6ц�� o�����// '/9/K/]/o/�/�/�/��/�/�/�/�/�DEV�*0�?Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O>�OPALTB��A ���O�O__,_>_P_ b_t_�_�_�_�_�_�_��_oo(o:o�OGRI�p��ra�OLo�o�o �o�o�o�o*< N`r������`o��RB���o� >�P�b�t��������� Ώ�����(�:�L��^�p����PREG �N��.�������� *�<�N�`�r������� ��̯ޯ���&��Ϳ�$ARG_��D ?	���i���  �	$��	[�}�]}���Ǟ�\�S�BN_CONFIOG i��������CII_SA_VE  ��۱�Ҳ\�TCELLSETUP i��%HOME_I�O�͈�%MOVq_�2�8�REP����V�UTOBAC�K
�ƽ�FRA:\�� ��Ϩ���'` ��������  ����$�6�c�Z�lߙ��Ĉ���������� ���!凞��M�_�q� ����2�������� �%�7���[�m���� ����@�������!3E$���Jo��������INI��@��ε��MESSAG����|q��ODE_D$����O,0.��P�AUS�!�i� ((Ol��� ����� /�/ /$/Z/H/~/l/�/�'�akTSK  �q�����UPDT�%�d0;WS�M_CF°i��еU�'1GRP Y2h�93 |�B���A�/S�XSCRDv+11
1; ����/�?�?�? OO $O��߳?lO~O�O�O �O�O1O�OUO_ _2_�D_V_h_�O	_X���G�ROUN0O�SU�P_NAL�h�	��ĠV_ED� 1�1;
 �%-BCKEDT-�_0`�!oEo$���a(��o�����ߨ���e2no_˔o�o�b���ee�o"�o�oED3�o�o ~p[�5GED4� n#�� ~�j���ED5Z��Ǐ6� ~p���}���ED6�� ��k�ڏ ~G���!�3�ED7��Z��~� ~p�V�şןED8F�&o��Ů}����i�{�ED9ꯢ�W��Ư
}3�����CRo�����3�տ@�����P�PNO_D�EL�_�RGE_U�NUSE�_�TLA�L_OUT �q�c�QWD_AB�OR� �΢Q��IT_R_RTN����ONONSe����CAM_PAR�AM 1�U3
� 8
SONY� XC-56 2�34567890��H � @����?���( SАV�|[r؀~�X�HR5k�|U�Q��߿�R57����A�ff��KOW�A SC310M�|[r�̀�d @6�|V��_�X� ����V��� ���$�6���Z�l��CE_R�IA_I857�F�1��R|]]��_LIO4W=V� ��P<~�F<��GP 1�,����_GYk*Cg*  ��C1� �9� @� G� �CVLC]� d� l� Es�R� ��[�Um� v� � �� _�� C�� �"��|W��7�HEӰO�NFI� ��<G_�PRI 1�+ P�m®/���������'CHKPA�US�  1E� ,�>/P/:/t/^/ �/�/�/�/�/�/�/?�(??L?6?\?�?"OƩ����H�1_MkOR�� �0�5 	 �9 O�?�$OOHO6K�2	��H�=9"�Q?55��CR�PK�D3P����>��a�-4�O__|Z
�OG_�7�P O�� ��6_��,xV�A�DB���='�)
�mc:cpmidcbg�_`��S:�(�	���Yp�_)o�S`�BBi�P�_mo8j�(�Koo�oV9i�(��og�o�o�m�of�oGq:�I�ZDEF �f8��)�R6pbuf.txtm�]nd�@����# 	`(н��A=L���zM-C�21�=��9����4�=�n׾�C�z  BHBCCo��C|��Cq�D��C�?��C�{iSZE@�D��F.���F��E⚵F,E�ٙ��E@F�N�IU���I?O�I<�#I6�I�I�SY���vqG����Em�(�.���(�(��<�q�G�)x2��Ң �� a��D�j���E�e��E�X�EQ�E�JP F�E�F� G�ǎ�^F E�� F�B� H,- Ge��H3Y����  >�33 ����xV  n42xQ@��5Y��8B� A�AST<#�
�� �_'�%��wR_SMOFS���~�2�yT1�0DE ��O c
�(�;�"�  <�6�z��R���?�j�C4R��SZm� W���{�m�C��B-G�CR�`@$�q��T{��FPROG %i����c�I��� �����f�KEY_TB�L  �vM�u� ��	
�� �!"#$%&'(�)*+,-./0�1c�:;<=>?�@ABC�pGHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������p���͓���������������������������������耇�������������������s��!j�LCK��x.�j���STAT����_AUTO_D�O���W/�IND�T_ENB߿2R���9�+�T2w�XS�TOP\߿2TRL^l�LETE�����_SCREEN �ikcs�c��U��MMEN�U 1 i  <g\��L�SU+� U��p3g������ ������2�	��A�z� Q�c������������� ��.d;M� q������ N%7]�m ���/��/J/ !/3/�/W/i/�/�/�/ �/�/�/�/4???j? A?S?y?�?�?�?�?�? �?O�?O-OfO=OOO �OsO�O�O�O�O�O_��O_P_Sy�_MA�NUAL��n�DB;COU�RIG��ٟDBNUM�p���<���
�QPXWO_RK 1!R�ү��_oO.o@oRk�Q_�AWAY�S��G�CP ��=��df_CAL�P�db�RY��������X_�p 1">�� , 
�^����o xvf`MT�I�^�rl@�:sONT�IM�������Zv�i
õ�cMOT�NEND���dRECORD 1(R�qa��ua�O��q ��sb�.�@�R��x Z�������ɏۏ� ����#���G���k�}� ����<�ş4��X�� �1�C���g�֟���� ����ӯ�T�	�x�-� ��Q�c�u�������� ��>����)Ϙ�M� ��F�࿕ϧϹ���:� ������%�s`Pn&�]� o��ϓ�~ߌ���8�J� ����5� ��k��� �ߡ��J�����X�� |��C�U�������� ���0�����	��db�TOLERENC�qdBȺb`L����PCS_CFG �)�k)wdM�C:\O L%04�d.CSV
�Pcl�)sA �CH� z�P)~���h�MRC_OUT �*�[�`+P S�GN +�e�r���#�10-MA�Y-20 10:�18*V17-FE�Bj9:09�k? PQ�8���)~�`pa�m��PJPѬ�VERSION� SV2�.0.r3wEFLOGIC 1,�[/ 	DX�P7)��PF."PROG_�ENB�o�rj UL�Sew �T�"_WRSTJNEp�V�r�`dEMO_OPT?_SL ?	�es�
 	R575)s7)�/??*?<?|'�$TO  �-د�?&V_@pEX�Wd�u�3PAT�H ASA\p�?�?O/{ICT�a-Fo`-�gds�egM%&ASTBF_TTS�x@�Y^C��SqqF�P�MAU� t/XrMS%WR.�i6.|
S/�Z!D_N�O0_�_T_C_x_g_�_�tSBL_FAUL"y0�[3wTDIAU �16M6p�A�1234567G890gFP? BoTofoxo�o�o�o�o �o�o�o,>Phb�S�pP�_ ���_s�� 0`�� ���)�;�M�_�q� ��������ˏݏ��|�)UMP�!� �^�TR�B�#+�=��PMEfEI�Y_T�EMP9 È�3p@�3A v�UNI�.�(YN_BRK �2Y)EMGDI_STA�%WЕ�NC2_SCR 3��1o"�4�F� X�fv���������#��ޑ14�����)�;�����ݤ5�����x�f	u�ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/߭P�b�t� � ��xߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N���r����� ����������& 8J\n���� ����"`�F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ 4?,?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�O �O�O?�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�O�O�o�o �o
.@Rdv �������� �*�<�N�`�r����o ����̏ޏ����&� 8�J�\�n����������ȟڟ����H�ETMODE 16���� ���ƨ
R�d�v�נRR�OR_PROG �%A�%�:߽� � ��TABLE  A������#��L�RRSEV_N�UM  ��Q���K�S���_A�UTO_ENB � ��I�Ϥ_NONh� 7A�{�R�_  *������%������^�+��Ŀ8ֿ迄�HISO�͡�I�}�_ALM 1]8A� �;�����+�e�wωϛ�ȭϿ��_H���  �A���|��4�T�CP_VER �!A�!����$EX�TLOG_REQ���{�V�SIZ�_�Q�TOL  �͡Dz��A Q�_BWD����r����n�_DI�� 9��}�z�͡m���STEP����4���OP_DO����ѠFACTOR_Y_TUN�dG��EATURE �:����l��Handling�Tool ��  �- CEng�lish Dictionary���ORDEAA� Vis�� Ma�ster���96� H��nalog� I/O���H5�51��uto S�oftware �Update  ���J��matic Backup��Part&�g�round Ed�it��  8\a�pCamer�a��F��t\j6�R�ell���LO�ADR�omm��syhq��TI" ���co��
! o����pane�� �
!��tyl�e select.��H59��nD���onitor��4�8����tr��Re�liab���ad�inDiagnos"����2�2 �ual Chec�k Safety� UIF lg\�a��hanced� Rob Ser}v q ct\���lUser Fr�U��DIF��Ext. DIO ��fiA d��e�ndr Err L,@��IF�r�� � �П�90��FCTN MenuZ �v'��74� TPw In��fac�  SU (�G=�p��k Ex�cn g�3��Hi�gh-Sper S�ki+�  sO�H�9 � mmunic�!�onsg�teu�r� ����V�����conn��2���EN��Incr�stru���5�.fdKAR�EL Cmd. ML?uaA� O��Run-Ti� E�nv����K� ��+�%�s#�S/W��7�4��Licens�eT�  (Au�* ogBook(�Sy��m)��"�
MACRO�s,V/Offsme��ap��MH� ܷ���pfa5�Me�chStop Pgrot��� d�zb i�Shif��^��j545�!xr x��#��,��b �ode Swit�ch��m\e�!o�4.�& pro��4��g��Multi-T7G���net.Po=s Regi��z��P��t Fun����3 Rz1��NCumx �����9m�|�1�  Adjuj���1 J7�7�* x����6tatuq1�EIKRDM�tot��scove�� ��@By- �}uest1�$Go�� � U5\SNPX b"���YA�"Libr���Ŀ#�� �$~@h�pd�]0�Jts in VCCM�����0��  �u!��2 RL�0�/I�08��TMILIB�M �J92�@P�Ac�c>�F�97�TP�TX�+�BRSQe9lZ0�M8 Rm���q%��692��Un�exceptr m�otnT  CV1V�P���KC������+-��~K  II�)�VSP CSXC�&.c�� e�"��{ t�@WewΌAD Q�8bvr� nmen�@�i%P� a0y�0�pf�GridAplay !� nh�@*�3R��1M-10iA(_B201 �`2V"�  F���scii��load��83� M��l����Gu{ar�d J85�0��mP'�L`���st�uaPat�&]$Cyqc���|0ori_ �x%Data'Pqu���ch�1��g`ڂ j� RLJam��5���IMI D�e-B(\A�cP" �#^0C  et�kc^0asswo\%q�)650�Ap�U�Xnt��Pve�n�CTqH�5�0�YELLOW �BO?Y��� Arc�0vis��Ch��WeldQciail4Izt�Op� X��gs�` 2@�a��poG yRjT11 NE�#HT� 3xyWb��! �pB�`gd`���p\� =P���JPN ARC�P*PR�A�� wOL�pSup̂fil�p��J�� ��7cro�670�1CX~E�d��SS�pe��tex�$ �P� S�o7 t� ssagN5 <Q�BP:� �9 "0�QrtQC��9P�l0dpn�笔��rpf�q�e�ppm�ascbin4�psyn�' pt�x]08�HELN�CL VIS P�KGS �Z@MBq &��B J8@�IPE GET_�VAR FI?S �(Uni� LU�OOL: ADD�@_29.FD�TCm���E�@DVp���`�A�ТNO WTW�TEST �� �x�!��c�FOR �ЯECT �a!� ALSE ALA`��CPMO-130���� b D: HANG FROMg���2��R709 �DRAM AVA�ILCHECKS� 549��m�VP�CS SU֐LI/MCHK��P�0x��FF POS� F��� q8-1�2 CHARS�E}R6�OGRA ���Z@AVEH�AME���.SV��Вאn�$��9�m "y�T�RCv� SHAD~P�UPDAT k�}0��STATI�~�� MUCH ����TIMQ MO?TN-003���@OBOGUIDE DAUGH��p�b��@$tou� �@C� �0��PAT�H�_�MOVET��� R64��VM�XPACK MA�Y ASSERT�jS��CYCL`�T�A��BE CORg 71�1-�AN���RC OPTIO�NS  �`��AP�SH-1�`fix��2�SO��B��XO�����_T��	�i��0�j��du�byz p� wa��y�٠HI�������U�pb XS�PD TB/�F� /\hchΤB0����END�CE�06\�Q�p{ smay� n@�pk��L >��traff#�	�� ��~1from� sysvar scr�0R� ��d�'DJU���H�!A���/��SET E#RR�D�P7�����NDANT SC�REEN UNR?EA VM �PD�MD��PA���R�?IO JNN�0��FI��B��GRO;UNנD Y�Т�٠�h�SVIP �53 QS��DIGIT VERS���ká�NEW�� P�06�@C�1IMA�G�ͱ���8� D�I`���pSSUE��5��EPLAN {JON� DEL����157QאD��CALLI���Q��m�ޥ�IPND}�IM�G N9 PZ�1�9��MNT/��EsS ���`LocR �Hol߀=��2�PnN� PG:��=�M���can����С:� 3D mE2vi?ew d X���ea1 �0b�pof� Ǡ"HCɰ�A�NNOT ACC�ESS M cp�ie$Et.Qs a�� loMdFlex�)a:��w$qmo G�sA9�-'p~0���h0pa��eJ A�UTO-�0��!i�pu@Т<ᡠIAB�LE+� 7�a FP�LN: L�pl� m� MD<�VI��и�WIT HO�C�Jo~1Qui���"��N��USB��@�Pt & re�mov���D�vAx?is FT_7�P�GɰCP:�OS�-144 � h �s 268QՐOS�T�p  CRASoH DU��$P���WORD.$�L�OGIN�P��P:�	�0�046 is�sueE�H�: �Slow st
�c�`6����໰�IF�IMPR��S?POT:Wh4����N1STY��0VM�GR�b�N�CATZ��4oRRE�� N� 58�1��:%�'RTU!Pe -M a�SE:�@pp���A�GpL��m@acll��*0a�OCB� WA���"3 C�NT0 T9DWr}oO0alarm�ˀm0d t�M�"0��2|� o�Z@OM�E<�� ��E%  #�1-�SRE��M�s�t}0g    } 5KANJI5?no MNS@��INISITAL�IZ'� E�f�w�e��6@� dr�@ �fp "��SCI�I L�afail�s w��SYS�TE[�i��  �� Mq�1QGro8�m n�@vA�����&��n�0q��RW{RI OF Lk�>�� \ref"�
��up� de-re�la�Qd 03.��0SSchőbe�twe4�IND �ex ɰTPa�D�O� l� �ɰG�igE�soper�abil`p l,�HcB��@]�le<�Q0cflxz������OS {����v�4pfigi GLA��$�c2�7H� l�ap�0ASB� I�f��g�2 l\c��0�/�E�� EOXCE 㰁�P��H�i�� o0��Gd`�]Ц�fq�l lx9t��EFal��#�0�i�O�Y�n�CLO�S��SRNq1NT
^�F�U��FqKP�A?NIO V7/ॠ�1�{����DB ��0��ᴥ�ED��DSET|�'� �bF��NLINEb�BU�G�T���C"RLI�B��A��ABC �JARKY@��� orkey�`IL����PR��N��ITGAR� D$�R �Er *�T��a�U�0x��h�[�ZE V�� TASK p.vr�P2" .�Xf�J�srn�S谥dIcBP	c���B/��wBUS��UNN�A j0-�{��cR'�v��LOE�DIVS�CULs$cb����BW!��R~�W`P�L����IT(঱tʠ��OF��UNEXHڠ+���p�FtE���SVEMG3`NM_L 505� D*�CC_SAFE�P�*� �ꐺ� PETp��'P�`�F  !�F��IR����c i �S>� K��K�H GUNCHG���S�MECH��M$��T*�%p6u��t�PORY LEA�K�J���SPExgD��2V 74\�GRI��Q�g��C7TLN��TRe @��_�p ���EN'�IN������$���r��sT3)�i�STO�IA�s�L��͐X	����q��Y� ��T!O2�J m��0F<�K�L���DU�S��O��I3 9�J F��&���SSVGN-q1#I���RSRwQDAU�Cޱ� �T6�g���� 3�]���BRK�CTR/"� �q\j�5��_�Q�S�qIN=VJ0D ZO�Pݲ ���s��г�Ui ɰ̒��a�DUAL� �J50e�x�RVO_117 AW�TH!pHr%�N�247%��52��|�&aol @���R���at�Sd�cqU���P,�LER���iԗQ0�ؖ  ST����Md�Rǰt� /\fosB�A�0Np��c����{�U��ROOP 2�b�pB��ITP4M��b� !AUt c0< � p�lete�N@�� z1^qR635 �(AccuCal�2kA���I) "P�ǰ�1a\�Ps�� ǐ� bЧ0P򶲊����ig\cbacul "A3p_ �1���ն���etacea��AT���PC�`������_p�.p�c!Ɗ��:�cir1cB���5�tl��B���:�fm+�Ί�V��b�ɦ�r�upfr�m.����ⴊ�xepd��Ί�~�pedA��D �}b�ptliabB�� �_�rt��	Ċ�_\׊ۊ�6�fm�݊�oޢ�e��̈�Ϙ���c�Ӳ�5�j>�����tcȐ��	�Qr����mm 1��FT�sl^0��T�m�L��#�rm3��ub �Y�q�std}��pl;�&�ckv�=�r��vf�䊰��9�vi����ul�`�0fp��q �.f��� �daq; i Dat�a Acquisi��n�
��T`���1�89��2�2 DMCM R�RS2Z�75��~9 3 R710�o59p5\?���T "��1 (D�T� nk@���������E Ƒȵ��Ӹ�egtdmm ��ER�����gE��1�q\mo?۳�=(G����[(

�2�` !� �@JMACR�O��Skip/Offse:�a��V��4o9� &qR66!2���s�H�
 E6Bq8����9Z��43 J77� 6�J783�o ���n�"v�R5I�KCBq2 PTL�C�Zg R�3 (�s, �������03�	зJԷ�\sfmnmc "MNMC����ҹ��%mnf�FMC�"Ѻ0ª etmc�r� �8����� ,��D���   87?4\prdq>,�jF0���axis�HProcess� Axes e�r;ol^PRA
�Dp~� 56 J81j�[59� 56o6� ئ��0w�690 98� [!IDV�1��2q(x2��2ont�0 �
����m2���?�C��etis "�ISD��9�� FpraxRAM�P� D��defB�,�G��isbasic�HB�@޲{6�� 7�08�6��(�Ac w:������D
�/,��AMOX�� ��DvE���?;T��>Pi� RAF!M';�]�!PAM�V �W�Ee�U�Q'
bU��75�.�ceNe�� nterfac�e^�1' 5&!54x�K��b(Devam ±�/�#���/<�Ta=ne`"DNEWE����btpdnui �AI�_s2�d_r�sono���bAsf�jN��bdv_ar�Fvf�xhpz�}w��h9kH9xstc��g�AponlGzv{�ff��r���z��3{q'Td>pch'ampr;e�p� ^5977��	܀�4}0��mɁ�/�����lf�~!�pcchmp]a�MP&B�� �mp�ev�����pc�s��YeS�� Ma�cro�OD��16 Q!)*�:$�2U"_,��<Y�(PC ��$_�;������o��J�ge�gemQ@GEMS�W�~ZG�gesndxy��OD�ndda���S��syT�Kɓ�s!u^Ҋ���n�m���L���  ���9:p�'ѳ޲��spotplusp���`-�(W�l�J�s��t[�׷p�key�ɰ�$���s�-Ѩ�m���\fewatu 0FEAWD��oolo�srAn'!2 p���a�A�s3��tT.� (N. A.)��!eP!�J# (j�,��0�oBIB�oD -�.�mn��k9�"K���u[-�_���p� "�PSEqW����wop "sEЅ�&� :�J������y�|��O 8��5��Rɺ���ɰ [��X�������%�@(
ҭ�q HL�0 k�
�z�a!�B�Q�"(g�Q�����]� '�.�����&���<�!��_�#��tpJ�H�~Z ��j�����y������ �2��e������Z���� V��!%���=�]�͂���^2�@iRV� o%n�QYq͋JF0� !8ހ�`�	(^�dQueue���X\1��ʖ`�+F1tpvt�sn��N&��ftp:J0v �RDV�	f�H�J1 Q���v��en��kvstk✐mp��btkc�lrq���get����r��`�kack�XZ�sctrŬ�%�stl��~Z�np:!�`�@��q/�ڡ6!l�/HYr�mc�N+v3��_� ����.v��/\jF��� ��`Q�΋ܒ�N50 (FRA��+��͢fraparm���Ҁ�} 6�J64�3p:V�ELSE�
#�VAR $S�GSYSCFG.�$�`_UNITS 2�DG~°@�4Jg�fr��4A�@FRL -��0ͅ�3ې���L �0NE�:�=�?@�8�v�9~Qx304��;�BPRSM~QA�5�TX.$VNUM�_OL��5��DJ5�07��l� Functʂ"qwAP��琎��3 H�ƞ�kP9jQ�Q5ձ� ��@jLJzBJ[�6N�kAP�����S��"TPP�R���QA�prn�aSV�ZS��AS8Dj�510U�-�`cr �`8 ��ʇ�DJR`jY�ȑH  ژQ �PJ6�a21���48AAVgM 5�Q�b0 lBު`TUP xb�J545 `b�`6�16���0VC�AM 9�CL�IO b1�59 ���`MSC8�
r�P R`\sS�TYL MNIN��`J628Q  ��`NREd�;@�`S�CH ��9pDCS�U Mete�`O�RSR Ԃ�a04� kREIOCu �a5�`542�b9vpP<�nP�a�`�R��`7�`�MA�SK Ho�.r7y �2�`OCO :��r3��p�b�p���r�0X��a�`13\m�n�a39 HRM�"�q�q��LC�HK�uOPLG \B��a03 �q.�pOHCR Ob�pCp�Posi�`fP6 {is[rJ554��N�pDSW�bM�D�p�qR�a37 }Rjr0� �1�s4 �R6�76��52�r5 �2�r�7 1� P6���R_egi�@T�u/FRDM�uSaq%��4�`930�uSN{BA�uSHLB̀�\sf"pM�NP�I�SPVC�J�520��TC�`"{MNрTMIL�{IFV�PAC W��pTPTXp6.�%�TELN N �Me�09m3�UECK�b�`UFyR�`��VCOR���VIPLpq89qSsXC�S�`VVF��J�TP �q��R6�26l�u S�`G�ސ�2IGUI\�C��PGSt�\ŀH863�S�q����ւq34sŁ68�4���a�@b>�3 �:B��1 T��96u .�+E�51 yf�q53�3�b1 ��f�b1 n�jr9 ��`VAT ߲�q7�5 s�F��`�sAW�SM��`TOP �u�ŀR52p���a8s0 
�ށXY q�澢0 ,b�`885�QXрOLp}�"p�E࠱tp�`LCM<D��ETSS����6 �V�CPE 9oZ1�VRCd3
��NLH�h��001m2Ep��3 f��p��4 /165C���6l���7PR��0�08 tB��9 -�200�`U0�pFL�1޲1 ��޲2L"����p��޲4��5� \hmp޲6 RBCF�`ళ�fsః8 �Ҋ��~�J�7� rbcfA�L�8`\PC����"�32m0�u�n�K�Rٰn�5 �5EW
n�9 �z��40 kB��3� ��6ݲ�`00iKB/��6�u��7�u���8 µ������sU�0�`�t �1 05w\rb��2 E� ��K���j���5˰���60��a�HУ`:�6�3�jAF�_���F�7 ڱ݀H�8�eHЋ��c�U0��7�p��1�u��8u��9 713������D7� �ҹ5t�97 ��8�U�1��2��1�1:���h��1np�"���8(�U1��\py�l��,࿱v ��B�8�54��1V���D�4��im��1�<��H�>br�3pr�4@pGPr�6 B���цp���1����1�`͵1{55ض157 �2��62�S����!1b��2����1Π"��2���B6`�1�<c�4 7B�5 �DR��8_�B/��1�87 uJ�8 0�6�90 rBn�1� (��202 0EW,ѱ2^��2��90�U2�p�2��2� b��4��2�a"�RB����9\�U2�`w�l���4 60Mp��7������b�s
5 ��3����pB"9 3 ����`6ڰR,:7 �2��V�2��5���2^��$a^9���qr����n�5����5᥁"��8a�Ɂ}�5B���5����`UA���� ��Y86 �6 S�0���5�p�2�#�529A �2^�b1P�5~�2`���&P5��8��5��u�!ѹ5��ٵ544��5��R�ąP nB^z�c (�4������U5J�V�5��1��1^��%�����5 b21��gA���58W82� rbr��5N�E�5890tr� 1�95 �" ������c8"a��|�PL ���!J"5|6��D^!�6��B�"8�`#��+�8%�6B�AyME�"1 iC��'622�Bu�6V��dڸ 4��84�`AN�RSP�e/S� C�5� �6� ��� �\� �6� �V� 3t~��� T20CA�R��8� Hf� 1DH��� AOE� ��� ,�|�� ��0\�� �!64K���ԓrA� �1 (M-=7�!/50T�[PM��P�Th:1�C�@#Pe� �3�0� 5`M75T"� �D8pC� �0Gc� u�4��>i1-710i�1� �Skd�7j�?6�:-HS,� �RN�@�U�B�f�X�=m75!sA*A6an���!/C,B�B2.6A �0;A �CIB�A�2�QF1�UBu2�21� /70�S� �4����Aj1�3�p���r#0 B2\	m*A@C��;bi"i1�K�u"A~AAU� imm7c7��ZA@I$�@�Df�A�D5*A�EF� 0TkdR1�35Q1@�"*�@�Q�1�QC)P �1*A�5*A�EA�5B,�4>\77
B7=Q�D��2�Q$B�E7�C�D/qAHEE�W7�_|`j�z@� 2�0�Ejc7P�`�E"l7�@7�A 
1�E�V~`�W2%Q�R�9ї@0L_�#�@���"A���b��H3s=rA/2�R5nR4��74rNUQ1ZU�A�s\;m9
1M92L2�!�F!^Y�ps� 2ci��-?�qhimQ�t   w043�C�p2�mQ�r�H_ �H20�Evr�QHs�XBSt62�q`s������ ��Pxq350_*A3I)�2�d�u�0�@� '4TX�06�pa3i1A3sQ�25�c��st�r�VR1%e�q0
��j1� �O2 �A�UEiy�.� ‐ �0Ch20$CXB79#A�ᓄM Q1]�~�� 9�Q��?PQ ��qA!Pvs� 5	15 aU���?PŅ���ဎ�Q9A6�zS*�7��qb5�1����Q��00P(��V7]u�ait E1���ïp?7� !?��z��rbUQRB1PM=�Qa9��H��QQ�25L�������Q��@L��8ܰ��y�00\ry�"R2�BL�tN  ��� �1D�� �2�qeR�5����_b�3�X]1m1lcBqP1�a�E�Q� 5F�䥒�!5���@M-16Q�� f���r��Q��e� ��� PN�LT�_�1��i1��9453���@�e�|�b1l >F1u*AY2�
��R�8�Q����RJ�J3�D}T� 85
Qg�/0 ��*A!P�*A�Ð𫿲��2ǿپ6t�6�=Q���Pȓ��� AQ� g�*ASt]1^u �ajrI�B����~�|0I�b��yI�\m�Qb�I�uz�A�c3Apa9q.� B6S��S��m����}�85`N�N�  �(M���f 1���6����161��55�s`�SC��U���A����5\setg06c����10�Fy�h8��a6��6��<9r�2HS ���Er���W@}�a��I�lB@���Y�ٖ�m�u� C����5�B��B��h`�F���X0���A:���C�M��AZ��@��4�6i����� e�O�-	���f1��F ��ᱦ�1F�Y	���T#6HL3��U66~`����U�dU�9D20L f0��Qv� ��fjq�� N������0v
� ��pi	�	��72lqQ�2������� \c�hngmove.�V��d���@2l_arf	�f~ ��6������9C�Z�`��~���kr41 S ���0��V��t���p���U�p7nuqQ`%�A]��V�1\�Qn�BJ�2W��EM!5���)�#:�6q4��F�e50S� \��0�=�PV���e ������E����޵�m7shqQSH"U��)��9�!A��(����� ,狟�ॲTR1�!��,�60e=�4�F�����2��	 R- ������������ ���4���LSR�)"�!lOA��Q�) ,%!� 16�
U/� �2�"2�E�9p���2X� SA/i��'�
7F�H�@!B�0��D ���5V��@2cVE֐�p��T��pt갖�1AL~E�#�F�Q��9E��#De/��RT��59 ���	�A�EiR������9\m20�2A0��+�-u�19r4�` �E1�=`O9`�1"ae��O�2��_$W.}am41�4�3�/~d1c_std��1)�!�`_T��r�_? 4\jdg�a�q �PJ%!~`-�r�+bpgB��#c300�"Y�5j�QpQb1�bq0��vB��v25�U��8����qm43� �Q <W�"PsA��e� ���t�i�P�W.� �c�FX.�e�k�E14�44�~67\j4�443sj<��r�j4up���\E19�h�PA�T�=:o �APf��coWo!\��2a��2A;_2��QW2�bF�(�V11�23�`��X5�Ra21�J*9�a:8�8J9X�l5�m1�a첚��*���(85 �&�������P6���R,52&A����q,fA9IfI50\u�z�OV
�v��}E֖aJ���Y>� 16r@�C�Y��;��1��L�� �Aq�&ŦP1��vB)�e�m�����1p�] �1D���27��F�KAREL U�se S��FCTyN��� J97�FA+�� (�Q޵�p�%�)?�Vj9F?(�j��Rtk208 "!Km�6Q�y�j��iÄ�Pr�9�s#��v�kwrcfp�RCFt3����Q��kcctme�!ME�g����6�main�dV�� ���ru��kDº�c`���o����J�dt�rF �»�.vrT�f�����E%�!��5�.FRj73B�K����UER�HJ�O  JF�� (ڳF���F�q �Y�&T��p�F�z��19�tkvBr���V�h�!9p�E�y�<�k�������;�v���"CT ��f����)�
І�� )�V	�6���!��q FF��1q���=����ҀO�?�$"���$��j�e���TCP Au�t�r�<520 H�5�J53E193Z��9��96�!8��q9��	 �B574��52�Je�(�� Se%!Y�����u��m|a�Pqtool����������con�rel�Ftrol� Reliabl�e�RmvCU!��H5�1����� a5�51e"�CNRE¹I�c�&��i�t�l\sfutst "UTա��"X�\u��g@�i�6Q"]V0�B,Eѝ6A� �Q�)C���X��Y�f�I�1|6s@6i��T6IU��vR�d��
$e%1��2�C58�E6��8�Pv�iV4OFFH58SOeJ� mvB7M6E~O58�I�0 �E�#+@�&�F�0�� �F�P6a���)/++�|</N)0\tr1��<���P ,��ɶ�r�maski�mskH�aA���ky'd�h	A�	�P�sDispl/ayIm�`v����?J887 ("A���+HeůצprdsP��Iϩǅ�h�0pl�E2�R2��:�Gt�@��PRD�TɈ�r�C��@Fm��D�Q�Asc	aҦ� V<Q&��bVvbrl�eې@���^S��&5Uf�j8710�yl	��Uq���7�&�p�p��P^@<�P�firmQ��ǀ�Pp�2�=bk�6�r�3x��6��tppl���PL���O�p<b�ac �q	��g1J�U�d�J��gait_9e���Y�&��Q���	�Sh�ap��erati�on�0��R67�451j9(`sGe�n�ms�42-f��r��p�5����2�rsg�l�E��p�G���qF�205p�5S���Ձ�r'etsap�BP�O��\s� "GCR��ö? �qngda��G��V��st2a�xU��Aa]��ba�d�_�btput�l/�&�e���tplcibB_��=�2.��8��5���cird�v��slp��x�hex���v�re?�Ɵx�k3ey�v�pm���x�us$�6�gcr���F������[�q27j�92�v�ollismqSk�9O�ݝ� (pl.���t��	p!o��29$Fo8���cg7no@�tptc;ls` CLS�o�b��\�km�ai_
�s>�v�o	�t�b����<��E�H��6�1�enu501�[m���utia|$ca�lmaUR��Cal�MateT;R51%�i=1]@-��/V� �@�Z�� �fq1�9 "K9E�L����2=m�CLMTq�S#f��et �LM3�!} �F�c�nspxQ�c���c_moq��� ��c_e�����#su��ޏ �_ �@�<5�G�join�i� j��oX���&cWv	� ���N�ve��C�c�lm�&Ao# �|$f�inde�0�STD ter �FiLANG4���R��
��n3���z0Cen���r,������J�����  ���K��Ú�=����_Ӛ��r� "F�NDR�� 3��f>��tguid�䙃0N�."��J�tq�� � ������������J����_������c��	�m�Z��\fnd�r.��n#>
B2p|��Z�CP Ma�����38A��� c��6� (���N�B������ 2�$�8�1��m_���"e x�z5�.Ӛ��c��`�bSа�efQ�p��	��RBT;�?OPTN �+# Q�*$�r*$��*$r*$ %/s#C�d/.,P�/0*>ʲDPN��$،��$*�Gr�$k �Exc�'IF�$M�ASK�%93 H�5�%H558�$5/48 H�$4-1�$���#1(�$�0 E��$��$-b�$���!UPDT �B�4�b�4�2�49�0�4a�3�9�j0"M�49�4  ��4�4tps�h���4�P�4- DQ� �3�Q�4�R�4�p�R%0�2�r�4.b
E\����5�A�4��3ad�q\�5K979"�:E�ajO l "DAQ^E^�3i�Dq �H�4ҲO ?R�? ���q�5��T��3rAq��O�Lst�5~��7p��5��REJ#�2�@av@^Eͱ�F���4��.�5�y N� �2il(�in�4��31 J0H1�2Q4�251ݠ�4Ormal� �3)� REo�Z_�æOx����4p��^F�?onorTf ��7_ja�UZҒ4l�5rmsAU�Kkg���4�$HCd\�fͲ�eڱH�4�REM���4yݱx"u@�RER5932f�O��47Z��5lit�y,�U��e"Di#l\�5��o ��7�987�?�25 �3hk910�3��FE��0=0P_�Hl\mhm�5��qe�=$�^��
E��u�IAymp�tm�U��BU��vste�y\�3��me�b� DvI�[�Qu�:F�Ub�`*_�
E,�su��_ Er��ox�<��4huse�E-�?�sn�������FE���,�box�����c ݌,"�������z���M��g��pdspw)�	��9���b���(��1���c ��Y�R�� �>�P����W��������'�0�ɵ�[��͂���  � ,�@�� �A�bWumpšf��B*��Box%��7Aǰ6�0�BBw���MC� (�6�,f�t I�s� ST��*��}B������w��"BBF
�>�`���)���\bbk968 a"�4�ω�bb��9va69����et�bŠ��X�����ed	�F��u�f� �sea"������'�\��,���b�ѽՑo6�H�
�x�$�f����!y���Q[�! �tperr�fd�� TPl0o� Recov,��3D��_R642 � 0��LC@}s� N@��(U�'rro���yu2r���  �
�  ����$$C�Le� ���t���������$z�?_DIGIT��������.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_� oo$j��+c:P�RODUCTM�0\PGSTKD��qV&ohozf99���D���$FE�AT_INDEX���xd���  
�`ILECOMP ;����#��`�cSETUP2 <�e��b�  N� �a�c_AP2B�CK 1=�i � �)wh0?{%&c����Q�xe %�I�m��� 8��\�n����!��� ȏW��{��"���F� Տj���w���/�ğS� ��������B�T�� x������=�үa��� ���,���P�߯t��� ���9�ο�o�ϓ� (�:�ɿ^���Ϗ� ��G���k� �ߡ�6� ��Z�l��ϐ�ߴ��� U���y����D��� h��ߌ��-���Q��� ������@�R���v� ���)�����_����� *��N��r� �7��m�&��3\�i
pP� 2#p*.VRc�*��0� /��PC/1/>FR6:/].��/+T�`�/�/�F%�/�,�`r/?�G*.F�8?	H#�&?e<�/�?;STM �2�?�.K �?�=�iPend�ant Pane	l�?;H�?@O�7.Op�?y?�O:GIF�O��O�5�OoO�O_:JPG _J_�56_�O_��_�	PANELO1.DT�_�0 �_�_�?O�_2�_So@�WAo�_o�o�Z3qo��o�W�o�o�o)�Z4 �o[�WI���
TPEINS.�XML��0\����qCusto�m Toolba�r	��PASS�WORDyF�RS:\L�� %�Passwor�d Config ���֏e�Ϗ�B0� ��T�f���������� O��s������>�͟ b��[���'���K�� 򯁯���:�L�ۯp� ����#�5�ʿY��}� �$ϳ�H�׿l�~�� ��1�����g��ϋ� � ����V���z�	�s߰� ?���c���
��.�� R�d��߈���;�M� ��q������<���`� �����%���I����� ���8����n�� �!��W�{ "�F�j|� /�Se��/� /T/�x//�/�/=/ �/a/�/?�/,?�/P? �/�/�??�?9?�?�? o?O�?(O:O�?^O�? �O�O#O�OGO�OkO}O _�O6_�O/_l_�O�_ _�_�_U_�_y_o o �_Do�_ho�_	o�o-o �oQo�o�o�o�o@ R�ov��;� _���*��N�� G������7�̏ޏm� ���&�8�Ǐ\�돀� �!���E�ڟi�ӟ� ��4�ßX�j������ ��įS��w�������B�#��$FILE�_DGBCK 1�=��/���� ( ��)
SUMMAR�Y.DGL���M�D:�����D�iag Summ�ary��Ϊ
CONSLOG��������D�ӱConsole logE��ͫ��MEMCH�ECK:�!ϯ����X�Memory �Data��ѧ��{)��HADO�W�ϣϵ�J���S�hadow Ch�angesM�'�-���)	FTP�7Ϥ�3ߨ���Z�m�ment TBD���ѧ0=4)ETHERNET��������T�ӱEthernet \��figurati�onU�ؠ��DCSVRF�߽߫������%�� verify all���'�1PY���DI�FF�����[���{%��diff]������1R�9�K���� ���X��CHGD�������c��r����2pZAS� ��GD���k���z��FY3pbI[� �/"GD���s/�����/*&UP?DATES.� �/~��FRS:\�/��-ԱUpdates List�/���PSRBWLD'.CM(?���"<?��/Y�PS_ROBOWEL��̯�?�? ��?&�O-O�?QO�? uOOnO�O:O�O^O�O _�O)_�OM___�O�_ _�_�_H_�_l_o�_ �_7o�_[o�_lo�o o �oDo�o�ozo�o3 E�oi�o��� R�v���A�� e�w����*���я`� ��������O�ޏs� �����8�͟\��� ��'���K�]�쟁�� ��4���ۯj������ 5�įY��}������ B�׿�x�Ϝ�1��� *�g�����Ϝ���P� ��t�	�ߪ�?���c� u�ߙ�(߽�L߶��� ����(�M���q� � ���6���Z������ %���I���B������2�����h����$�FILE_� PR�� ��������MDONLY 1=.~�� 
 ��� q���������� ~%�I�m �2��h�� !/�./W/�{/
/�/ �/@/�/d/�/?�//? �/S?e?�/�??�?<? �?�?r?O�?+O=O�? aO�?�O�O&O�OJO�O �O�O_�O9_�OF_o_~
VISBCKL|6[*.VDv_|�_.PFR:\�_��^.PVisi�on VD file�_�O4oFo\_jo T_�oo�o�oSo�owo �oB�of�o �+������ �+�P��t������ 9�Ώ]�򏁏��(��� L�^�������5��� ܟk� ���$�6�şZ���~�����
MR_GRP 1>.�L��C4  ;B���	 W������*u����RHB ���2 ��� �?�� ���B��� ��Z�l���C���D������Ŀ��K�E�jJ�d5I��(T�N8F�5UP��* ���ؿ�E�M.G��E$��;n߇�:G��@O����@��
@�f��fe@�k�@�H~*λ� F@ ��������J��NJk��H9�Hu���F!��IP��s�?����(�9��<9�8�96C'6<?,6\b��+�@&�(�a�L߅�p�A��A��߲�v���r��� ���
�C�.�@�y�d� �������������`�?�Z�lϖ�BH�� �Ζ��������
0�PS@�P��Rh��ܿ� �B�x��/ ��@�33:���.�gN�UUU�U��q	>u.�?!rX���	�-=[z��=�̽=V6�<�=�=��=$q�����@�8�i7G���8�D�8@9!�7�:�����D�@ D�Ϡ Cϥ��C�
�����'/0-��P/ ����/N��/r��/�� �/�??;?&?_?J? \?�?�?�?�?�?�?O �?O7O"O[OFOOjO �O�O�O�O�гߵ��O $_�OH_3_l_W_�_{_ �_�_�_�_�_o�_2o oVohoSo�owo�o�i ��o�o�o��); �o_J�j��� ����%��5�[� F��j�����Ǐ��� ֏�!��E�0�i�{� B/��f/�/�/�/���/ ��/A�\�e�P���t� �������ί��+� �O�:�s�^�p����� Ϳ���ܿ� ��OH� �o�
ϓ�~ϷϢ��� �������5� �Y�D� }�hߍ߳ߞ������� �o�1�C�U�y��� ������������� -��Q�<�u�`����� ����������; &_J\����� �����ڟ�F� j4������� ��!//1/W/B/{/ f/�/�/�/�/�/�/�/ ??A?,?e?,φ?P� q?�?�?�?�?O�?+O OOO:OLO�OpO�O�O �O�O�O�O_'__K_ �o_�_�_�_l��_0_ �_�_�_#o
oGo.oko Voho�o�o�o�o�o�o �oC.gR� v�����	�� �<�`�*<��` �����ޏ��)�� M�8�q�\�������˟ ���ڟ���7�"�[� F�X���|���|?֯�? �����3��W�B�{� f�����ÿ������� ��A�,�e�P�uϛ� b_�����Ϫ_��߀� =�(�a�s�Zߗ�~߻� ��������� �9�$� ]�H��l������ ������#��G�Y� � B�������z������� 
ԏ:�C.gRd ������	� ?*cN�r� ����/̯&/� M/�q/\/�/�/�/�/ �/�/�/?�/7?"?4? m?X?�?|?�?�?�?�? ��O!O3O��WOiO�? �OxO�O�O�O�O�O_ �O/__S_>_P_�_t_ �_�_�_�_�_�_o+o oOo:oso^o�o�op� �o�� ��$�� o�o�~��� ����5� �Y�D� }�h�������׏�� ��
�C�.�/v�<� ��8������П��� �?�*�c�N���r��� �����̯��)��? 9�_�q���JO����� ݿȿ��%�7��[� F��jϣώ��ϲ��� ����!��E�0�i�T� yߟߊ��߮��߮o�o ��o>�t�>�� b�����������+� �O�:�L���p����� ��������'K 6oZ�Z�|�~�� ���5 YD i�z����� �/
//U/@/y/@� �/�/�/�/���/^/? ??Q?8?u?\?�?�? �?�?�?�?�?OO;O &O8OqO\O�O�O�O�O��O�O�O_�O7_���$FNO ����VQ_�
F0fQ kP� FLAG8�(�LRRM_CHKT_YP  WP��^P�WP�{QO=M�P_MIN�P�����P�  �XNPSSB_CF�G ?VU ��_���S� ooIUTP_DEF_OW  ���R&hIRCOM��P8o�$GENO�VRD_DO�V��6�flTHR�V �d�edkd_ENB�Wo k`RAVC_GRP 1@�WCa X"_�o_ 1U<y�r� ����	��-�� =�c�J���n������� �ȏ����;�"�_�pF�X���ibROU�`�FVX�P��&�<b&�8�?���埘�������  D?�јs���@@g�B�7�p�)�ԙ���`SMT�cG��mM���� �LQHoOSTC�R1H����P��at�S5M��f�\���	127.0��=1��  e��ٿ �����ǿ@�R�d��vϙ�0�*�	ano?nymous���������z��[�� � �����r����� �ߺ�����-���&� 8�[�I�π���� ��1�C��W�y� ��`�r������ߺ��� ����%�c�u�J\ n�������� �M�"4FX��i ������7/ /0/B/T/���m/ ��/�/�/??,? �/P?b?t?�?�/�?� �?�?�?OOe/w/�/ �/�?�O�/�O�O�O�O �O=?_$_6_H_kOY_ �?�_�_�_�_�_'O9O KO]O__Do�Ohozo�o �o�o�O�o�o�o
 ?o}_Rdv���_ �_oo!�Uo*�<� N�`�r��o������̏ ޏ�?Q&�8�J�\����>�ENT 1I��� P!􏪟  ����՟ğ�� �����A��M�(�v� ��^�����㯦��ʯ +�� �a�$���H��� l�Ϳ�����ƿ'�� K��o�2�hϥϔ��� ���ϰ�������F� k�.ߏ�R߳�v��ߚ� �߾���1���U��y��<�QUICC0 ��b�t����1�����%���2&���u��!ROUTER�v�R�d���!PC�JOG����!�192.168.�0.10��w�NA�ME !��!�ROBOTp�S_CFG 1H��� �A�uto-star�ted�tFTP�������  2D��hz� ���U��
// ./�v���/�� �/�/�/�/�/�!?3? E?W?i?�/?�?�?�? �?�?�?���AO�? eO�/�O�O�O�O�?�O �O__+_NO�OJ_s_ �_�_�_�_
OO.Oo B_'ovOKo]ooo�oP_ >o�o�o�o�oo�o 5GYk}�_�_�_ ��8o��1�C� U�$y��������ӏ f���	��-�?��� ��Ə���ϟ�� ���;�M�_�q��� .�(���˯ݯ��P� b�t�����m������� ��ǿٿ�����!�3� E�h��{ύϟϱ��� �$�6�H�J�/�~�S� e�w߉ߛ�jϿ����� ���*߬�=�O�a�s����YT_ERR �J5
���PDU�SIZ  ��^�J����>��WR�D ?t�� � guest}��%�7�I�[��m�$SCDMNG�RP 2Kt������V$��K�� 	P0�1.14 8�� _  y�����B    �;����� ���������
 �������������~����C.�gR|���  �i  �  k
�������� �+�������_
���l .r+���"�l��� m
d������__GROU��L�� �	����0�7EQUPD  �	պ�J�TY�a ����TTP�_AUTH 1M��� <!iP�endany���6�Y!KAR�EL:*��
-�KC///A/ V�ISION SE!TT�/v/�"�/ �/�/#�/�/
??Q?�(?:?�?^?p>�CTRL N����5��
�FFF�9E3�?�FR�S:DEFAUL�T�<FANU�C Web Se/rver�:
��� ��<kO}O�O�O�O�O���WR_CONF�IG O�� ��?��IDL_C_PU_PC@�sB��7P�BHU�MIN(\��<TGNR_IO�������PNPT_SIM�_DOmVw[TPMODNTOLmV} �]_PRTY�X�7RTOLNK 1P����_o!o3o�EoWoio�RMAST�ElP��R�O_C3FG�o�iUO��o>�bCYCLE�o�d�@_ASG 1Q����
 ko,> Pbt����������sk�bNU�M����K@�`IP�CH�o��`RTRY_CN@oR��b�SCRN����Q�b�� �b�`�bR����Տ��$J23_DSP_EN	�����OBPR�OC�U�iJOG�P1SY@��8��?�!�T�!�?>*�POSRE�zV?KANJI_�`��o_�� ��T�L�6x͕����CL_LGP�<�_���EYLOGWGIN�`����LANGUAGgE YF7RDY w���LG��U�?V⧈�x� ���j��=P��'0����$ NMC:�\RSCH\00�\��LN_DISP V��
���������OC�R.RDz�VTA{�OGBOOK W
{��i��ii��X����� ǿٿ�����"��6	h�����e��?�G_BUFF K1X�]��2	� �ϸ���������� �!�N�E�W߄�{ߍ� �߱�����������J���DCS }Zr� =���� ^�+�ZE��������a��IO 1[
{ ُ!� �!�1�C� U�i�y����������� ����	-AQc�u�������E^fPTM  �d�2 /ASew�� �����//+/ =/O/a/s/�/�/���SEV����TYP�/??y͒�RS@"��×��FL 1\
������?�?�?�?�?�?L�?/?TP6��"}>�NGNAM�ե�U`�UPS��G�I}�𑪅mA_L�OAD�G %��%DF_MO�TN���O�@MAXUALRM<��J� �@sA�Q����WS �
�@C �]m�-_���M�P2�7�^
{ �Z��	�!P�+ʠ1�;_/��Rr�W�_�WU�W�_��R	o �_o?o"ocoNoso�o �o�o�o�o�o�o�o ;&Kq\�x� ������#�I� 4�m�P���|���Ǐ�� �֏��!��E�(�i� T�f�����ß��ӟ�� �� �A�,�>�w�Z� ������ѯ����د� ��O�2�s�^����� ��Ϳ���ܿ�'��B�D_LDXDIS�AX@	��MEMO�_APR@E ?�+
 � *�~� �Ϣϴ����������@�ISC 1_�+ ��IߨT��Q�c� Ϝ߇��ߧ�����w� ���>�)�b�t�[�� ��{���������� :���I�[�/������ ������o�����6! ZlS��s� ���2�AS '�w����g���.//R/d/�_MSTR `�-~w%SCD 1am��L/�/H/�/�/?�/ 2??/?h?S?�?w?�? �?�?�?�?
O�?.OO RO=OvOaO�O�O�O�O �O�O�O__<_'_L_ r_]_�_�_�_�_�_�_ o�_�_8o#o\oGo�o ko�o�o�o�o�o�o�o "F1jUg� �������� B�-�f�Q���u������ҏh/MKCFG �b�-㏕"LT�ARM_��cL�;� σQ�|N�<�METPUI��ǂ���)NDS?P_CMNTh��8�|�  d�.���ς�ҟܔ|�PO�SCF����PS�TOL 1e'�4=@�<#�
5�́ 5�E�S�1�S�U�g��� ����߯��ӯ���	� K�-�?���c�u������|�SING_CH�K  ��;�ODAQ,�f��Ç��DEV 	L�	�MC:!�HSI�ZEh��-��TA�SK %6�%$�12345678�9 �Ϡ��TRI�G 1g�+ l6�%���ǃ����ό8�p�YP[� ��E�M_INF 1h�3� `�)AT&FV0�E0"ߙ�)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ������H�� ���A���AI�q� ,��|���� ��� �ߵ�����J���n��� ����W����������� "����X��/�� ��e������0 �T;x�=�a s��/�,/c=/ b/�/A/�/�/�/�/ ��?���^?p? #/�?�/�?s?}/�?�? O�?6OHO�/lO?1? C?U?�Oy?�O�O3O _ �?D_�OU_z_a_�_玿ONITOR��G� ?5�   	?EXEC1Ƀ�RU2�X3�X4�X5�XT���V7�X8�X9Ƀ�RhBLd�RLd�RLd �RLd
bLdbLd"bLd@.bLd:bLdFbLc2ShU2_h2kh2wh2�hU2�h2�h2�h2�hU2�h3Sh3_h3�R��R_GRP_SOV 1in���(�����C?BPP��A4�>%���gY�>rﳌ�x�_D=R^��P�L_NAME �!6��p�!D�efault P�ersonali�ty (from� FD) �RR�2eq 1j)TU�X)TX��q��X dϏ8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|������2'�П�����@*�<�N�`�r��<�� ������ү������,�>�P�b� �Rdr �1o�y �\�,� �3���� �@D�  ��?�ĸ���?䰺��A'�6����;�	�lʲ	 ��xJ������ �<w �"�� �(���pK�K ���K=*�J����J���JV�`��Z�����r���́p@j�@T;;f���f��ұ�]�l��I���������������b��3��´  ��`�>����b����z��ꜞ����Jm��
� B�H�˱]���q��	� p�  �P�pQ�p��p|  Ъ�g���c�	'� � ���I� �  �����:�È~
�È=���"��nÿ�	�ВI  ?�n @B�c���\��ۤ��q�y��o�N���  '������@2��@Ǔ����/�C���C�C�@ C�������
��A�W�@<�P�JR�
h�B�b�A�Єj�����:��Dz۩��߹������j��( �� -��C���'�7�����q�Y������ �?�ff� ��gy ����o�:a�:�
>+�  PƱj�(����7	�ü�|�?����x�Z�p<
6b<�߈;܍�<��ê<� <�#&Jσ�AI�ɳ�+���?fff?�I�?&�k�@�.���J<?�`�q�.�˴fɺ� /��5/����j/U/ �/y/�/�/�/�/�/?0�/0?q��F�? l??�?/�?+)�?�?~�E�� E�I�?G+� F��? )O�?9O_OJO�OnO�Of�BL޳B�?_h� .��O�O��%_�OL_�? m_�?�__�_�_�_�_��
�h�Îg>��_Co�_goRodo�o�GA�ds�q��C�o�o�o|���A�$]Hq���D���pC���pC!HmZZ7t���6q�q���ܶN'�3A��A�AR1AO��^?�$�?��K/�±
=���>����3�?W
=�#�W���e��9������{����<�����(�B�u���=B0������	L���H�F�G����G��H�U�`E���C�+����I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3�l� W���{��������՟ ���2��V�A�z��� w�����ԯ������ ��R�=�v�a����� �������߿��<� '�`�Kτ�oρϺϥ� �������&��J�\� G߀�kߤߏ��߳��� ����"��F�1�j�U� ��y���������� ��0��T�?�Q�����(���3/E�y���u����<��q3�8�����q4Mgs&�IB+2D�a���{�^^	�@�����uP2	P7Q4_A��M00bt��R��`����/   �/�b/P/�/t/�/  *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?��?�?O 2 F;�$�vGb�/�Aa��@�a�`�qC��C�@�o�Ot���KF�� DzH@�� F�P D���O�O�ys<O!_3_E_�W_i_s?���@U@pZ�422�!2~
  p_�_�_�_	oo-o?o Qocouo�o�o�o�o��Q ��+��1���$MSKCF�MAP  �5?� �6�Q��Q"~�cONREL7  
q3��bEXCFENB�?w
s1uXqFNC�_QtJOGOVLKIM?wdIpMrd�bWKEY?w�u�bWRUN�|�u�bSFSPDTY�xavJu3sSIGN?>QtT1MOT�Nq��b_CE_GRoP 1p�5s\r���j�����T�� ⏙������<��`� �U���M���̟��� ���&�ݟJ��C��� 7�������گ��������4�V�`TCOM_CFG 1q}��Vp�����
P�_/ARC_\r
jyUAP_CPL���ntNOCHECK� ?{  	r��1�C�U�g� yϋϝϯ����������	��({NO_WA�IT_L�	uM�NMTX�r{�[m�o_ERRY�2sy3� &��������r�c� ��T_�MO��t��,  �E�$�k�3�PAR�AM��u{��	�[���u?�� =�9@345678901��&���E�W� 3�c�����{������������=��UM_RSPAC�E �Vv��$ODRDSP���jx�OFFSET_C�ARTܿ�DIS���PEN_FI�LE� �q��c֮�O�PTION_IO���PWORK kv_�ms � P(�R�Q
�j.j�	 ��Hj&6$�� RG_DSBL'  �5Js�\���RIENTTO>p9!C��PqfA�� UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?p]a]�D�WcUa쪋l;�	�lmb�`�x7J�`�p����a�< ���`� ��b��H(���H3k7HS�M5G�22G�?��Gp
��
�ƨ��'|��CR�>�>q�GsuaT��3���  �4spBpyr  ]o��*SB_����=j]��t�q� ��rna �,��~�6  ��UPQ�|N��M�,k���	'�� � ��I�� �  ��%�=��ͭ����ba	���I  �n @��~����p�������N	 W�  '!o�:q:�pC	 C�@@sBq��|��� m�
�T!�h@ߐ�n��$��*�B	 �A����p� �-�qbz ��P��t�_�������( �� -��恊�n�ڥD[A]Ѻ�b4�'!5�~(p �?�ff� ��
����OZ�R�*�85�z���>΁  Pia��(5���@����ک�a�c�dF#?˙�5�x��*�<
�6b<߈;����<�ê<�? <�&�o&ς)�A�lcΐI�*�?offf?�?&c�ޒ�@�.uJ<?�`��Yђ ^�nd��]e��[g��G� �d<����1��U�@� y�dߝ߯ߚ����߼� 	���-������&��~"�E�� E��?G+� Fþ��� ��������&��J�(5��bB��AT�8� ђ��0�6���>���J� n�7��[m��0��h��1��>�M�I
�@��A�[���C-�)��?Ƀ��� /�Y���Jp��vav`CH�/������}!@�I�Y�'�3A��A�AR1A�O�^?�$�?�����±
=�ç>����3�W
=�#�����+e��ܒ������{����<���.(�B��u��=B0�������	��*H�F�G����G��H��U`E���C��+�-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�? O�?3OOWOBOTO�O xO�O�O�O�O�O�O_ /__S_>_w_b_�_�_ �_�_�_�_�_oo=o (oaoLo�o�o�o�o�o �o�o�o'$] H�l����� ��#��G�2�k�V� ��z���ŏ���ԏ� ��1��U�g�R���v� ����ӟ�������-�:�(���������a����xQ�c�,!3�8�}�<��,!4Mgs�����ɢIB+կ篴a?���{����A�/�e�S���w��P!�P�������7�`�ӯ�ϑ�R9��Kτ�oχϓϥ�  ���χ����)�� M������z���{߉�����ߒߤ�������  )�G�q��_���2 wF�$�&Gb����n�[ZjM!C��s�@j/�A�S�=�F�� Dz���� F�P D��W����)������������x?��ͫ@@
9�=��=��=��
 v����� ��*<N`ܷ*P ���˨��1��$PARA�M_MENU ?�-�� � DEF�PULSEl	�WAITTMOU�T�RCV� �SHELL_�WRK.$CUR�_STYL��,OPT�/PT�B./("C�R_DECSN���,y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?��USE_PROG %�%�?�?�3CCR�����7�_HOST !F�!�44O�:T̰�?PCO)ARC�O�;_TIME�XB��  �GDEB�UGV@��3GINP_FLMSK�O��IT`��O�EPGA�P �L��#[CH��O�HTYPE����?�?�_�_�_�_ �_oo'o9obo]ooo �o�o�o�o�o�o�o�o :5GY�}� ���������1�Z��EWORD �?	7]	RS�`�	PNS��$��JOE!>�T�Es@WVTRACE�CTL 1x-�]� ������ɆDT Q�y-���D 7� ��,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�T�(� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ j��_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�_����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v��������//"#�$PGT�RACELEN � #!  ���" �8&_�UP z��e�g!o S!h �8!_CFG {Fg%Q#"!x!�$�J �#|"DEFSP/D |�,!!J ��8 IN TR�L }�-" 8��%�!PE_CON�FI� ~g%��g!�$�%�$L�ID�#�-74G�RP 1�7Q!��#!A ����&ff"!A+33�D�� D]� ?CÀ A@+6�!�" d�$�9�9*1*0?� 	 +9�(8�&�"�? ´	C�?�;B@3AO�?OIO�3OmO"!>�T?��
5�O�O�N�O �=��=#�
 �O_�O_J_5_n_Y_��O}_�_y_�_�_�_ G Dzco" 
o Bo�_Roxoco�o�o�o �o�o�o�o>)�bM��;
V7�.10beta1��$  A��E�rӻ�A �" �p?!G��q>����r��0�q{�ͻqBQ��q�A\�p�q�4�q�p
�"�BȔ2�D�V��h�w��p�?�?)2 {ȏw�׏���4� �1�j�U���y����� ֟������0��T� ?�x�c�������ү�� ��!o�,�ۯP�;�M� ��q�����ο���ݿ �(��L�7�p�+9��sF@ �ɣͷ� ��g%������+�!6 I�[߆������ߵߠ� ��������!��E�0� B�{�f�������� �����A�,�e�P� ��t���������� ��=(aL^� ������' 9$]�Ϛ��ϖ� ������/<�5/`� r߄ߖߏ/>�/�/�/ �/�/?�/1??U?@? R?�?v?�?�?�?�?�? �?O-OOQO<OuO`O �O�O�O�O���O_�O )__M_8_q_\_n_�_ �_�_�_�_�_o�_7o Iot���o�o�� �o�o�o(/!L/^/p/ �/{*o����� ����A�,�e�P� b����������Ώ� �+�=�(�a�L���p� �����Oߟ񟠟� � 9�$�]�H���l�~��� ��ۯƯ���#�No`o ro�on��o�o�o�oԿ ���8J\ng� ���vϯϚ������� 	���-��Q�<�u�`� r߫ߖ��ߺ������ �;�M�8�q�\���� ����z������%�� I�4�m�X���|����� ������:�L�^��� Z���������� �$�6�H�Sw b������� //=/(/a/L/�/p/ �/�/�/�/�/?�/'? ?K?]?H?�?��?�? f?�?�?�?O�?5O O YODO}OhO�O�O�O�O �O�O&8J4_F_� ���_�_��_�_ "4-o�O*ocoNo�o ro�o�o�o�o�o�o )M8q\�� �������7� "�[�m��?����R�Ǐ ���֏�!��E�0� i�T���x�������� _$_V_ �2�l_~_�_������R�$PLI�D_KNOW_M�  �T������SV ��U͠�U��
��.�ǟR��=�O�����mӣM_?GRP 1��!`U0u��T@ٰo�
ҵ�
���Pзj� �`���!�J�_�W� i�{ύϟϱ�������X��߱�MR�����1T��s�w� s��� �޴߯߅��ߩ߻��� ��A���'���� �����������=� ��#���������}�������S��ST��1W 1��U# ���;0�_ A .�� ,>Pb���� ����3(i L^p������2*���	<-/3/)/;/M/�4f/x/�/�/5 �/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?M_AD  d#�`PARNUM  w�%OWSCH?J ME
�Gp`A�Iͣ�EUPD`O�rE
a�OT_CM�P_��B@�P@'�˥TER_CHK'U��˪?R$_6[�RSl�¯��_MO�A@�_�U_�_RE_R/ES_G �� >�oo8o+o\oOo�o so�o�o�o�o�o�o�o�W �\�_%�U e Baf�S� �� ��S0����SR0 ��#��S�0>�]�b���S�0}������RV �1�����rB@c]���t�(@c\�����D@c[��$���RTHR_�INRl�DA��˥d�,�MASS9� Z�M�MN8�k�MON�_QUEUE a���˦��x� RDNPUbQN{�P[���END���_ڙEX1E�ڕ�@BE�ʟ>��OPTIOǗ�[���PROGRAM7 %��%��ۏ��O��TASK_I�AD0�OCFG ኞ�tO��ŠDATuA���Ϋ@��27�>�P�b�t���,� ����ɿۿ�����#�x5�G���INFOU���������ϭϿ� ��������+�=�O� a�s߅ߗߩ߻���������^�jč� �yġ?PDIT �ίc���WERF�L
��
RGADoJ �n�A��¹�?����@���IOORITY{�QV���MPDSPH������Uz����OTO�Ey�1�R� (/!AF4�E�P]�~��!tcph�>��!ud��!icm��ݏ6�XY_ȡ�R�=�ۡ)� *+/ ۠�W:F �j����� �%7[B�=*��PORT#�BC�۠����_C?ARTREP
�R�> SKSTAz��Z�SSAV���n�	�2500H86A3���r�$!�R����q�n�}/x�/�'� URGE��B��rYWF� DO{�rUVWV��$�A��WRUP_DEL�AY �R��$RO_HOTk��%O�]?�$R_NORM�ALk�L?�?p6SE�MI?�?�?3AQS�KIP!�n�l#x 	1/+O+ O ROdOvO9Hn��O�G�O �O�O�O�O_�O_D_ V_h_._�_z_�_�_�_ �_�_
o�_.o@oRoo vodo�o�o�o�o�o�o �o*<Lr`���n��$RCgVTM�����p�DCR!�L���qB��C*J��C$�>�$� >5?-;���04M¹�O���ǃ��������~��9On�Y�<
�6b<߈;����>u.�??!<�&{�b� ˏݏ��8�����,� >�P�b�t��������� Ο���ݟ��:�%� 7�p�S������ʯܯ � ��$�6�H�Z�l� ~�������ƿ���տ ���2�D�'�h�zϽ� �ϰ���������
�� .�@�R�d�Oψߚ߅� �ߩ���������<� N��r������� ������&�8�#�\� G�����}��������� ��S�4FXj| ������� ��0T?x�u ����'//,/ >/P/b/t/�/�/�/�/ �/�/�?�/(??L? 7?p?�?e?�?�?��? �? OO$O6OHOZOlO ~O�O�O�?�?�O�O�O �O __D_V_9_z_�_ �?�_�_�_�_�_
oo�.o@oRodovo�X�qG�N_ATC 1��� AT�&FV0E/� �ATDP/6/�9/2/9�hA�TA�n,A�T%G1%B96}0/�+++�o�,�aH,�qIO�_TYPE  �u�sn_�oREFPOS1 1�P{� x�o�X h_�d_����� K�6�o�
���.���R�x���{{2 1�P{���؏V�ԏz����q3 1��$�6��p��ٟ���S4 1�����˟���n�|��%�S5 1�<��N�`�����<���S6 1�ѯ���/�𭿘�ѿO�S7 1�f�x���ĿB�-�f�>�S8 1������Y�������y�SM�ASK 1�P � 
9�G��XNO�M���a~߈ӁqMOTE  h�~t��_CFG �������рrPL_RA�NG�ћQ��POW_ER ��e����SM_DRYP_RG %i�%���J��TART ��
�X�UME_P�RO'�9��~t_E�XEC_ENB � �e��GSPD�������c��TDB����RM��MT�_!�T���`O�BOT_NAME� i���iO�B_ORD_NU�M ?
�\q�H863  a�T��������b�PC_TIMEO�UT�� x�`S2�32��1��k �LTEACH PENDAN ��ǅ�}���`�Maintena�nce ConsțR}�m
"{�dKCL/Cg��Z ���n� No Use}�	���*NPO��х����(CH_�L�������	��mMAVAILȰ�{��ՙ�SPACE1 2��| d��(>���&���p��M,8�?�ep/eT/ �/�/�/�/�W//,/ >/�/b/�/v?�?Z?�/ �?�9�e�a�=??,? >?�?b?�?vO�OZO�?��O�O�Os�2� /O*O<O�O`O�O�_��_u_�_�_�_�_[3 _#_5_G_Y_o}_�_ �o�o�o�o�o[4.o@oRodovo$�o �o����"�	�7�[5K]o��A� ���	�̏�?�&�T�[6h�z������� ^�ԏ���&��;�\�C�q�[7�������� ͟{���"�C��X�y�`���[8����Ư دꯘ��0�?�`�#��uϖ�}ϫ�[G ��i� �ϋ
G� ����$�6� H�Z�l�~ߐ��8 ǳ�@����߈��d(� ��M�_�q���� ��������?���2� %�7�e�w��������� �����������!�R E�W�����������?Q; `�� @0�@�ߖrz	�V_ �����
/L/^/ |/2/d/�/�/�/�/�/ �/?�/�/�/*?l?~? �?R?�?�?�?�?�?�?�?2O�?
��O[�_MODE  ��˝IS ���vO,*ϲ�O-_���	M_v_#dCWO�RK_AD�M\{1�%aR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/$��:	d/JaR��WY��^���^R�^	r  P��� �  8��P�	�D��GYk}�� ������Qp/@/R//)P;�o\T��Q�pg-�t�_�DiKT��[  � lv%������/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OWW�#�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_olO~O d+No`oro�o�o�o�o �o�o�o&8J \n������u�  0�"0g�/� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q�����$o��˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�����Do ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������w
�  58�J�\�n߀� �ߜկ���������	� �-�?�Q�c�u������ ��-�� ��� �2�D�V�h�z���������������v���& ���%	12345�678�" 	�
�/� `r�������� (:L^p�� ����� //$/ 6/H/Z/l/~/��/�/ �/�/�/�/? ?2?D? V?h?�/�?�?�?�?�? �?�?
OO.O@Oo?dO vO�O�O�O�O�O�O�O __*_YON_`_r_�_ �_�_�_�_�_�_oo C_8oJo\ono�o�o�o �o�o�o�oo"4 FXj|���������	��s�3�E�W�{�Cz � Bp��   ��2���z�$S�CR_GRP 1��(�U8(�\�x^ @�  �	!�	 ׃���"� $� ��-��+��R�nw����D~������#����O����M-10iA 78909905 Ŗ~5 M61C >P4��Jׁ
� ���0�����#�1�	"�z�������4¯Ҭ ���c� ��O�8�J��� ����!�����ֿ��B�y�������r��A��$�  @���<� �R�?��d���H�y�u�O���F@ F�`�§�ʿ�϶� ������%��I�4�m� �<�l߃ߕߧ߹�B���\����1�� U�@�R��v����� �������;���*<=�
F���?�d�<��>7�����@��:��� B����ЗЙ���EL_D�EFAULT  ������B�MIPOWERFL  �x$1 WFDO� $��ERVE�NT 1������"�pL!D?UM_EIP��8���j!AF_I�NE �=�!FIT���!���4 ��[!�RPC_MAIN�\>�J�nVI�Sw=���!�TP�PU��	d��?/!
PMON?_PROXY@/�Ae./�/"Y/�fz/��/!RDM_S�RV�/�	g�/#?!#R C?�h?o?K!
pM�/�i^?��?!RLSYN�C�?8�8�?O!�ROS�.L�4 �?SO"wO�#DOVO�O �O�O�O�O_�O1_�O U__._@_�_d_v_�_ �_�_�_o�_?ooco�iICE_KL �?%y (%SVCPRG1ho 8��e���o�m3�o�o"�`4 �`5(-"�`6PU�`7x}��`���l9��{ �d:?��a�o��a�o E��a�om��a���a B���aj叟a�� �a�5��a�]��a� ���a3����a[�՟�a �����a��%��aӏM� �a��u��a#����aK� ů�as���a��mob �`�o�`8�}�w����� ��ɿ���ؿ���5� G�2�k�VϏ�zϳϞ� ���������1��U� @�y�dߝ߯ߚ��߾� ������?�*�Q�u� `���������� ��;�&�_�J���n������������sj_�DEV y	��MC:�ջ_OUT"�,REC 1q�Z� d   w 	�    ��@��� ���A�����
 �PSD#O6 r��O� ��� �� `�� ��Z�{� �� �*�  +X- � I- �- !- �� �X�YZ�PS�J;4 �?j  (�  Q� ��R ���� E- � b�/e/�l4H�/��� X� (�,/>/P/�/�/�""J4� =�!� � ؀  ?"S1��Z'!�/���("- ��\?�?$=�=�?�? �?"OOFO4OjO|O^O �O�O�O�O�O�O�O_  __T_B_x_f_�_�_ �_�_�_�_�_ooo Po>oto�oho�o�o�o �o�o�o(
L:�\�p���w ,����4�"�X� F�|���p�����֏ď ����0��@�f�T� ��x�����ҟ�Ɵ� ��,��<�b�P���h� z������ί��(� :��^�L�n�p����� ��ܿ�п� �6�$� Z�H�jϐ�rϴϢ��� �������2�D�&�h� Vߌ�z߰ߞ������� ����
�@�.�d�R��ZjV 1�w �P����j 
?�� ����
�TYPEVFZ�N_CFG ��5d�4�?GRP 1�A�c/ ,B� A� �D;� B����  B4R�B21HELL":�(
��?���<%RS'!�� H3lW�{� �����2XVh������%w����#!0�1�����7��2�0d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he��_ &_8_J_\_B_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}4xcopy �fr:\*.* �virt:\tm�pback�Q=>�192.168.�4�P46:165�2 �R�_�_�_�K}5�Ua�_�_�V�_go�yo�o}9�Ts:o�rderfil.dat.l@oVo�o�o�}0�Rmdb: +o�o�R�ocu�b �_2o?U��
�o���Sod�v����
�xyzrate 61 +�=�O�����������5012 ��ҏc�u����o �o56�ٟ���"���5�џb�t����6ܠ���emp:�81�88 W������.��*.d��Ʈϯ`�r�����1 +�=�O� ����)�Ҳ��ҿ c�uχϚ���5�ͧ�� �����"���̩��c� u߇ߚ����R�U��� ��
������T���h� z��ϱ�:������� 
�߸�A���d�v��� ��.�;�������� ����O�`r���� 2������'�� K�\n�����8�� ���#�G/ j/|/����3/E/W/�/��/�/��w2244 ?��/b?t?�?��4 58�?�?�?"�?58 �?bOtO�O���?���p9120 WO�O�O �O��O�J�Oa_s_�_ �/��<_N_�_�_o? (?�S�_�_couo�o�? �?5O�G�o�o�oO"O �o�H�obt���/ �/QcU��
�/� �Nq�h�z���o�o :����
���A�ӏd�v������$S�NPX_ASG �1�������� P 0� '%R[?1]@1.1����?���%֟��&� 	��\�?�f���u��� �����ϯ��"��F� )�;�|�_�������ֿ ��˿���B�%�f� I�[Ϝ�Ϧ��ϵ��� ����,��6�b�E߆� i�{߼ߟ�������� ���L�/�V��e�� �����������6� �+�l�O�v������� ��������2V 9K�o���� ���&R5v Yk�����/ ��<//F/r/U/�/ y/�/�/�/�/?�/&? 	??\???f?�?u?�? �?�?�?�?�?"OOFO )O;O|O_O�O�O�O�O �O�O_�O_B_%_f_ I_[_�__�_�_�_�_ �_�_,oo6oboEo�o io{o�o�o�o�o�o �oL/V�e� �������6� �+�l�O�v��������PARAM ������ �	U��P�����OFT_KB_CFG  ⃱����PIN_SIM  ���C�U�g������RVQSTP/_DSB,�򂣟|����SR �/��� &  AR������TOP__ON_ERސ����PTN �/�@�A�	�RING_PR�M� ��VDT_GRP 1�ˉ�  	������ ������Я����� *�Q�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߣߠ߲������� ����0�B�i�f�x� ������������� /�,�>�P�b�t����� ����������( :L^p���� ��� $6H Z�~����� ��/ /G/D/V/h/ z/�/�/�/�/�/�/? 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_�__\_��VPRG_�COUNT��8@���RENBU��U�M�S��__UPD� 1�/�8  
s_�oo*oSoNo `oro�o�o�o�o�o�o �o+&8Jsn �������� �"�K�F�X�j����� ����ۏ֏���#�� 0�B�k�f�x������� ��ҟ������C�>� P�b���������ӯί������UYSDOEBUG�P�P�)��d�YH�SP_PA�SS�UB?Z�L�OG ��U��S)�#�0�  ���Q)�
MC:�\��6���_MPC ���U���Qñ8�� �Q�SAV ������ǲ%��ηSV;�TEM_TIME 1��[W (�P �Ty��ؿT1SVGUNYS�P�U'�U����ASK_OPTICON�P�U�Q�Q���BCCFG Ì�[u� n�X�G�`a�gZo��߃ߕ��� ��������:�%�^� p�[���������  �����6�!�Z�E�~�@i���������%��� ����&8��nY �}�?��ԫ � �(L:p^ �������/  /6/$/F/l/Z/�/~/ �/�/�/�/�/�/�/2? 8 F?X?v?�?�?? �?�?�?�?�?O*O<O 
O`ONO�OrO�O�O�O �O�O_�O&__J_8_ n_\_~_�_�_�_�_�_ �_o�_ o"o4ojoXo �oD?�o�o�o�o�oxo .TBx�� j������� �,�b�P���t����� Ώ��ޏ��(��L� :�p�^�������ʟ�� o��6�H�Z�؟ ~�l�������د��� ʯ ��D�2�h�V�x� z���¿���Կ
��� .��>�d�Rψ�vϬ� ���Ͼ�������*�� N��f�xߖߨߺ�8� ��������8�J�\� *��n�������� ����"��F�4�j�X� ��|����������� ��0@BT�x �d����� >,Ntb��� ���/�(//8/ :/L/�/p/�/�/�/�/ �/�/�/$??H?6?l? Z?�?~?�?�?�?�?�? O�&O8OVOhOzO�? �O�O�O�O�O�O
__ �O@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<o^o�oro�o�o�o �o�o�o J8 n$O�����X ���4�"�X�B�v���$TBCSG_�GRP 2�B���  ��v� 
 ?�  ������׏����叀��1��U�g�z����~��d, ����?v�	 HC���d�>����e�CL  B���Пܘ���\)>��Y  A�ܟ$�3B�g�B�Bl�i��X�ɼ���X��  �D	J���r�����C ����үܬ���D�@v�=�W�j�}�H�Z� ��ſ����������v�	V3.�00��	m61c�	*X�P�u�Lg�p�>���v�(:��� ��p͟�  O����p������z�JCFG ȖB��� ����������=��=�c�q�K�qߗ߂� �ߦ��������'�� $�]�H��l����� ��������#��G�2� k�V���z��������� �����p*<N ���l����� ��#5GY} h����v�b�� >�// /V/D/z/h/ �/�/�/�/�/�/�/? 
?@?.?d?R?t?v?�? �?�?�?�?O�?*OO :O`ONO�OrO�O�O� �O�O�O_&__J_8_ n_\_�_�_�_�_�_�_ �_�_�_oFo4ojo|o �o�oZo�o�o�o�o�o �oB0fT�x �������,� �P�>�`�b�t����� Ώ�������&�L� �Od�v���2�����ȟ ʟܟ� �6�$�Z�l� ~���N�����دƯ� � �2��B�h�V��� z�����Կ¿���� .��R�@�v�dϚψ� ���Ͼ�������<� *�L�N�`ߖ߄ߺߨ� ���ߚ�������\� J��n������� ���"���2�X�F�|� j��������������� .TBxf� ������ >,bP�t�� ���/�(//8/ :/L/�/�ߚ/�/�/h/ �/�/�/$??H?6?l? Z?�?�?�?�?�?�?�? O�?ODOVOhO"O4O �O�O�O�O�O�O
_�O _@_._d_R_�_v_�_ �_�_�_�_o�_*oo No<oro`o�o�o�o�o �o�o�o&�/>P �/������ ���4�F�X��(� ��|�����֏���� Ə0��@�B�T���x� ����ҟ������,� �P�>�t�b������� ��������:�(� ^�L�n�������2d �����̿�$�Z�H� ~�lϢϐ��������� �� ��0�2�D�zߌ� �߰�j���������� 
�,�.�@�v�d��� �����������<� *�`�N���r������� ������&J\ �t��B��� ���F4j| ��^����/��  2 6# �6&J/6"�$TB�JOP_GRP �2���?  ?�X,i#��p,� �xJ� ��6$�  �<� �� �6$ �@2 �"	 �C��� �&b  C�x�'�!�!>���
5�59>�0+1�33=�CL� �fff?+0?�ffB� J1�%Y?d7�.���/>��2�\)?0�5����;��hCY� ��  @� �!B� � A�P?�?�3EC�  D�!�,�0�*BOߦ?�3JB���
:���Bl�0��0�$�1�?O6!?Aə�AДC�1sD�G6�=q�E�6O0�p��B�Q�;�A�� �ٙ�@L3D	��@�@__�O�O>BÏ\JU�OHH�1ts}�A@33@?1� C�� �@�_�_&_8_>��D�UV_0��LP�Q30<{�zR� @�0�V�P!o3o �_<oRifoPo^o�o�o �oRo�o�o�o�oM (�ol�p~���p4�6&�q5	�V3.00�#m761c�$*(��$�1!6�A� Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,IR�C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^S@;Q��|8�E`rz@/&�8�6&�<��1�w�^$ES�TPARS  �*({ _#HR��AB_LE 1�p+Z�6#|�Q� � 1�|��|�|�5'=!|�	�|�
|�|�˕6!�|�|�|���RDI��z!ʟܟ� ��$���O������ ¯ԯ�����S��x# V���˿ݿ��� %�7�I�[�m�ϑϣ� �����������U-�� ��ĜP�9�K�]�o���-�?�Q�c�u���6�N�UM  �*z!� >  Ȑ�����_CFG ������!@b IMEBF_TT����x#��a�VER��b�w�a�R 1�p+
' (3�6"1 ��  6!����������  �9�$�:�H�Z�l�~� ���������������^$��_��@x�
�b MI_CHAN�m� x� kDBGLV;0o�x�a!n �ETHERAD �?�� �y��$"�\&n ROUmT��!p*!�*�SNMASK��x#�255.�h�fx^$OOL�OFS_DI���[ՠ	ORQCTRL �p+;/�� �/+/=/O/a/s/�/ �/�/�/�/��/�/�/�!?��PE_DET�AI��PON_�SVOFF�33P_MON �H��v�2-9STRTC_HK ����42VTCOMPA�Ta8�24:0FPR�OG %�%�CA)&O�3ISP�LAY��L:_IN�ST_MP GL�7YDUS���?�2L�CK�LPKQUIC�KMEt �O�2SC�RE�@�
tps��2�A�@�I���@_Y���9�	S�R_GRP 1Ҿ� ��� \�l_zZg_�_�_�_�_�_�^�^�oj�Q'O Do/ohoSe��oo�o �o�o�o�o�o! WE{i�������	1234�567��!���X��E1�V[
 �}�ipnl/a�g?en.htmno���������ȏ~�P�anel setup̌}�?��0�B�T�f� ��񏞟 ��ԟ���o���� @�R�d�v������#� Я�����*���ϯ ůr���������̿C� �g��&�8�J�\�n� ����϶��������� uϣϙ�F�X�j�|ߎ� �����;��������0�B��*NUALR�Mb@G ?�� [���������� �� ��%�C�I�z�m�������v�SEV � ����t�E?CFG Ձ=]�/BaA$   B�/D
 ��/C� Wi{�����@�� PRց;C �To\o�I�6?K0(%����0 �����//;/ &/L/q/\/�/�/�/lƇD �Q�/I_��@HIST 1׾�9  ( � ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1?v?�?�?ά?�� >?P=962c?�?
OO.O�?�?�136�?|O�O�O�O AOSOeO�O__0_�H M___q_�_�_�_�_H_ �_�_oo%o7o�_[o moo�o�o�oDo�o�o@�o!3E ��a 81�ou����� �o���)�;�M�� q���������ˏZ�l� ��%�7�I�[��� ������ǟٟh���� !�3�E�W�������� ��ïկ�v���/� A�S�e�Pb������ ѿ������+�=�O� a�s�ϗϩϻ����� ��ߒ�'�9�K�]�o� ��ߥ߷��������� ��#�5�G�Y�k�}�� ������������� 1�C�U�g�y���v��� ��������	�? Qcu��(�� ��)�M_ q���6��� //%/�I/[/m// �/�/�/D/�/�/�/? !?3?�/W?i?{?�?�? �?�����?�?OO/O AOD?eOwO�O�O�O�O NO`O�O__+_=_O_ �Os_�_�_�_�_�_\_ �_oo'o9oKo�_�_ �o�o�o�o�o�ojo�o #5GY�o}������?��$�UI_PANED�ATA 1������  	�}�0�B�0T�f�x��� )���� mt�ۏ����#�5� ��Y�@�}���v����� ן�������1��U�pg�N������ �1��Ïȯگ���� "�u�F���X�|����� ��Ŀֿ=������ 0�T�;�x�_ϜϮϕπ�Ϲ������,ߟ� M��j�o߁ߓߥ߷� �����`��#�5�G� Y�k��ߏ������ ��������C�*�g� y�`���������F�X� 	-?Qc��� �߫���� ~;"_F��| �����/�7/ I/0/m/�����/�/�/ �/�/�/P/!?3?�W? i?{?�?�?�??�?�? �?O�?/OOSOeOLO �OpO�O�O�O�O�O_ z/�/J?O_a_s_�_�_ �_�O�_@?�_oo'o 9oKo�_oo�oho�o�o �o�o�o�o�o#
G Y@}d��&_8_ ����1�C��g� �_��������ӏ��� ^���?�&�c�u�\� ������ϟ���ڟ� )��M��������� ��˯ݯ0�����7� I�[�m���������� ٿ�ҿ���3�E�,� i�Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#��� ���� ��$�6��Z� A�~�e�w������ �����2��V�h�O������v�p��$UI�_PANELIN�K 1�v��  � � ��}1234?567890���� 	-?G ���o �����a��@#5G�	����4p&���  R� ����Z��$/ 6/H/Z/l/~//�/�/ �/�/�/�/�/
?2?D? V?h?z??$?�?�?�? �?�?
O�?.O@OROdO vO�O O�O�O�O�O�O _�O�O<_N_`_r_�_�_�0,���_�X�_ �_�_ o2ooVohoKo �ooo�o�o�o�o�o�o ��,>r}��� �������� �/�A�S�e�w���� ����я���tv�z� ���=�O�a�s��� ����0S��ӟ���	� �-���Q�c�u����� ��:�ϯ����)� ��M�_�q��������� H�ݿ���%�7�ƿ [�m�ϑϣϵ�D��� �����!�3�Eߴ_i� {�
�߂����߸��� ���/��S�e�H�� ��~��R~'�'�a� �:�L�^�p������� �������� ��6 HZl~���#� 5��� 2D�� hz�����c �
//./@/R/�v/ �/�/�/�/�/_/�/? ?*?<?N?`?�/�?�? �?�?�?�?m?OO&O 8OJO\O�?�O�O�O�O �O�O�O[�_��4_F_ )_j_|___�_�_�_�_ �_�_o�_0ooTofo ��o��o��o�o�o ,>1bt� ���K���� (�:����{O���� ��ʏ܏�uO�$�6� H�Z�l���������Ɵ ؟����� �2�D�V� h�z�	�����¯ԯ� �����.�@�R�d�v� �������п���� ��*�<�N�`�rτ��O �Ϻ�Io��������� 8�J�-�n߀�cߤ߇� ���߽����o1�o X��o|�������� �����0�B�T�f� �������������S� e�w�,>Pbt� �'���� �:L^p��# ���� //$/� H/Z/l/~/�/�/1/�/ �/�/�/? ?�/D?V? h?z?�?�?�???�?�? �?
OO.O��ROdO�� �OkO�O�O�O�O�O�O _�O<_N_1_r_�_g_��_7OM�m�$�UI_QUICK�MEN  ���_AobR�ESTORE 1��  �|��Rto�o�im�o�o�o�o �o:L^p�%� �����o��� �Z�l�~�����E�Ə ؏���� �ÏD�V� h�z���7�������/� ��
��.�@��d�v� ������O�Я���� �ßͯ7�I���m��� ����̿޿����&� 8�J��nπϒϤ϶� a�������Y�"�4�F� X�j�ߎߠ߲����� �ߋ���0�B�T�goSCRE`?#mu1sco`Wu2��3��4��U5��6��7��8��bUSERq�v��Tp���ks����4���5��6��7��8���`NDO_CFoG �#k  n`� `PDATE� ���N�onebSEUFRAME  �T�A�n�RTOL_�ABRTy�l��E�NB����GRP �1�ci/aCz  A�����Q�� $6HRd���`U�����MSKG  �����Nv�%�U�%���b�VISCAND_wMAX�I���FAIL_IM)G� �PݗP#���IMREGNUMr�
,[SIZ��n`�A�,VO�NTMOU���@���2��a���a�����FR:\ �� MC:\ޚ\LOG�B@F� !�'/!+/�O/�Uz M�CV�8#UD1&r&EX{+�S�P�PO64_��0n'fn6PO��CLIb�*�#V����,f@�'�/� �=	�(SZV�.�;���'WAI�/STAT ���B�P@/�?�?�:$�?��?��2DWP  ��P G@+b=��� H�O�_JMPERRw 1�#k
  ��2345678901dF�ψO{O�O�O �O�O�O_�O*__N_�A_S_�_
� MLO�Wc>
 �_TI�=�'MPH?ASE  ��F���PSHIFT֗1 9�]@< �\�Do�U#oIo�oYo ko�o�o�o�o�o�o�o 6lCU�y ����� ��	��V�-�e2����	�VSFT1�2	uVM�� �5�1�G� ���%A� W B8̀̀�@ pكӁ˂�у��z�#ME@�?�{��!�c>&%�aM1��k�0�{ �$`0T?DINEND���\�O� �z����Sp��w��P���ϜRELE�Q��Y����\�_ACTIV���:�R�A �`�e���e�:�RD� ����YBOX ��9�د�6��02����190�.0.�83���254��QF�	 �X�j��1��robo�t���   �p�૿�5pc��̿�����7���x��-�f�ZABC�����,]@U��2ʿ� eϢωϛϭϿ�����  ���V�=�z�a�s�$��E�Z��1�Ѧ