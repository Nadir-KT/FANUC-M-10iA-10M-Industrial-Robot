��   I�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���B�IN_CFG_T�   X 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �ET�H_FLTR.�� $�  � �FTP_C�TRL. @ ?$LOG_8	��CMO>$DN�LD_FILTE�� � SUBDIR�CAP�j� HOv��NT. 4� �H_NAME �!ADDRT�YPA H_LE�NGTH' ��z +LS �D $ROBO�TIG PEER�^� MASKM�RU~OMGDEuV#� RDM*��DISABL�&� TCPI�G/ 3 $AR�PSIZ&_I{PF'W_MC�ދF_IN� FA�~LASSs�H{O_� INFO���TELK P�V�b	 WO�RD  $A�CCESS_LV�L?TIMEOU=TuORT � ��ICEUS= ���$#  �����!�� � � VIRTUAL�/�!'|0 �%
���F�����$�%����+ ������$�� �-2�%;�SHARED� 1�)  CP!�!�?���!|? �?�?�?�?O�?%O�? 1OOZOOBO�OfO�O �O�O�O_�O�OE__ i_,_�_P_�_t_�_�_ �_o�_/o�_SooLo �oxo�opo�o�o�o�o �o*Os6� Z�~����� 9��]� ���D�V��� z�ۏ����#����Y�H�}�@���)7z _LIST 1=_x!1.ܒ0���d�ە1�d�25c5.$������%ړ2��X���+�=�O�3Y��Р�������O�4ѯ�H���	��-�O�5I���� o�������O�6����8������ �$ ���-� ���-� ��&�%��&!Ò�)��0H!� ����rj3_tpd����! � �!!KC� e�0ٙ��&W�!Cm ��w߉�~S�!CON� ���1�=�smon��W�