��   D�A��*SYST�EM*��V7.5�0122 8/�1/2   A �
  ���C�ELLSET_T�   w$�GI_STYSEL_P 7_T  7ISAO:iRibDi�TRA�R��I_INI; ���t�bU9ARTaRSRPNS1Q�2345*678Q
�TROBQACKSNO��) �7�E�S�a@�o�z2 U3 4 5 6 �7 8awn&GINm'D�&��)%� �)4%��)P%��)l%3SN�{(OU��!|7� OPTNA�73�73.:B<;}a6�.:C<;CK;CaI?_DECSNA�38R�3�TRY1���4��4�PTHC�N�8D�D�INCYC@HG�KD�?TASKOK�{D �{D�7:�E�U:�C h6�E�J�6�C�6U�J��6O�;0U��:IAT�L0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T��T�@REQ�d��drG�:Mf�GJO_HFAUL�Xd�dvgALE� �g�c�g�cvgE� �H�dvg�NDBR�H�dgR�GAB�Xtb   �CLMLIy@�   $�TYPESIND�EXS�$$CL�ASS  �S��lq����apVIRTUALi�{q'61ION  �����q�t+ UP0 �u�q�Style� Select �	 ;p��r�uRe�q. /Echo:���yAck����sInitiaQt�p�r�s�t@�$O�a�p���	�� � ������
�����q��������q��sOption bit A���B����C�D�ecis�cod�;��zTryout� mL��Path� segJ�ntikn.�II�yc:���Task OK���!�Manual� opt.r�pA�ԖBޟԖC�� ?decsn ِ��Robot interlo�"�>�� isol3��C⚒i/�"�z�ment��z�ِ����_��status�	�MH Faulty:��ߧAler�p�%��p@r 1�z L��[�m�+�; �LE_COMNT� ?�y�   ��䆳�Ŀֿ��� ��0�B�T�g�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ߀�������������Up������   ��ENAB  ���u�������<�ꐵMENU>�y���NAME ?%��(%$*4���D� ;p2�k�V���z����� ��������1U @Rdv���� ���*<u `������� �/;/&/_/J/f/n/ �/�/�/�/�/?�/%? ?"?4?F?X?j?�?�? �?�?�?�?�?�=