��   38�A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���U�I_CONFIG�_T  T �($NUM_MENUS  9�* NECTCRE�COVER>CCOLOR_CRR�:EXTSTAT���$DUMMY�36CMEM_L�IMIR$DB�GLVL�POPUP_MASK��zA  �7��ODE�
8CF�OCA �9CP�S)C��g 
H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � �NU_FAVB ?� 
$HLP> 7_DIQ?� m�ELEMV}URȥ h� So�$7HMI�RO'X�W ADONLY�� �TOUCH�PROOMM�O?$�ALA�R< �FILVE9W�ENB=�!%bC -"USE�R6)FCTN6)W�I�� I* _E�D�h"R!_TIT�L�  &US�TOM0 t �$} RT_SP�ID��$C�$*P�AG� ?ZDE�VICE�)SCR�EqEF���'N~�@$FLAG��@�"USRVI| 1  < \ +2�,1PR-I�m� A� K0�TRIP�"m�$�$CLASS  ����l1��Rz��Ra0VIRTO1�j?|0'2 )�E��)�O`R�	 �%,��;����2�0��3�3�1�� ,� �  <�?��
 ��s1,O@>OPObOtO�O�O (O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ ���@���� �/��S�e�w����� ��<�я�����+��=� TPT�X��͈`�r� � sH���$/s�oftpart/�genlink?�help=/md�/tpmenu.dg?�ٟ����ȏ 3�E�W�i�{������ ïկ�������A� S�e�w�����*���ѿ`�������9����F�6�3C�($ ��p���^ϗςϻ���s1�1���?K�����q�̛3�" 1�5ޱ2 \�6 �REC VE�D��U�g�who�lemod.ht}m{�singl���doub���trip��brows�߯�h�
� �.���R�d�v������R�<�v߈�dev�.s��l���(�1�	t?���(����� ������|�������G� �0_q ������� @[0Bf x��I�B<�� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ?��??B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�OT �O�O�O�O	__-_?_ Q_c_^�_�_h_z_�_ �_���O)o$o6oHo qolo~o�o�o�o�o�o �o IDV$? vp������ 
��.�@�R�d�v��� ������Џ⏰O�/� A�S�e�w��������� �_���ğ֟+�=��_ o쏅�������ͯȯ گ���"�4�]�X� j�|��������ҿ̿ ����0�B�T�f�x� �ϜϮ���������� �,�>��yߋߝ߯� ��������	���?� Q� �2���P�b�H� ������ �)�$�6�H� q�l�~����������� ��ܿ.(Vh z������� 
.@Rdv� �h����//// A/S/e/w/r�/�/|/��/�/�/:�$UI�_USERVIE�W 1��R 
���6?H?�mg?�?�? �?�?�?{?�?O O2O DO�?hOzO�O�O�O[? �O�O�OSO_._@_R_ d__�_�_�_�_�_�_ �_oo*o<oNo�O[o moo�_�o�o�o�o �o&8J\n� �����o��� }/�X�j�|�����C� ď֏������0�B� T�f�x�#�������� �����,�ϟP�b� t�������M�ί�� ����#�5�G����� ������ʿm�� �� $�6�ٿZ�l�~ϐϢ� M�W�����E��� �2� D�V�h�ߌߞ߰��� ��w���
��.�@��� M�_�q��߬������ ����*�<�N�`�r� ��������������� ����J\n�� 5������" 4FXj�� ���//0/� T/f/x/�/�/?/�/�/ �/�/?�(