��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 W �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$� � NO�P�S_SPI_IN[DE��$�X��SCREEN_NAME �/SIGN��~� PK_FIL�	$THKYMP�ANE�  	�$DUMMY �� u3|4|GR�G_STR1 � $TITP_$I��1�@{�����5�U6�7�8�9�0��z������1�1�1 '1�
'2"GSBN_�CFG1  8� $CNV_J�NT_* |$D�ATA_CMNT��!$FLAGS|�*CHECK�!��AT_CELL�SETUP � P $HOM�E_IO,G�%��#MACRO�"R�EPR�(-DRU�N� D|3SM�5H UTOBAC�KU0 � �$ENAB��!E�VIC�TIk � D� DX!2�ST� ?0B�#$INTERVAL!2�DISP_UNI�T!20_DOn6E{RR�9FR_F�!2IN,GRES��!0Q_;3!4C�_WA�471�8GW�+0�$Y $DB\� 6COMW!2�MO� H.	 �\rVE�1$F8�RA{$O�UD�cB]CTMP1_FtE2}G1_�3�B�2�FXD�#
 �d $CARD�_EXIST4�$FSSB_TY�P!AHKBD_YSNB�1AGN Gn� $SLOT�_NUM�APR{EV4DEBU� �g1%�;1_ED�IT1 � *1G=� S�0�%$EP�$�OP�U0LE�TE_OK�BUSބP_CR�A$�;4AV� 0LACIw1�R�@k �1$@�MEN�@$D �V�Q`PvVA{G �BL� OU&R A,A�0�!� B� OLM_O�
eR�"�CAM_;1 �xr$ATTqR4�@� ANNN@�5IMG_HEI�GH�AXcWIDTMH4VT� �UU0F_ASPEC�Aw$M�0EXP�v.@AX�f�CF�D� X $GR�� � S�!.@B�PN�FLI�`�d� UI�RE 3T!GITC�H+C�`N� S�d_�LZ`AC�"�`EDTp�dL� J�4S�0@� <za�!p;G0� � 
$WARNM�0f�!�@� �-s�pNST� CO�RN�"a1FLTR^{uTRAT� T}p�  $ACC�a1�p��|{�rOR�I�P�C�kRT0_YS~B\qHG,I1 [ T�`�"3I�pTYD�@*2 3`#@� �!�B*�HDDcJ* Cd�2�_�3_�4_�5_�6*_�7_�8_�94�0w�CO�$ <� ��o�o�hK3 1#`O_�Mc@AC t 2� E#6NGPvABA� �c1�Q8��`,��@nr1�� d��P�0e�]p� cvnpUP&Pb26���p��"J�p_R�rPBCb��J�rĘߜJV�@ U� B��s}�g1�"Yt�P_*0OFS&R; @� RO_K8T��aIT�3T�NOM	_�0�1p�3� >��D �� Ќ@��hPV��mEX�p� �0�g0ۤ�p�r
$TyF�2C$MD3i��TO�3�0U� F� ���Hw2tC1(�Ez�g0#E{"F0�"F�40CP@�a�2 �@$�PPU8�3N)ύR&ևAX�!DU��;AI�3BUF�F=�@1 |pp���pkPIT� PP�EM�M�y��F�SIMQSI�"ܢ�VAڤT��@�w 	T�`(zM��P�B�q�FACTb�@E�W�P1�BTv?�M]C� �$*1�JB`p�*1DEC���F��ňP���� �H0CHNS�_EMP1�$G��8��@_4�3�p|@P��3�TCc�(r/� 0-sx��ܐ� MBi���!����JR� i�S/EGFR��Iv �a�R�TpN�C��P�VF4>�bx &��f{uJc!�Ja ��� !28�ץ�AJ����SIZ�3S�c�B�T�M���g��JaRSINFȑb���q�۽��н����L�3�B����CRC�e�3CC p����c��mcҞb��1J�cѿ�.����D
$ICb�Cq�5r�ե�0�@v�'���EV���zUF��_��F,pN��
ܫ�?�4�0A�! �r���h�Ϩ� �p�2�͕a�� �د��A	�Cx �Ϗ��o"27�!ARtV�O`C�$LG�pV�B�1�P��@�t�a!A�0'�|�+0Ro�� MEp`"1 C3RA 3 AZV�g46p�O �FCCb�`��`F�`K������ADI��a�A�bA�'�.p��p�`�c�`S04PƑ�a�AMP��-`IY�3P�M�]pUR���QUA1  $@TITO1/S@S�!�����"0�DBPXW�O��B0!5�$SK���C�x q�!�"�"�PR�� �
� =����!# l@q1$2�$z�
��L�)$�/���� )%�/�$C�!&?�$gENE�q.'*?��Ú RE�p2(�H ��O�0#$L|3$$�#�B[h�;���FO_D��ROSr�#�������3RIGGER��6PApS����ET�URN�2�cMR_�8�TUw��0EkWM��M�GN�P����BLAH�<E��<�P��&$P� �'P@�Q3�CkD{���DQ���4�11��FG�O_AWAY�BM�O�ѱQ#!�D�CS_�)  �PIS� I gb {s �C��A��[ �B$�@S��AbP�@�EW-�NTNTVճ�BV�Q�[C�(c`�UWr�P�J���P�$0��SAFE܇��V_SV�bEX�CLU��nONL2��SY�*a&��OT�a'�HI_V��4��B���_ �*P0� 9�_z��p� �TSG�� +nrr�@6Acc*b��G�#@E�V.iHb?fANNUN$0.$fdKID�U�2�SC@��`�i�a��j�f���z��@I$2,O�$1FibW$}�OT9@�1� $DUMMAYT��da��dn�f0|� �E- ` ͑HE4(sg�*b�SAB���SUFFIW���@CA=�c5r�g6�abMSW�E�. 8Q�KEYI5���TM�10s�qAF�vIN��#�p�D��/ D��HOST_P!�rT��ta�`�tn��tsp�pEMӰ�V�����pLc UL>I�0  8	=�ȳ��f0Tk0�!1 ϴ $S��ESAMPL��j�۰f璱�f���I�0��[ $SUB�k�#0�C��8T�r#a�SAVʅ���c���C��P�fP�$n0E�w YN_�B#2 0Q�DI�{dlpO(��9#$��R_I�� �?ENC2_S� �3  5�C߰��f�- �SpU����!4��"g�޲�1T���5X�j`ȷg��0�0�K�4�AaŔAVE�R�qĕ9g�DSP�v��PC��r"��x(���ƓVALUߗ�HE�ԕM+�IP\ճ��OPP ��CTH��֤��P�S�$ �۰F��df�J�l �qRS�ET+�6 H�bLL_DUs�~a3@{��3:���OTX"���s�a�0NOAUT5O�!7�p$)�$�*��c4�(�C� �8�C, �p�&�L��� 8H *8�LH <6����c"� �`, `Ĭ�kª�q��@q��sq��~q��7���8��9��0����1���1̺1ٺ1�1��1 �1�1�2R(�2����2̺2ٺU2�2�2 �2�U2�3(�3��3���̺3ٺ3�3�3� �3�3�4(�%���?��!9 A<�9�&�z��I��01���M��QFE@'@΂ : ,6��Q?3 �@P?9��
5�9�E�@A�a�A�� ;p$TP~�$VARI:��ʠ��@P2�P< ���TDe���K`�Q���OP��BAC�"= T�p��e$�)_,�bn�kp+ IF�IG�kp�H  ��Pİ!�F@`�!>Gt ;E��sC�ST�D� D���c�<� 	C��{�� _���l���R  ���FORCEUP?b^��FLUS�`H��N>�F ���RD_CM�@E������ ��@vMP��REMr F �Q��1k@���7Q
�K4	NJ�5EFF�ۓ:�@IN2Q��O�VO�OVA�	TgROV���DTՀ�DTMX� � �@�
ے_PH"p��CL��_TpE�@d�pK	_(�Y_T��Tv(��@A;QD� ������!0tܑ&0RQ���_�a��2��M�7�CL�dρ�RIV'�{��EAmRۑIOHPC�@d����B�B��CM9@����R �GCLF�e!DYk(M�a6p#5TuDG��8� �%�qFSSD �s�? P�a�!�1����P_�!�(�!1��E��3�!3�+5�&�GSRA��7�@��;ᚔPW��ONn��EBUG_SD2H�P�{�_E A ��p�=��TERM�`5Bi5��O�RI#e0Ci5�p�GSM_�P��e0Di5����TA�9E��9UP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1젎4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ3Q�E�p %B`�'EC����@R$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"��A��?���ERV��XQ�Y�� mG>@�BN��U\���R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`� 0SMT6�G�3�GR��13�aPA�L@��p�q�uH �� ���TOC$A�`P	P�`������p�ѡ�`0O,��RE�`R4C�A�O�p낎Be�`R��Eu�h�A��e$P�WR�IMu�RR�_�cN��q=B I�&2H���p_ADD�R��H_LENG��B�q�q�q$�R��S��JڢSS��SK�N��u\��u̳�uٳS�E�A�jrS��MN�!K�����b����OLX��p�<���`ACRO3pJ� �@��X�+��Q��6�OUP3�b_�IX��a�a1��}򚃳� ��(��H��D��ٰ���氋�IO2S��D�����	�7��L $d��`Y!_O�FFr��PRM_���b��HTTPu_+�H:�M (|p�OBJ]"�p��$���LE~Cd���N� � ��֑AB%_�TqᶔS�`6H�LVh�KR"u�HITCOU��B-G�LO�q����h�����`��`SS� ���HW�#A:��Oڠ<`INCP}U2VISIOW� ͑��n��to��to�ٲ� �IOLN��P� 8��R��r�$�SLob PUTM_n�$p��P& x¢��Y F_AS�"Q��$L������DQ  U�0	P4A��^���ZPHY��-���y��UOI �#R `�K����$�u�"pPpk����$�����Y�UJ5�S�-���NE6WJOG�KG̲DIS���K�p���#T (�uAV8F�+`�CTR�C
��FLAG2��LG�dU ���؜�13?LG_SIZ����`b�4�a��a�FDl�I`�w� m�_�{0a� ^��cg���4�����������{0��� SCH�_���a7�N�9�V
W���E�"����4�"�UM�Aљ`LJ�@�7DAUf�EAU�p��d|�r�GH�ba����BOO��WL ?�6 IT��y0��REC��SCR� ܓ�D
�\���MARGm�!��զ ���d%�����S����Wp���U� �JGM[��MNCHJ���FN�KEY\�K��PR�G��UF��7P��F�WD��HL��STP��V��=@��А�RS��HO`����C�9T��b ��7�[�U L���6�(RD� ����Gt��@PO������z��MD�FOCU���RGEX��TUI��I��4�@� L�����P����`���P��NE��CAN�A��Bj�VAIL�I�CL !�UDCS�_HII4��s�O��(!�S���Sܿ�%��_BWUFF�!X�?PTH$m���v`��ķ���AtrY��?P��j�3��`OS1
Z2Z3Z8��`Z � ��[aE�Ȥ��ȤIDX�dP�SRrO���zA�S�T]�R}�Y&�� _Y$E�C����K�&&���ѿ![ LQ��+00�	P�� �`#qdt
�U�dw<���?_ \ �`4Р��\��Ѩ#\0C4�]{ ��CLDP]�>�UTRQLI��d8ڰ�)�$FLG&�� �1�#�D���'B�LqD�%�$�%ORGڰ 5�2�PVŇVY8�s�T8�r�$}d^ ���$(6��$�%S�`T� ��B0�4�6RCLM�C�4]?o?�9세�M9I�p}d_ d=њ�RQ��DSTB�p� ;F�HH�AX�R JHdLE�XCESr��BM!p�a`��/B�T�F���`a�p=F_A@7Ji��KbOtH� K�d�b \Q���v$M�BC�LI|�)SREQUIR�R�a.\o��AXDEBUZ�AL
t M��c�b�{P��8��2D�MNDRѧ`®`d;�2�ȺSDC��N�INl�K�x`찄�X� N&��aZ���EL�SPST� �ezrLOC�RYIrp�EX<fA�px�9AAODAQ��7f XY�OND��"MF,Łf�s"��`}%�e/� ���FX3@�IGG�� g ��t"��ܓs#N�s$R�a%��i]��h�]�v�@�DATA#?pE�%�tR��Y��Nh t $+MD`qI}�)nv� ytq�ytHP`�Pxu��<(�zsANSW)�yt(@��yuD+�)\b��ܵ0o�i �@CU�w�V�p 0XeRR2��j Du�{Q��7B?d$CALIA@���G��2��RIN���"�<6�INTE��Ck�r^�آXb]���_N�qlk���9��D���Bm��DIVFFDH�@���qnI�$V,��S�$��$Z�X�o��*����oH ?�$BELT�u!_ACCEL�.�~�=�IRC�� ����D�T�8�$PS�@�"L1 �r��#�^�S�Eы T�PAT!H3���I���3x�p�A_W��ڐ���2n�C��4�_MG��$DD��T���$FW�Rp9��I�4���DE7�PPAB�N��ROTSPE!E�[g�� J��[��C@4�1 $US�E_+�VPi��S�YY���1 �aYNr!@A�ǦOFF�qnǡMOU��NG����OL����INC �tMa6��HB��0HBENCS+�8q9Bp�X4�FDm�IN�Ix�0]��B��VE��#�>y�23_UP񕋳/LOWL���p� B���Du�9B#P`��x ���BCv�r�MO3SI��BMOU��@��7PERCH  ȳOV��â
ǝ� ���D�ScF�@MP����� Vݡ�@y�j��LUk��Gj�p�UPp=ó���ĶTRK�>�AYLOA�Qe� �A��x�����N`�F��RTI�A$��MO UІ�HB�BS0�p7D5����ë�Z�DU�M2ԓS_BCKLSH_Cx�k�� ��ϣ���=���ޡ< �	ACLAL"q�p�1м@��CHK� :�S�RTY���^�%E1Qq_�޴_�UM�@�C#��S�CL0�r�LMT_OJ1_L��9@H��qU�EO�p�b�_�e�k�e�SPC��u�L��N�PC�N�Hz �\P��C�0~"XT\��CN_:�N9�L�I�SF!�?�V����U�/���x�T���CB!�SH�:��E� E1T�T����y���T�f�PA ��_P��_� =������!����J6 L�@���OG�G�TORQU��ONֹ��E�R0��H�E�g_W2��ā_郅���I*�I�I��Ff`xaJ�1�~1�VC3�0BD:B�1�@SBJRKF9~�0DBL_SM�:�2M�P_DL2GRV�����fH_��d���CcOS���LNH ��������!*,�aZ���fcMY�_(�TH���)THET0��N�K23���"��C-B�&CB�CAA�B��"��!��!�&SB8� 2�%GTS�Ar�CIMa�����,4#<97#$DU���H�\1� �:Bk62�:AQ�(rSf$NE�D�`I ��B+5��$̀�!�A�%�5�7���LCPH�E�2���2S C%C%�2-&FC0JM&̀V�8V�8߀LUVJV!KV/KV=KUVKKVYKVgIH�8@FRM��#X!KH/KUH=KHKKHYKHgI�O�<O�8O�YNO�JO!KO/KO=KO*KKOYKOM&F�2�!�+i%0d�7SPBA?LANCE_o![c�LE0H_�%SP�c� &�b&�b&PFULC�h�b�g�b%�p�1k%�UTO_<��T1T2�i/�2N��"�{�t#�Ѡ�`�0�*�.�T��O�À<�v INSEG"�ͱREV4vͰl�gDIF�ŕ�1lzw6��1m�0OBpq�ь�?�MI{���nL�CHWARY���A�B��!�$MEC�H�!o ��q�AX���P����7Ђ�`n� 
�d(�U�RO�B��CRr�H���N��SK_f`�p� P �`_��R /�k�z�����1S�~��|�z�{���z��qIN�Uq�MTCOM�_C� �q  ����pO�$NO�REn����pЂ7r 8p GRe�u�SD�0AB�$?XYZ_DA�1a���DEBUUq�������s z`$��COD�� L���p��$BUFIwNDX|�  <��MORm�t $فUA��֐����y��rG��u �� $SIMUL�  S�*�Y�̑a�OB�JE�`̖ADJUyS�ݐAY_I�S�D�3����_F-I�=��Tu 7� ~�6�'��p} =�C�}pt�@b�D��FRIrӚ�T��RO@ \�E�}'�8c�OPWO�Yq�v0Y�SY�SBU/@v�$SO!Pġd���ϪUΫ}p�PRUN����PA�D���rɡL�_O�Uo顢q�$^)�IMAG��w���0P_qIM��L�I�Nv�K�RGOVCRDt��X�(�P*�J�|��0L_�`]�L�0�RB1�0��M��ED}��p ʚ�N�PMֲ��u%��w�SL�`q�w� x $OVS�L4vSDI��DEX����#���-�	V} *�N4�\#�B�P2�G�B�_�M����q�E� x Hxw��p��ATUSWЅ��C�0o�s���BSTM�ǌ�I�k��4��x�԰q�y DBw�E&���@E�r���7��жЗ�EXE ��ἱ�����f q�gz @w���UP'�f�$�pQ�XN����������� �P�G΅{ h $GSUB����0_��|�!�MPWAIv�P7ã�LOR�٠F�\p˕$RCVF�AIL_C��٠B�WD΁�v�DEF�SP!p | L�w���Я�\���UCNI+�����H�R�,p}_L\pP��x�t���p�}H�> �*��j�(�s`~�N�`KE)TB�%�J�PE Ѓ�~��J0SIZE�����X�'���S�O�R��FORMAT��`��c ��WrEM2�t��%�UX��G���PLI��p� � $ˀP_S�WI�pq�J_PL~��AL_ ���J��A��B��� C���D�$E���.�C_�U�� � � ���*��J3K0����TIA�4��5��6��MOM��������ˀB��AD��������6��PU� NR��������m��?� A$PI�6q� �	�����K4��)6�U��w`��SPEEDgPG���� ����Ի�4T�� �� @��SAM�r`��\�]��MOV_�_$�npt5��5$���1���2���� ����'�S�Hp�IN�'�@�+�����4($4+T+GA�MMWf�1'�$G#ET`�p���Da���=

pLIBR>�I]I2�$HI=�_g�Ht��2�&E;��(A�.� �&LW�-6<�)@56�&]��v�p��V���$PDCK����q��_?���� �q�&���7��4����9+� �$I/M_SR�pD�s�r�F��r�rLE���O0m0H]��0�6c��ܬpq��PJqUR_SCRN�FA����S_SAVE_DX��dE@�NOa�CA A�b�d@�$q�Z�Iǡ s	�I� �J�K� ��� �H�L��>�"hq� �����ɢ�� �bW^US�A�-M4���a��)q`��3��WW�I@v�_�q�.M�UAo�� � $sPY+�$W�P�vNG�{��P:��R`A��RH��RO�PL��@���q� ��s'�X;�	OI�&�Zxe ���m�G� p��ˀ�3s��O�O�O�O�O�aa�_т� |��q�d@�� .v��.v��d@��[wFv���E���%s�t;B��w�|�tP���P�MA�QUa ���Q8��1٠QTH��HOLG�QHY�S��ES��qUE��pZB��Oτ�  ـPܐ(�A����v�J!�t�O`�q��u��"���FA��IROG�����Q2���o�"�x�p��INFOҁ��׃V����R���O�I��� (�0SLEQ������Y�3�H���Á��P0Ow0Ԟ��!E0NU���AUT�A�COPY�=�/�'��@Mg�N��=�}1������� ��RG��Á�f��X_�P�$;�(���`��W��P��@������EXT_CYC bHᝡRprÁ�r��_NAec!А���ROv`~	�� � ���POR_�1�E2��SRV �)_�I�DI��T_�k�}�'����dЇ�����5��6J��7��8i�2ASdBZ���2�$��F�p���GPLeAdA
�TAR�Б@���P���裔d� ,��0FL`�o@YN���K�M��Ck��P�WR+�9ᘐ��D�ELA}�dY�pA�D�a�RQSKIPN4� �A�$�OB`�NT����P_ $�M�ƷF@\bIpݷ� ݷ�ݷd����빸���Š�Ҡ�ߠ�9���J2R� ���� 4V�EX� TQ Q����TQ������ ���`�#�RDC�V�S �`��X)�R�p������r��m$RGoEAR_� IOBT��2FLG��fipE	R�DTC���Ԍ��ӟ2TH2NS}� �1���G TN\0 ���u�M\��`I�dG�REF:�1Á� l�h���ENAB��cTPE�04�]����Y�]� �ъQn#��*��"�������2�Қ�߼��߸����� ��3�қ'�9�K�]�o��
�4�Ҝ�������(�����5�ҝ!�3��E�W�i�{��6�Ҟ��������������7�ҟ-?Qcu
�8�Ҡ����x���SMSKÁ%�l��a��EkA��oMOTE6������@�݂TQ�IO�}5�ISTP��PO9W@��� �pJ� ���p����E�"�$DSB_SIG!N�1UQ�x�C\��/S232���R�i�DEVICEUS��XRSRPARIT|��4!OPBIT�Q�I�OWCONT�R+�TQ��?SRCU�� MpSUXTAS�K�3N�p�0p$TATU�PE#�0������p_XPC)��$FREEFRO�MS	pna�GET\�0��UPD�A�2ΙqRSP� :���� !$US�AN�na&����ER1I�0_�RpRYq5*"�_j@_�Pm1�!�6WRK9KD���6��~QFRIEND�Q��RUFg�҃�0TO�OL�6MY�t$�LENGTH_VT\�FIR�pC�@�ˀE> +IUFINt-RM��RGI�1�ÐAITI�$GX�ñ3IvFG2v7G1`���p3�B�GPR�p�1F�O_n 0��!�RE��p�53҅U�T�C��3A�A�F �G((��":���e1n! ��J�8�%���%]���%�� 74�X TO0�L��T�3H&���8���%b453GE�W$�0�WsR�TD�����T��M����Q�T]�=$V 2����1��а91�8�02�;2
k3�;3�:ifa�9�-i�aQ��NS��ZR$)V��2BVwEV�	V�B;�����&�S��`��F�"�k�@�2a�P5S�E��$r1C���_$Aܠ6wP!R��7vMU�cS�t 8'�/89�� 0G�aV"`��p�d`���50��@��-�
25S�� ��aRW����iB�&�N�AX�!��A:@LAh��rTHIC�1I���X��d1TFEj��q�uIOF_CH�3�qI܇7�Q�pG1RxV����]��:�u�_JF�~�PRԀƱ�RV{AT��� ��`0���0RҦ�DOfE���COUԱ��AXI|���OFFSE׆TRIGNS���c�� ��h�����H�Y��IGMA0PA�p�J�E�ORG_U�NEV�J� �S������d �$�CА�J�GROU�����TOށ�!��D;SP��JOGӐ�#&��_Pӱ�"O�q�����@�&KEP�I�R��ܔ�@M}R��A	P�Q^�Eh0��K��SYS�q"K�PG2�BRK�B��߄��pY�=�d����`A�D_�����BSOC����N��DUMMgY14�p@SV�P�DE_OP�#SFSPD_OVR-����C��ˢΓOR$٧3N]0ڦF�ڦ6��OV��SF��p���F+�r!���CC�|�1q"LCHDL��RECOVʤc0���Wq@M������ROȮ#��Ȑ_+��� �@0�e@VER�o$OFSe@CV/ �2WD�}��Z2,���TR�!����E_FDO�MB�_CM���B��BAL�bܒ#��adtVQ R�$0p���G$�7�AM5��� eŤ�σ_M;��"'����8�$CA��'�E�8�8�$HBK(1���I�O<�����QPPA������
��Ŋ��~��DVC_DBhC�;��#"<Ѝ�r!S�1�[ڤ�S�3[֪�AT�IOq 1q� ʡU8�3���CABŐ�2��CvP��9P^�B���_�� �SUBCPU�ƐS�P �M�)0�NS�cM�"r�$HW_C��U��S@���SA�A�pl$UNkITm�l_�AT��x�e�ƐCYCLq��NECA���FLTR_2_FIO�07(��)&B�LPқ/��.�_SCT�CF_�`�Fb�l���|�FS8(!E�e�CHA�1��p4�D°"3�RSD��`$"}����_Tb��PRO����� EM�i_��a�8!�ac !�a��DIR0~�RAILACI�)RMr�LO��C����Qq��#q�դ�P�R=�S�A�pC�/�c 	��FUNCq�0rRINP�Q�0���2�!RAC �B ���[���[WARn���BL�Aq�aA����DAk�0\���LD0����Q��qeq�T�I"r��K�hPRIYA�!r"AF��Pz! =�;��?,`�RK����MǀI�!�DF_�@B�%1n�LM�F=Aq@HRDY�4_�P@RS�A�0� �MULSE@���a ��ưt�m�m�$�1$�1�$1o����o� x*�EG� ����!AR���Ӧ��09�2,%� 7�AX]E��ROB��WpA2��_l-��SY[�W!4‎&S�'WRU�/-91��@�STR����t��Eb� 	�%��J��AB� ���&9������OTo0 	$��ARY�s#2��4�Ԓ�	ёFI@��?$LINK|�qJC1�a_�#���%:kqj2XYZ��t;�rq�3�C1j2^8'0B��'�4����+ �3FI���7�q����'��_Jˑ��⣜O3�QOP_�$;5����ATBA�QBCL��&�DUβ�&6��TURN߁"r�E110:�p��9GFL�`_� ��* �@�5�*7��Ʊ� 1�� KŐM��&8���"r��ORQ��a�(@# p=�j�g�#qXU������mTOVEtQ:�M ��i���U��U��VW�Z�A�Wb��T{�,  ��@;�uQ���P\�i� �UuQ�We�e�SSERʑe	��E� O���UdAas��4S`�/7����AX�� B�'q��E1�e��i ��irp�jJ@�j�@�j �@�jP�j@ �j�!�f ��i��i��i��i ��i�y�y�'y��7yTqHyDEBU8�$32���qͲ0f2G + AB�����رnSVS�7� 
 #�d��L�#�L��1W� �1W�JAW��AW��AW� QW�@!E@?D2�3LAB�29U4�AӼ���C (o�E�Rf�5� � $��@_ A��!�PAO��à�0#���_MRAt�� d� � T��ٔER1R����;TY&����I��V�0�cz�TO	Q�d�PL[ �d�"��� 
��C! � pp`T)0���_V1Vr�aӔ�����2ٛ2�E����@�8H�E���$W���j��V!��$�P@��o�cI��aΣ	 �HELL_CFG�!� 5��Bo_BASq�SR3�\�� a#Sb�T��1�%��2��U3��4��5��6��e7��8���RO�����I0�0NL�\CAqB+�����ACK4� ����,�\@2@�&�?�7_PU�CO. U�OUG�P~ ����m�ذ�����TPհ_KcAR�l�_�RE*��P���7QUE����uP����CST?OPI_AL7�l��k0��h��]�l0SE�M�4�(�M4�6�T�YN�SO���DI�Z�~�A�����m_T}M�MANRQ���k0E����$KEYSWITCH��ص�m���HE��BE�AT��E- LE(~�����U��F!Ĳ�|��B�O_HOM=�OGREFUPPR�&��y!� [�C��O��-ECOC��Ԯ0_IOCMWD
�a����m��� � �Dh1���UX���M��βgPgCFORC<��� ^%>�m��OM.  � @��5(�U�#P, 1(��, 3��45���NPX_ASt��; 0��ADD����$SIZ��$�VAR���TIPR/�.��A�ҹM�@ǐ��/�1�+ U"S��U!Cz���FRIF���J�S���5Ԓ�N�F�� �� � x6p`SI��TE�C��.�CSGL��TQ2�@�&����� ��ST�MT��,�P �&ByWuP��SHOW4�Α�SV�$�w� �Q�A00�@ Ma}���� �����T&���5��6��7��8��9��A��O ��@�Ѕ�Ӂ���0��F�� � G��0G���0G����@G��PG��1�	1	1	1+	1�8	1E	2��2��2���2��2��2��2���2��2��2��2�	2	2	2+	2�8	2E	3��3��3���3��3��3��3���3��3��3��3�	3	3	3+	3�8	3E	4�4��4���4��4��4��4���4��4��4��4�	4	4	4+	4�8	4E	5�5��5���5��5��5��5���5��5��5��5�	5	5	5+	5�8	5E	6�6��6���6��6��6��6���6��6��6��6�	6	6	6+	6�8	6E	7�7��7���7��7��7��7���7��7��7��7�	7	7	7+	7�8	7E��VP��U�PDs�  �`NЦ�
>�YSL}Ot�� � L�`��d���A�aTA�80d��|�ALU:ed��~�CUѰjgF!aIgD_L�ÑeHI�j�I��$FILE_���d��$2�
�c;SA>�� hO��`?E_BLCK��b|$��hD_CPUy M�yA��c�o�d�b��ކ�R �Đ
P�W��!� oqLA®�S=�ts�q~tRUN�qst�q~t���p�qst�q~t �T���ACCs��Xw -$�qLEN;� �tH��ph�_�I��ǀLOW_AXI�SF1�q�d2*�MZ���ă��W�Im�ւ�a�R�TOR��pg�Dx�Y���LACEk��ւ�pV�ւ~�_MA�2�v�������TCV��؁��T��ي���@��t�V����V�Jj�R�MA�i�J��m�u�)b����q2j�#аU�{�t�K�JK��V�K;���H���3��J�0����JJ��JJ��AAL��ڐ��ڐ�Ԗ4Օ5���N1����ʋƀW�LP�_�(�g����pr��{ `�`GROUw`���B��NFLI�C��f�REQUI;RE3�EBU��qB���w�2����p��x�q5�p�� \��/APPR��C}�Y��
ްEN٨CLO7��S_M��H����u�
�qu�� ���MC�����9�_MG��C�Co��`M��в�N�BRKL�N�OL|�N�[�R��_CLINђ�|�=�J����Pܔ�����������������6ɵ�̲�8k�+��q����# ��
��q)��7�PATH3�L�BàL��H�wࡠ�J�CN�CA�Ғ�ڢB�IN�rUCV�4a��-C!�UM��Y,����aE�p����ʴ�~��PAYLOA���J2L`R_AN�q�Lpp���$��M�R_F2LSHR��N�LOԡ�R����`ׯ�ACRL_@G�ŒЛ� ��Hj`�߂$HM���FL�EXܣ�qJ�u� :�����׀�������1�F1�V�j�@�R�d�v�������E����ȏڏ ����"�4�q���6� M���~��U�g�y����T��o�X��H��� ���藕?�����ǟ ِݕ�ԕ����%��7��P��J�� � �V�h�z���`AT؃採@�EL�� �S��J|�Ŝ�JE�y�CTR��~�TN��FQ��HAND_VB-���v`�7� $��F2M��,��ebSW�q\�'��� $$MF�:�Rg�(x�,4�%��0&A�`�=��aM)�F�AW�Z`i�Aw�A���X X�'pi�Dw�Dʆ�Pf�G�p�)ST�k��!x��!N��DY �pנM�9$`%Ц�H� �H�c�׎���0� ��Pѵڵ����������J��� ����1��R�6��QA'SYMvř���v���J���cі�_SH >��ǺĤ�ED����������J�İ%��C��IDِ�_VI��!X�2PV_UNIX�FThP�J��_R�5 _Rc�cTz�pT�V��@�@��İ�߷��U ��������Hqpˢ���aEN�3�DI�����O4d�`J�S� x g"IJAA�a z�aabp�coc�`a�p�dq�a� ��OMME��� �b�RqAT(`PT�@� S��a7�;�Ƞ�@�h�a�i�T�@<� $D�UMMY9Q�$�PS_��RFC� 9 S�v �p���Pa� XƠ����STE���SBR�Y�M21_VF�8�$SV_ERF�O���LsdsCLRJtA���Odb`O�p �� D $GgLOBj�_LO����u�q�cAp�r�@aS;YS�qADR``�`TCH  �� ,��ɩb�W_NA���7����SR���l ���
*?�&Q�0" ?�;'?�I)?�Y)��X� ��h���x������)�� Ռ�Ӷ�;��Ív�?�ДO�O�O�DE�XS�CRE栘p��f��ST��s}y`�����/_HAΗq� TơgpTYP�b���G�aG�j��Od0IS_i䓀d�UEMdG� ����ppS�q�aRSM_�q*eU?NEXCEP)fW�`S_}pM�x���g�pz�����ӑCOU��S�Ԕ 1�!�U�E&��Ubwr��PR�OGM�FL@7$CUgpPO�Q���5�I_�`H� �� 8�� �_HE��PS�#��`RY ?�qp�b��dp��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI@m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1 �ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS���>4�VSHIF��Nc�P�`ג�E�ȐyR����OSUR��=Wk`RADILѮ��_�a��:�9a��`a��r��LULQ$O�UTPUT_BM����IM�AB �@��rTILSC	O��C7��� ����&��3��A����q���m�I�2$G�ϑV�pLe�}��y�DJU��N�WAIT֖�}��{��%! NE�u�YB�O�� �� c$`�t�SB@wTPE��NECp��J^FY�nB_T��R�І�a$�[Y��cB��dM���F�� �p�$�pb�OP�?�MAS�_DO*�!QT�pD��ˑ�#%��p!"DELA1Y�:`7"JOY�@( �nCE$��3@ �xm��d�pY_[�!"�`��"��[���P? {T`ZABC%�?�  $�"R���
ϐ�$$CL�AS�������!pϐ� � VIRqT]��/ 0ABS�����1 5�� < �!F?X?j?|?�?�? �?�?�?�?�?OO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�o�o�o  $6HZi{0-�GAXL�p��"�637  �{tIN��q�ztPRE�����v��p�uLARMRE?COV 9�r�wtNG�� .;	? A   �.��0PPLIC��?�5�p��Handling�Tool o� �
V7.50P/�23-�  �Pz���
��_SW�t� UP�!� �x�F0��t�Qz�Aϐv� 8[64�� �it��y�2�2 �7DA5�� [�� d��@���o�Noneisͅ�˰ ��T����!�Ayx�>�_l�V�uT��s9�UTO�"�Њt�y~��HGAPON
0�g�1��Uh�D 1-581�����̟ޟry����Q 1���p�,�� ����;�@��q_��"��" ��c�.�H���D�?HTTHKYX��" �-�?�Q���ɯۯ5� ���#�A�G�Y�k�}� ������ſ׿1���� �=�C�U�g�yϋϝ� ������-���	��9� ?�Q�c�u߇ߙ߽߫� ��)�����5�;�M� _�q�������%� ����1�7�I�[�m� ���������!���� -3EWi{� �����) /ASew��� �/��/%/+/=/ O/a/s/�/�/�/�/? �/�/?!?'?9?K?]? o?�?�?�?�?O�?�?`�?O#O]���TO��E�W�DO_CLE�AN��7��CNM ; � �_�_/_A_S_�DSP�DRYR�O��HIc��M@�O�_�_�_�_ oo+o=oOoaoso�o`�o���pB��v �u���aX�t������9�PLUGG���G���U�PRCvPB�@"��_�orOr_^7�SEGF}�K[ mwxq�O�O����8�?rqLAP�_�~ q�[�m��������Ǐ�ُ����!�3�x�T�OTAL�f yx�U�SENU�p�� ��H���B��RG_S�TRING 1~u�
�Mn��S5�
ȑ_ITwEM1Җ  n5� � ��$�6�H�Z�l� ~�������Ưد����� �2�D�I/�O SIGNAL�̕Tryou�t Modeӕ�Inp��Simu�latedבO�ut��OVE�RR�P = 10�0֒In cy�cl��בPro?g Abor��ב���Status�Փ	Heartb�eatїMH �Faul��Aler'�W�E�W�i�{���ϟϱ������� �CΛ�A����8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j�|���WOR{pΛ�� (ߎ����� ��$�6� H�Z�l�~���������������� 2PƠ�X ��A{� ������ /ASew���8��SDEV[� o�#/5/G/Y/k/}/ �/�/�/�/�/�/�/?�?1?C?U?g?y?PALTݠ1��z?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O8�O_�?GRI�`Λ DQ�?_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o2_l�R��a\_�o"4 FXj|���� �����0�B�T��oPREG�>��  f���Ə؏���� � 2�D�V�h�z��������ԟ���Z��$A�RG_��D ?	����;���  	]$Z�	[O�]O���Z�p�.�SBN_�CONFIG �;�������C�II_SAVE � Z�����.�T�CELLSETU�P ;�%H?OME_IOZ�Z�?%MOV_���
�REP�lU�(�U�TOBACKܠ���FRA;:\z� \�z�Ǡ'`�z���n�WINI�0z����n�MESSAG༠�ǡC���ODEC_D������%�O��4�n�PAUSX!��;� ((O >��ϞˈϾϬ����� �����*�`�N߄��rߨ߶�g�l TSK�  w�Կ׿q�UgPDT+��d!�~A�WSM_CF���;���'�-�G�RP 2:�?� �N�BŰA��%�XS�CRD1�1
7� �ĥĢ������ ����*�������r� ����������7���[� &8J\n��|*�t�GROUN�|UϩUP_NA��:�	t��_E�D�17�
 ��%-BCKED�T-�2�'K�`�Ƣ�-t�z��q�q�z���2 t1�����q�kp�(/��ED3/ ��/�.a/�/;/M/ED4�/t/)?�/.p?p?�/�/ED5`? ?�?<?.�?O�?�?ED6O�?qO�?.pMO�O'O9OED7�O `O_�O.�O\_�O�O�ED8L_,�_�^�-�_ oo_�_ED!9�_�_]o�_	-9o�oo%oCR_  9]�oF�o�k� � ?NO_DEL���GE_UNUSE���LAL_OU�T ����W?D_ABORﰨ~���pITR_RT�N��|NONS�k���˥CAM�_PARAM 1�;�!�
 8
�SONY XC-�56 23456�7890 �~��@���?��( А\�
����{����^�HR5pq�̹��ŏR57ڏ��Aff��K�OWA SC31�0M
�x�̆�d @<�
��� e�^��П\�����*�<��`�r�g�CE�_RIA_I�j!�=�F��}�vz� ��_LIU�Y]�����<���FB�GP 1��Ǯ�M�_�q��0�C*  ����CU1��9��@��G��Z�CR�C]��d��l��s��R�����U[Դm��v����}����� C���ő(�����=�HE�`ONFIǰ�B��G_PRI 1�{V���ߖϨϺ�����������CHK�PAUS�� 1K� ,!uD�V�@� z�dߞ߈ߚ��߾��� ���.��R�<�b���O��������_MOR�� y�6��� 	 �� ���*��N�<����"���?��q?;�;�I���K��9�P����ça�- :���	�

��M����pU�ð��<��,,~��DB���튒�)
mc:cpm�idbg�f�:����q���c�p��/�  �*9 �9 �� ��s>�0��0�ҰU�?��pH��pIUg�/��
�p�Uf�M/w�O/~�
DEF l���s)�< buf.txts/�t/��ާ�)�	`���ޛ�=L���*MC��1����?43���1��t�īC�z  B�J�B���_C|��Cq�CG�eC�?��CTyY
K��D6��F.���F��E⚵F,E�ٟ��K�F6�*IU���I?O�I<�#I6�I慴Y	?3���#w�1����s���.*�p������BDw��M@x8�K�C�C�����D�p@�E�YK�EX�E�Q�EJP F��E�F� G���>^F E��� FB� H�,- Ge��H�3Y��:�  >�33 ���N~  n8�~@��#5Y�E>�ðA��Yo<#�
"Q ����+_�'RSMOF�S�p�.8��)T1>��DE ��F� 
Q��;�(P � B_<_��R��X��	op6C4P�Y
�s@ ]AQ�2s@CR�B3�MaC{@@*c�w��UT�pFPROG %�z�o�o�igI�q���v��ldK�EY_TBL  ��&S�#� �	
��� !"#�$%&'()*+�,-./01i�:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������vq���͓���������������������������������耇���������������������p`LCK�l4�p`�`�STAT ��S_A�UTO_DO����5�INDT_ENB!���R�Q?�1��T2}�^�STOP�b���TRLr`LE�TE��Ċ_SCREEN �Z�kcsc��U���MMENU 1� �Y  < �l�oR�Y1�[���v� m���̟�����ٟ� 8��!�G���W�i��� �����ïկ��4�� �j�A�S���w����� 迿�ѿ����T�+� =�cϜ�sυ��ϩϻ� ������P�'�9߆� ]�o߼ߓߥ������ ��:��#�p�G�Y�� ����������$��� �3�l�C�U���y��� �������� ��	V�Y)�_MANUAyL��t�DBCO[��RIGڇ
�DBN�UM� ��B1 e
��PXWORK 1!�[�_U/�4FX�_AWA�Y�i�GCP r b=�Pj_AL� #�j�Y��܅ `��_�  1"�[ , 
�mt7�&/�~&lMZ�IdPx@|P@#ONTIMه�� d�`&�
��e�MOTNEN�D�o�RECOR/D 1(�[g2�/{�O��!�/ky "?4?F?X?�(`?�?�/ �??�?�?�?�?�?)O �?MO�?qO�O�O�OBO �O:O�O^O_%_7_I_ �Om_�O�_ _�_�_�_ �_Z_o~_3o�_Woio {o�o�_�o o�oDo�o /�oS�oL�o ����@��� +�yV,�c�u���� ����Ϗ>�P����� ;�&���q���򏧟�� P�ȟ�^������I� [����� ���$�6��������jTOL�ERENCwB����L�͖ CS_CFG )��/'dMC:\�U�L%04d.C�SV�� c��/#A� ��CH��z� �//.ɿ��(S�RC_OUT *���1/V�SGN �+��"��#��19-FEB-20 08:010�17l�19:09�+ PQ�8�ɞ�/.��f�pa��m��PJP�Ѳ��VERSI�ON Y��V2.0.84,E�FLOGIC 1�,� 	:�ޠ=�ޠL��PROG_ENB��"p�ULSk' ����_WRSTJNK ���"fEMO_O�PT_SL ?	��#
 	R575/#=������0�B����TO  a�ݵϗ��V_F �EX�d�%��P�ATH AY�A�\�����5+IC�T�Fu-�|j�#egS��,�STBF_TTS�(�	d���l#!w�� MAU��z�^"�MSWX�.�<�(4,#�Y�/�
!J� 6%ZI~m���$SBL_FAU�L(�0�9'TDI�A[�1<�<� ����1234567890
��P��HZl~�� �����/ /2/�D/V/h/�� P� ѩ�yƽ/��6 �/�/�/??/?A?S? e?w?�?�?�?�?�?�?8�?�,/�UMP����3 �ATR��Ӝ1OC@PMEl�OOY�_TEMP?�ÈÓ3F���G�|DUN�I��.�YN_BR�K 2_�/�EMGDI_STA���]�'�@NC2_S_CR 3�K7 (_:_L_^_l&_�_�_`�_�_)��C�A14_ �/oo/oAoԢ�B�T5�K�ϋo~o l�{_�o�o�o' 9K]o���� �����#�5��/ V�h�z��л`~����� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T��� x���������ү��� ��,�>�P�b�t��� ������ο���� (�f�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������:� �2�D�V� h�z���������� ��
��.�@�R�d�v� ������������� *<N`r�� �����& 8J\n����� �����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?��?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__�NoETMODE �16�5�Q �d�X
X_j_|Q��PRROR_PR�OG %GZ%��@��_  �UTAB_LE  G[�?�oo)oRjRRSE�V_NUM  <�`WP�QQY`��Q_AUTO_ENB  �eOS�Tw_NOna 7G[��QXb  *�*�`��`��`��`d`�+�`�o�o�o�dHI�SUc�QOP�k_AL�M 18G[ �2A��l�P+�ok@}�����o_Nb.�`  G[�a�R�
�:PTCP_VE/R !GZ!�_��$EXTLOG_7REQv�i\��SIZe�W�TOL�  �QDzr��A W�_BWD��p��xf́t�_DIn�� 9�5�d��T�QsRֆSTEP���:P�OP_D�Ov�f�PFAC�TORY_TUN�wdM�EATUROE :�5̀rQ�Handl�ingTool ��� \sfm�English �Dictiona�ry��roduAA Vis�� Master��ީ�
EN̐nalog I/O��ީ�g.fd̐ut�o Softwa�re Update  F OR��matic Ba�ckup��H59�6,�ground Editޒ�  1 H5�Camera�F���OPLGX�elyl𜩐II) X�7ommՐshw���7com��co����\tp���pan}e��  opl���tyle sel�ect��al C�nJ�Ցonit;or��RDE���tr��Relia�b𠧒6U�Dia�gnos(�푥�5�528�u��he�ck Safet�y UIF��En�hanced Rob Serv%��q ) "S�r�U?ser Fr[������a��xt. D�IO �fiG� �sŢ��endx�Ekrr�LF� pȐ�ĳr됮� ���� � !��FCTN /Menu`�v-�ݡ|���TP Inې�fac�  ER_ JGC�pב_k Exct�g���H558��igh�-Spex�Ski~1�  2
P���?���mmunic�'�ons��&�l�uqr�ې��ST Ǡ���conn��2ި�TXPL��nc=r�stru�����"FATKA�REL Cmd.� LE�uaG�54�5\��Run-T�i��Env��d�
!���ؠ++�s�)�S/W��[�LicenseZ��� 4T�0�ogB�ook(Syڐm�)��H54O�MA�CROs,\�/O�ffse��Loa��MH������r,� k�MechStop Prot����� lic/�MiвShif����ɒ�Mixx��)���,�e�S�Mode �Switch�� �R5W�Mo�:�.�� 74 ����g��K�2h�ult�i-T=�M���LN (Pos�Regiڑ������|d�ݐt Fun��⩐.�����Numx~����� lne�|�ᝰ Adjup������  - W���tatuw᧒T��RDMz�o}t��scove U�9���3Ѓ�uest 492�b*�o�����62;�?SNPX b ����8 J7`���Li3br��J�48����"�� �Ԅ�
�6O��� Parts i�n VCCMt�3�2���	�{Ѥ�J9�90��/I� 2� P��TMILI�B��H���P�A�ccD�L�
TE�$TX�ۨ�ap1�S�Te����pke�y��wգ�d���Unexcep=tx�motnZ���������є�� qO���� 90J��єSP CSXC`<�f��Ҟ� Py�sWe}���PRI��>vr�t�menz�� ��iPɰ�a�����vGri=d�play��v���0�)�H1�M-�10iA(B20�1 �2\� 0\}k/�Ascii��l�Т�ɐ/�Col���ԑGuar� �
�� /P-�ޠ"Kv��st{Pat �:�!S�Cyc��΂�orie��IFn8�ata- quҐ��� ƶ��mH57m4��RL��am����Pb�HMI D�e3�(b����PC�Ϻ�Passwo�+!��"PE? Sp�$�[���tp��� vKen��Tw�N�p��YELLOW B�OE	k$Arc��v�is��3*�n0W�eldW�cialh�7�V#t�Op�����1y� 2F�a�portN�(�p�T1�T� �� �ѳxy]�&TX��t�w�igj�1� b� �ct\�JPN �ARCPSU P�R��oݲOL� S;up�2fil� &�PAɰאcro�� �"PM(����O$SuS� eвtex�ԣ r���=�t�s'sagT��P���P@�Ȱ�锱�rt�W��H'>r�dpn��n1
t�!�� z ��ascbi?n4psyn��+A}j�M HEL��NCL VIS �PKGS PLOA`�MB �,�4�VW�RIPE �GET_VAR {FIE 3\t���FL[�OOL: �ADD R729.FD \j8'�iCsQ�QE��DVvQ��sQNO WTW�TE��}PD  D�p��biRFOR ���ECTn�`��ALSE ALAfP�CPMO-130�  M" #h�D�: HANG F�ROMmP�AQfr���R709 DR�AM AVAIL?CHECKSO!���sQVPCS SU��@LIMCHK �Q +P~dFF PO�S��F�Q R59�38-12 �CHARY�0�PR�OGRA W�SwAVEN`AME�P�.SV��7��$E�n*��p?FU�{�TR}C|� SHADV0�UPDAT KC|JўRSTATI�`~�P MUCH y��1��IMQ MO?TN-003��}��ROBOGUIDE DAUGH�a8���*�tou�����I� Šhd�ATH|�PepMOVET��ǔVMXPACK� MAY ASS�ERT�D��YCL�fqTA�rBE C�OR vr*Q3rA�N�pRC OPToIONSJ1vr̐PSH-171Z@-x�tcǠSU1�1`Hp^9R!�Q�`_T�P���'�j�d{tb�y app wac 5I�~d�PHI����p�aTEL�MX?SPD TB5bLu� 1��UB6@�qEN�J`CE2�61��p���s	�may n��0� R6{�R� >�Rtraff)��� 40*�p��fr���sysvar ?scr J7��cNj`DJU��bH �V��Q/�PSET �ERR`J` 68���PNDANT �SCREEN U�NREA��'�J`D��pPA���pR`IgO 1���PFI�p}B�pGROUN�P�D��G��R�P�QnRS�VIP !p�a�PD�IGIT VER�S�r}BLo�UEW~ϕ P06  �!��MAGp�abZV��DI�`� SS�UE�ܰ�EPL�AN JOT` D�EL�pݡ#Z�@D�͐CALLOb�Q �ph��R�QIPN�D��IMG�R7{19��MNT/�PWES �pVL�c���Hol�0Cq���tP�G:�`C�M�caynΠ��pg.v�S�: 3D mK�v_iew d�` �p���ea7У�b� o�f �Py���ANN�OT ACCESGS M��Ɓ*�t47s a��lok��Flex/:�Rw�!mo?�PA?�-�����`n�pa S�NBPJ AUTO-�06f����TB���PIABLE1q �636��PLN:Y RG$�pl;pNW7FMDB�VI���t�WIT 9x�0@o���Qui#0�ҺPN� RRS?pUSB��� t & remov�@ )�_��&�AxEPFT_=� �7<`�pP:�OS�-144 ��h qs�g��@OST� �� CRASH �DU 9��$�P�pW� .$��L/OGIN��8&�J���6b046 issue 6 Jg���: Slow ��st��c (HCos`�c���`IL`�IMPRWtSPO�T:Wh:0�T�S�TYW ./�VMGqR�h�T0CAT��hos��E�q���� �O�S:+pRSTU' k�-S� ����E:��pv@�2�N� t\hߐ��m ���all��0�  �$�H� WA͐��3 CNT0 T��� WroU�alacrm���0s�d � @�0SE1���r R{�OMEBp���K� �55��REàSEs�t��g    } �KANJI��no���INIS?ITALIZ-p�d�n1weρ<��dr�� lx`�SCI�I L�fail�s w�� ��`�YSTEa���o��PvЧ IIH���1W�G�ro>Pm ol\�wpSh@�P��Ϡn� cflxL@АW{RI �OF Lq���p?�F�up��d�e-rela�d� "APo SY�c}h�Abetwe:0IND t0$gb#DO���r� `��GigE�#ope�rabilf  P�AbHi�H`��c�le{ad�\etf�P8s�r�OS 030��&: fig��GL�A )P ��i��7�Np tpswx�B��If�g�������5aE�a EXC�E#dU�_�tPCLO�S��"rob�NTdpFaU�c�!����PNIO V750�Q1��Qa��'DB ��P M�+Pv�QED�DET���-� \rk��ON�LINEhSBUG�IQ ߔĠi`Z�IB�S apABC �JARKYFq� ����0MIL�`� R��pNД �p0GAR��D*pR��P�"'! jK�0cT�P��Hl#n�a�ZE V��� TASK�$VP2(�4`
�!�$�P��`WIBPK05��!FȐB/��BUSY RUNN��C "�򁐈��R-p��LO�N�DIV�Y�CUL��fsfoaBW�p����30	V��ˠIT�`�a505.�@O=F�UNEX�P1bҬaf�@�E��SVwEMG� NMLq�� D0pCC_SA�FEX 0c�08"qD. �PET�`N@�#'J87����RsP�TA'�M�K�`K��H GUNCHG^۔MECH�pMcz� T�  y, g@��$ ORY LE�AKA�;�ޢSP�Em�Ja��V�tGR�Iܱ�@�CTLN�TRk�FpepR��j50�EN-`IN�����p �`�Ǒ�k!��T3/dqo�SKTO�0A�#�L�pA �0�@�Q�АY�&�;pb1TO8pP�s����FB�@Yp`�`D	U��aO�supk�t4� � P�F� Bnf��Q�PSVGN-18��V�SRSR)J�UP�a2�Q�#D�q� l O��QBRKCTR5Ұ�|"-��r�<pc�j!INVP�D ZO� ��T`�h#�Q�cHset,x|D��"DUAL� �w�2*BRVO117 A]�TNѫt�+bTa2473��q.?���r�{1 009�.fd8�y`j60�4.\P-�`han�c�U� F��eN8��  ��npJtPpd!q��`��� 5h'596p�!5d�� @"p�P�P�Q�0�P2�p �A� \P��R(}\\P�e� aʰI���E���1��p� j  �� ,e?�Dp� �A��A\P�q 5 sig:��a��"AC;a���
�bCe\Pb_p���.pc]l<bHbc?b_circ~h<n�`tl1�~`\P`o�d�\P�b]o2�� �cb��c�i\P�jupfr�m�d\P�o�`exe��a�oFd\Ptped�}o��u`�cptli1bxz\P�lcr�xr\P\�blsazEd\P_fm�}gc\P�x�� �o|sp�o�mc(��o'b_jzop�u6��wf��t��wms�1�q��sld�)��jm!c�o\�n��nuhЕ�ƭ|st�e��>�pl�qp�iwck���u�vf0uߒ��lvi�sn�CgaculwQ
E `RFciV\P�qiP��Data Acquisi��ynZU�SR631`���TR�QDMCM Z�2�P75H�1�P�583\P1��71֫�59`�5�P57@<P\P�Q����(����Q��o p\P!daq\�oA��@��� ge/�etdm~s�"DMER"؟�,�pgdD���.�mp���-��qaq.<ጡ�\Pmo��h���f�{�oR503��MA�CROs, Sk�saff�@lR���03��SR�Q(��Q6��1"�Q9ӡ�R�ZSh��P^\PJ643�@7ؠ�6�P�@�PRS�@����e �Q�UС PI�K�Q52 PTLqC�W��\P3 (��p/O��!�Pn ��\P5��03\s�fmnmc "M�NMCq�<��Q��\$AcX�FM���ci ,Ҥ�X����cdpq+�6
�sk�SK�\P�SH560,P���,�y�refp "GREFp�d�A�j\P6	�of�OFc�<g6y�to�TO_���<�ٺ���+je|�u��caxis2��\PE�\�e�q"IS�DTc��]�prax ��MN��u�b�isde܃h�\��iR\P! isba�sic��B� P�]��QAxes�R�6������.�(Ba�Q�ess��\P����2�D�@�z�atis���(�{����h��~��m��FMc��u�{�
ѩ�MNIS ��ݝ����x�����ٺ��jW75��De�vic�� Interfac�RȔQJ754��� \P�Ne`��\P�ϐ`2�б����dn� �"DNE���
t�pdnui5UI��ݝ	bd�bP>�q_rsofOb~
dv_aro��u�����stchkc��z	 �(�}onl��G!ffL+H�J(��"l"�/�n�b��z�h�amp��T�C�!i�a"�59��S�q��0 (�+P�o�u�!�2��xpc_2pcc{hm��CHMP_�|8бpevws��2�쳌pcsF��#C� Sen\Pacrao�U·�-�R6�P�d�\Pk�����p��g8T�L��1d M�2`���8�1c4ԡ�3 qem��GEM,\i(�>�Dgesnd�5��`�H{�}Ha�@sy����c�Isu�xD��Fmd��I��7�4���u����AccuCal �P�4t@��ɢ7ޠBU0��6+6f�6��C99\aFF q�S(�U��2�
X�p�!Bdf��cb_�SaUL��  �t@?�ܖt�o��otplus\tsrnغ�qb��Wp��t���1��T�ool (N. �A.)�[K�7�Z�(P�m����bfc�lst@k94�"Kp4p��qtpap�� "PS9H�stpswo��p�L7��t\�q����D�yt 5�4�q��w�q��t@��M�uk��rkey�����s��}t�sfoeatu6�EA��t@cf)t\Xq�����̜d�h5���LR0C0�md�!�587���aR�(����2V���8c?u3l\�pa�3}H�&r-�Xu���t,�t@�q "�q�Ot� �~,���{�/��1c�}����y�p�r��5� ��S�XAg�-�y���W�j874�- i�RVis���Queu�t@Ƒ�-�6H�1���(����u����tӑ����
�tp�vtsn "VTCSN�3C�+�t@v\p�RDV����*�pr�dq\�Q�&�vs�tk=P������n�m&_�դ�clrq8ν���get�TX��Bd���aoQϿ�0qstr�D[t@��at�p'Z����npv��@�enlIP0��`D!x�'�|���sc ����tvo/��2�q���vb����q ���!���h]��(�� Control^�PRAX�P5��g556�A@59�P[56.@56@5A��J69$@982� J552 IDVR7�hqA���16��H���La�� ���Xe�frlpa�rm.f�FRL��am��C9�@(F�����w6{���A<��QJ643�t@�50�0LSE
�_pVAR $SG�SYSC��RS_?UNITS �P�2��4tA�TX.$V�NUM_OLD �5�1�| {�50�+�"�` Funct���5tA� }��`#@��`3�a0�cڂ��9���@H5נt@�P���(�A����۶�}����ֻ}��bP�Rb�߶~ppr4�TPSPI�3�}�r�10�#;A� t�
`��2�1���96����@�%C�� Aف��J�bIncr�	����\����1o5qni4�MNINp	�t@���!��Hour�  � �2�21 ��AAVM���0y ��TUP ��J545 ���6162�V�CAM  (��CLIO ���R6�N2�MS�C "P ��STYL�C�2�8~ 13\�NRE "FHRM �SCH^�DC�SU%ORSR �{b�04 �oEIOC�1 j o542 � os| ~� egist������7�1��MASK�93�4"7 ��OCO) ��"3�8��12���� 0 HB���� 4�"39N� �Re�� �LCH=K
%OPLG%��3"%MHCR.%M�C  ; 4? ��6 6dPI�54�s� �DSW%MD� pQ�K!637�0�0p"��1�Р"4 �6~<27 CTN K V� 5 ���"7���<25�%/�T�%FRDM� �Sg!���930 FB( NB�A�P� ( HLB o Men�SM$@<jB( PVC ��s20v��2HTC�~CTMIL��~\@PAC 16U��hAJ`SAI \@EL�N��<29s�U�ECK �b�@FR3M �b�OR����IPL��Rk0CS�XC ���VVF�naTg@HTTP ��!26 ��G��@obIGUI�"%IPGS�r� H863 qb�!�07rΈ!34 �r�84 \so`! Qx`CC�3 Fb�21�!9s6 rb!51 ����!53R% 1!s(3!��~�.p"9js �VATFUJ775�"��pLR6^RP�W;SMjUCTO�@xT158 F!80���1�XY ta3!770� ��885�UO	L  GTSo
�{` �LCM �r| TS�S�EfP6 W�\@C�PE `��0VR�� l�QNL"��@001 imrb�c3 =�b�0���0�`�6 w�b-P- Ru-�b8n@5EW�b9 �Ґa� ���b�`�ׁ�b2 2000$��`3��`4*5�`A5!�c�#$�`7.%~�`8 h605? ;U0�@B6E"aRpm7� !Pr8 t��a@�tr2 iB�/�1vp3�vp5 �Ȃtr9Σ�a4@-�p�r3 F��r5`&�re`u��r7 ��r8�U�p9 \h�738�a�R2DK7"�1f��2&�y7� �3 7iCЊ�4>w5Ip�Or6�0 C�L�1bEN�4 I�pyL�uP��@LN�-PJ8�N�8Ne�N�9 H�r`�E"�b7]�|���8�В����9 2��a`0�qЂ5�%U097 0��@1�0����1 (�q�3 5R���0���mpU��0�0�7*�H@x(q�\P"RB6�q124�b;��@���f@06� x�3 p�B/x�u ��x�6 /H606�a1� ����7 6 ���<p�b155 ����}7jUU162 ��3 g��4*�6?5 2e "_��PF�4U1`���B1��z�`0'�174 �q���P�E186 R� ��P�7 ��P�8�&�3 (�90 B/�s191����@�202��6 30���A�RU2� d���2 b2h`��4Ģ᪂2�4���19�v Q�2��u2d�TRpt2� ��H�a2hPd�$�5���!U2�pD�p
�2�p��@5�0H-@��8 @�9��TX@�� �e5�`rb26Af�2^R�a�2 Kp��1y�b5Hp�`

�5�0@�gqGA��F�a52ѐ�Ḳ6�K60ہ5� ׁ2��i8�E��9�EU5@�ٰ\�q5hQ`S�2
ޖ5�p\w�۲�pJh �-P��5�p1\t�ZH�4��PCH�7j��phiw�@��P�x�~�559 ldu�  P�D���Q�@�������� �`.��P>��8��581�"�q58�!AM۲T�A iC�a589��@�x�����5 �a��12@׀0.�1���,�2��8��,�!P\h8��Lp� ��,�7��6�08�40\t� "T20C}A��p��{��ran��FRA ��Д�е���A% ���ѹ�Ҁ�����( ����Ѐ���З��� ������р����$�!G��1��ը���������� ,e�`q�  �����`�64��M��iC/50T-H������*��)p46��� C���N����m75s�֐� Sp�ѯb4�6��v����ГM-71?�7�З�����42������C��-��а�70�r�E��/h����O$���rD���c7c7C@�q��Ѕ���L���/��2\imm7c7�g������`���(��e����� "�������a r�L�c�T,�Ѿ�"��,�� ��x�Ex�m77t���k���a5�����)�iC��-HS-� B
_�@>���+�Т�7U��]���Mh7�s�7������-9~?�/260L_� �����Q������4��]�9pA/@���q�S�х鼔��h621��c��92������.�)92c0�g$�@ �����)$��5$����pylH"O"
�21p���t?�350� ���p��$�
��� �350!���0���9�U/0\m9��M9A3��4%� s�3M$��X%yu���"him98 J3����� i d�"m4~�103p�� �Ӏ�h794̂�&R���H�0����\���g� 5A���Ԝ��0���*2@��00��#06�`�АՃ�է!07{r ��������kЙ @����EP�#�� ����?��#!�;&�07\;!�B1P��߀A��/ЁCBׂ2��!�:/��?�ҽCD2C5L����0�"l�2BL
#��B��\20�2_�r�re ���X��1��N����A$@��z��`C�p0U��`�04��DyA�\�`fQ����sU���\�5  ���� p�Dp���<$85���+�P=�ab1l�1LT��lA8�!uDnE\(�20T��J�1 e�bH85���b����5[�16Bs��������d2��x��m6t!`Q�����bˀ���b#�(�6iB;S�p�!��3� � ��b�s��-`�_�Wa8�_����6I	$2�X5�1�U85��R�p6S����/�/+q��!�q��`�6o��58m[o)�m6sW��Q��?��set06�p ��3%H�5��10�p$����g/�JrH~��  ��A�856����F�� ���p/2��� ��܅�✐)�5��̑v0��(��m6��Y�!H�ѝ̑m�6�Ҝ���a6�DM����-S�+��H2������ ��� �r̑��✐0��l���p1���Fx���2�\t6h T6H����Ҝ�'V l���ᜐ�V7ᜐP/����;3A7��@p~S��������4�`@圐�V���!3��2�PM[��%ܖO�7chn��vel5�p���Vq���_arp#���̑�.���2l_�hemq$�.�'�6415���5���?�� ��F�����5g�L�ј[���1��𙋹y1����M7NU�@�М��eʾ����uq$D;��-�4��3&H�f�c�Ĝ�h����� �u���㜐��`ZS�!ܑ4���M-����S�$̑�ք �� �0��<�����07shJ�H�v�À�sF ��S*󜐳���̑�� �vl�3�A�T�#��`QȚ�Te��q�pr��,��T@75j�5�dd� ̑1�(UL�&�(�,����0�\�?���̑�a��? ,e����a��e�w�2��(�	�2�C��A/���\�+px�����21 (ܱ�CL S����B�̺��7F���?�<�lơ1L����c� ��b�u9�0����e/q���O���9�K��r9 (��,�Rs�ז�x5�G�m20c��i��w�2��:�0`�$��2�2l�0�k�X�S� ,�ι2��O����1!41w���2<T@� _std��G��y� �ң�H� jdgm����w0\� �1 L���	�P�~�W*�b��t 5������%3�,���E{�������L��5\L��3�L�|#~���~!���4�#��O����h�L6A������2璥���44������[6\j4s��·���#��ol�E"w�8Pk�����?0 xj�H1�1Rr�>��6]�2a�2Aw�P ��2��|41�8��ˡ���{� �%�A<���  +�?�l��0�&�"��|�`Am1�2��ػ��3�HqB��K�R� �ˑb�W���Fs��� �)�ѐ�!���a�1��ڛ�5��16�16�C��C����0\imBQ��d����b���\B5�-���DiL ���O�_�<ѠPEtL�E�RH�ZǠPgω�am1l��u���̑��b�<����<�$�T �̑�F����Ȋ�D�pb��X"��hr��pw� ��Dp����9�0\� j971\kckrcfJ��F�s�����c��e "CTME�r��������a�`main.p[��g�`run}�_vc�#0�w�1O�ܕ_u����bctm�e��Ӧ�`ܑ�j7�35�- KAREL Use {�	U���J��1��
�p� Ȗ�9�B@���L�9��7j[�a�tk208 "KP��Kя��\��9���a��̹����cKRiC�a�o ��kc�q J�&s�����Grſ� fsD��:y��s��A1X3\j|хrdtB�,� ��`.v�q�� ��sǑIf�Wfj52��TKQuto S�et��J� H5nK536(�932�Z��91�58(�9�BA�1(�74O,A$�?(TCP Ak��В/�)Y� �\t�pqtool.v��v���! co�nre;a#�Control Re��ble��CNRE (�T�<�4�2���D�)����S�552��q(g�� (򭂯4X�cO�ux�\sfuts�UTS`�i�栜����t�棂��? 68�T�!�SA OO+D6���������,!��6c+� ig.t�t6i��I0�TW8 ���la��vo58�o�bFå򬡯i�Xh��!Xk�0Y!�8\m6e�!6EC���v��6���������<16�A���A�6s����U�g�TX|ώ���r1�qR��˔Z4�T�����,#�eZp)g����<O NO0���uJ��tCR;�x�F�a� ,e��f���prdsuchk �1��2&&?���	t��*D%$�r(��@���娟:r��'�s�q8O��<scrc�C�<\At�trldJ"�o�\�V����Pa�ylo�nfir1m�l�!�87��7� �A�3ad�! ��?ވI�?plQ��3���3"�q��x p�l�`���d7��l�calC�uDu���;���mov�����i'nitX�:s8O�p�a�r4 ��r67A4�|�e GenerGatiڲ���7g2�q$��g R� (#Sh��c ,|�bE��$Ԓ\�:�"��4��4�4�. sg��5�F$d6�"e;Qp "SH�AP�TQ ngcr pGC�a(�&"<� ��"GDA¶��r6�"aW�/�$�dataX:s�"t�pad��[q�%tput;a__O7;a�o8(�1�yl+s�r�?�:H�#�?�5x�?�:c O��:y O�:�IO�s`O%g�qǒ�?�@08\��"o�j92;!�P�pl.Colli=s�QSkip#��@ 5��@J��D��@\ވP�C@X�7��7��|s2��ptclsF�LS�DU�k?�\_ ets�`�< \�Q��@���`dc�KqQ�FC;��J,�n��` (��4eN����T�{��� 'j(�c�����/IӸaxȁ��̠H������зa�e\mc�clmt "CL�M�/��� mate�\��lmpALM0�?>p7qmc?����2vm�q��%�3s���_sv90�_x_m#su�2L^v_� K�o�{in�8(3r<�c_logr�N�rtrcW� �v_3�~yc��d��<�te��derv$cCe� Fiρ�R��Q�?�l�enter߄|��d(Sd��1�TX�+�fK�r�a99sQ9x+�5�r\tq\�� "FNDR����STDn$�LANG�Pgui��D⠓�S����Ơ�sp�!ğ֙uf �ҝ�s����$�����e+�=����������ࠓ���w�H�r\f�n_�ϣ��$`x�tc�pma��- TC�P�����R638� R�Ҡ��38
��M7p,���Ӡ�$Ӏ��8p0Р�VS,�>�tk��99�a��B3�� �PզԠ��D�2�����UI��t���hqB���8��������p���rqe�ȿ��exe@ 4φ�B���e38�ԡG��rmpWXφ�var@�φ�3N������vx�!ҡ��q��RBT $cO�PTN ask �E0��1�R MA�S0�H593/�9�6 H50�i�48
0�5�H0��m�Q�QK��7�0�g�Pl��h0ԧ�2Ҧ�D�P��@"��t\mas��0�a��"�ԧ�����k�գR�����¹`m��b��7�.f���u�d��r��splayD�E���1>w�UPDT Ub���887 (��Di{���v�Ӛ�Ԛ⧔���#�B��㟳��o  ����a�䣣��60q��B����qscan��B����ad@�������q `�䗣�#��К�`2�� vlv��Ù�`$�>�b���! S���Easy/К�U�til��룙�51G1 J�����R7 Θ�Nor֠��inGc),<6Q�� �`�c��"4�[���98Q6FVRx So����q�nd6����P�� 4�a\ (��
  ����D���d��K�bdZ����men7���- Me`tyFњ�Fb¨0�TUa�57	7?i3R��\��5�u?��!� n����f������l\mh�Ц�űE|Ghmn�	��<\HO���e�1�� l!D��y��Ù�\|�p����B���Ћmh�@��:.aG! ���/�t�55�6�!X�l�.us��Y/k)�ensubL���eK�h�� �B\1;5�g?y?�?�?D��?*r�m�p�?Ktbox  O2K|?�G��C?A%�ds���?�P"�!� �TR��/��P�T6@@�`�U�P�V�P�Ue�P!0�U�PO��\3�U�P �f�Pk"�2}�4�T�P �f�P2�"�Q5�S�Q@���R?Ă�Q3t.�PF׀al��P+O�n�P517��IN0a���Q(}g��PES	Tf3ua�PB�l�i�g�h�6�aq��P �� ,e��` � n�0mbump�P�Q969g�69�Qq��P0�baAp�@>Q� BOX��,�>vche�s�>ve�tu㒣=wffse�3���]�;u`aW��:zol�sm<u�b�a-��]D�K�ib�Q�c����Q<twaǂ �tp�Q҄Taror Recov�br�O�P�642�����a�q��a⁠QErǃ�Qry��`�P'�T�`�aar�������	{'�pak971��71��m���>��`jot��PXc��C��1�adb -�ail���nag���b�QR629�a�Q��b�P�  �
 � �P��$$CL~[q ����������$�PS?_DIGIT���"�!�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v��������*璬1:P�RODUCT�Q0�\PGSTK�bV�,n�99�����$FEAT_INDEX��~~������ILECOM�P ;��)���"��SETUPo2 <��?�  N !��_AP2BCK �1=�  �)}6/E+%,/i/��W/�/~+/�/O/ �/s/�/?�/>?�/b? t??�?'?�?�?]?�? �?O(O�?LO�?pO�? }O�O5O�OYO�O _�O $_�OH_Z_�O~__�_ �_C_�_g_�_�_	o2o �_Vo�_zo�oo�o?o �o�ouo
�o.@�o d�o���M� q���<��`�r� ���%���̏[���� ���!�J�ُn����� ��3�ȟW������"� ��F�X��|����/� ��֯e������0��� T��x������=�ҿ �s�ϗ�,ϻ�9�b�t� P/ 2) *.VRiϳ�!�*���������Ɲ�PC�7�!�F'R6:"�c��χ��T��߽�Lը����x���*.F���>� �	N�,�k�x�ߏ��STM �⠸���Qа���!��iPendant? Panel���H��F���4������GIF�������pu����JPG&�P��<����	�PANEL1.D	T��������2�Y�G��
3w�����//�
4�a/��O///�/�
TP�EINS.XML�/���\�/�/�!�Custom T?oolbar?��PASSWOR�D/�FRS:�\R?? %Pa�ssword Config�?��? k?�?OH�6O�?ZOlO �?�OO�O�OUO�OyO _�O�OD_�Oh_�Oa_ �_-_�_Q_�_�_�_o �_@oRo�_voo�o)o ;o�o_o�o�o�o*�o N�or��7� �m��&���\� ����y���E�ڏi� �����4�ÏX�j��� �����A�S��w�� ���B�џf������� +���O��������� >�ͯ߯t����'��� ο]�򿁿�(Ϸ�L� ۿpς�Ϧ�5���Y� k� ߏ�$߳��Z��� ~�ߢߴ�C���g��� ��2���V����ߌ� ��?����u�
��� .�@���d������)� ��M���q�����< ��5r�%�� [�&�J� n��3�W� ��"/�F/X/�|/ /�/�/A/�/e/�/�/ �/0?�/T?�/M?�?? �?=?�?�?s?O�?,O >O�?bO�?�OO'O�O KO�OoO�O_�O:_�O ^_p_�O�_#_�_�_Y_��_}_o�_�_Ho)f��$FILE_DG�BCK 1=���5`��� ( �)
S�UMMARY.DyGRo�\MD:�o��o
`Diag� Summary��o�Z
CONSLOG�o�o�a
J�a�ConsoleO logK�[�`�MEMCHECK�@'�o�^qMe�mory Dat�a��W�)>�qHADOW����P��sShad�ow Chang�esS�-c-��)	FTP=��9�����w`qmmen�t TBD׏�W0�<�)ETHERNET̏�^�q��Z��aEther�net bpfiguration[���P��DCSVRF�ˏ��Ïܟ�q%��� verify� allߟ-c1P{Y���DIFFԟp��̟a��p%��diffc���q���1X�?�Q�� �����X��CH�GD��¯ԯi��px��� ���2`�G�Y��� ��� �GAD��ʿܿq��p���Ϥ�FY3h�O�aώ�� ��(�GAD������y��p�����0�UPDAT�ES.�Ц��[FORS:\�����a�Updates �List���kPS�RBWLD.CM�.��\��B��_pP�S_ROBOWEL���_����o��,o !�3���W���{�
�t� ��@���d�����/ ��Se����� N�r� =� a�r�&�J� ��/�9/K/�o/ ��/"/�/�/X/�/|/ �/#?�/G?�/k?}?? �?0?�?�?f?�?�?O �?OUO�?yOO�O�O >O�ObO�O	_�O-_�O Q_c_�O�__�_:_�_ �_p_o�_o;o�__o �_�o�o$o�oHo�o�o ~o�o7�o0m�o � ��V�z� !��E��i�{�
��� .�ÏR���������� .�S��w������<� џ`������+���O� ޟH������8���߯�n����$FIL�E_��PR����������� �MDONL�Y 1=4�� 
 ���w�į�� 诨�ѿ�������+� ��O�޿sυ�ϩ�8� ����n�ߒ�'߶�4� ]��ρ�ߥ߷�F��� j�����5���Y�k� �ߏ���B�����x� ���1�C���g���� ��,���P����������?��Lu�VI�SBCKR�<�a��*.VD|�4 OFR:\��4 �Vision VD file�  :LbpZ�# ��Y�}/$/� H/�l/�/�/1/�/ �/�/�/�/ ?�/1?V? �/z?	?�?�???�?c? �?�?�?.O�?ROdOO �OO�O;O�O�OqO_ �O*_<_�O`_�O�__�%_�_�MR_GR�P 1>4�L~�UC4  B�P�	 ]�ol`��*u����RHB ��2 ���� ��� ���He�Y�Q`ork bIh�oJd�o�Sc�o��oMr�J��v&J�F�{5U�aQ�D-�o��o^`��MFU��wD��8���	9 t>�� l}@��@�	�lq?�Ǝ�@~#@��}E�� F@� �r�d�a}J���NJk�H9��Hu��F!�_�IP�s}?�`��.9�<9��896C�'6<,6\�b�}AD��A�l�BN7A�1xA�fA��u� �&�A�P/�B(�@��g�A��VA�K��,.��PA�����|�ݏx����%��  @���A<L�@9�>`�>4��� j�����ǟ���֟���!��E�`r�UBH�P �a`�P��QA[a����Ư�Q�
6�PS@�PS�H}˯�o�oB�x�P5���@�33@����4�m�T�UUU�U�~w�>u.�?!x�^��ֿ����3��=[z��=�̽=V6�<�=�=��=$q~9��@�8�i7G���8�D�8@9!�7ϥ�@Ϣ����cD�@ D�O� Cϫo4z��P��P'�6��_V� m �o��To��xo�ߜo�� ����A�,�e�P�b� ������������ �=�(�a�L���p��� ������.�������* ��N9r]��� �����8# \nY�}���� ���/ԭ//A/� e/P/�/p/�/�/�/�/ �/?�/+??;?a?L? �?p?�?�?�?�?�?�? �?'OOKO6OoO�OH� �Ol��ߐߢ��O�� _ ��G_bOk_V_�_z_�_ �_�_�_�_o�_1oo Uo@oyodovo�o�o�o �o�o�oN u������ ���;�&�_�J��� n�������ݏȏ�� %�7�I�[�"/�描� ����ٟ�������3� �W�B�{�f������� կ�������A�,� e�P�b��������O�O �O��O�OL�_p� :_�����Ϧ������ ��'��7�]�H߁�l� �ߐ��ߴ�������#� �G�2�k�2��Vw� ����������1�� U�@�R���v������� ������-Q� u���r��6� �)M4q\ n������/ �#/I/4/m/X/�/|/ �/�/�/�/�/?ֿ� B?�f?0�BϜ?f��? ���/�?�?�?/OOSO >OwObO�O�O�O�O�O �O�O__=_(_a_L_ ^_�_�_�_���_��o �_o9o$o]oHo�olo �o�o�o�o�o�o�o# G2kV{�h �������C� .�g�y�`��������� �Џ���?�*�c� N���r��������̟ ��)��M�_�&?H? ���?���?�?�?��� �?@�I�4�m�X�j��� ��ǿ���ֿ���� E�0�i�Tύ�xϱϜ� ��������_,��_S� ��w�b߇߭ߘ��߼� ������=�(�:�s� ^��������� �'�9� �]�o���� ~������������� 5 YDV�z� �����1 U@yd��v�� ���/Я*/��
/� u/��/�/�/�/�/�/ �/??;?&?_?J?�? n?�?�?�?�?�?O�? %OOIO4O"�|OBO�O >O�O�O�O�O�O!__ E_0_i_T_�_x_�_�_ �_�_�_o�_/o��?o eowo�oP��oo�o�o �o�o+=$aL �p������ �'��K�6�o�Z�� ����ɏ��폴� � �D�/ /z�D/��h/ ş���ԟ���1�� U�@�R���v�����ӯ ������-��Q�<� u�`���`O�O�O��� ޿��;�&�_�J�o� �πϹϤ�������� %��"�[�F��Fo�� �����ߠo��d�!�� �W�>�{�b���� ����������A�,� >�w�b����������������=��$�FNO ����\��
F0l q  oFLAG>�(R�RM_CHKTY/P  ] ��d ��] ��OM�� _MIN� 	����� �  X�T SSB_CFG� ?\ �����OTP_DEF�_OW  	�|�,IRCOM� �>�$GENOV�RD_DO���<�lTHR� dz�dq_ENB]� qRAVC_?GRP 1@�I X(/ %/7/ /[/B//�/x/�/�/ �/�/�/?�/3??C? i?P?�?t?�?�?�?�? �?OOOAO(OeOLO�^O�OoROU�F\\� �,�|B,�8�?����O�O�O	__��� � DE_�Hy_�\@@m_B�=�vR/��I\�O�SMT�G��SUoo&oRHO7STC�1H�I� ���zMSM��l[bo��	127.0�`1�o  e�o�o�o #z�oFXj|��l60s	anonymous��������%ao�&�&��o�x��o���� ��ҏ�3��,�>� a�O����������Ο �U%�7�I��]���� f�x��������ү� ���+�i�{�P�b�t� ����������� S�(�:�L�^ϭ�oϔ� �ϸ������=��$� 6�H�Zߩ���Ϳs��� �������� �2��� V�h�z��߰����� ����
��k�}ߏߡ� ����߬��������� C�*<Nq�_�� �����-�?�Q� c�eJ��n��� ����/"/E �X/j/|/�/�/� %'/?[0?B?T? f?x?��?�?�?�?�? ?E/W/,O>OPObO�K~DaENT 1I�K� P!�?�O  �P�O�O�O�O�O #_�OG_
_S_._|_�_ d_�_�_�_�_o�_1o �_ogo*o�oNo�oro �o�o�o	�o-�oQ u8n���� ����#��L�q� 4���X���|�ݏ��� ď֏7���[���B�QUICC0��h�z�۟��1ܟ��ʟ�+���2,���{�!ROUTER|��X�j�˯!PCJ�OG̯��!1�92.168.0�.10��}GNAM�E !�J!R�OBOT�vNS_�CFG 1H�I� �Au�to-start{ed�$FTP�/���/�?޿#?�� &�8�JϏ?nπϒϤ� ǿ��[������"�4� �&����������濜� ���������'�9�K� ]�o��������� ����/�/�/G���k� �ߏ������������� 1T���Py� ����"�4�	H -|�Qcu�VD ����/�;/ M/_/q/�/����/ 
/�/>?%?7?I?[? */?�?�?�?�/�?l? �?O!O3OEO�/�/�/ �/�?�O ?�O�O�O_ _�?A_S_e_w_�O4_ ._�_�_�_�_oVOhO zO�O�_so�O�o�o�o �o�o�_'9K no�o�����o *o<oNoP5��oY�k� }�����pŏ׏��� �0���C�U�g�y����_�T_ERR �J;�����PDUS_IZ  ��^P�����>ٕWRD� ?z��� � guest���+�=�O�a�s��*�SCDMNGR�P 2Kz�Ð��۠\���K�� 	P01�.14 8�q �  y��B�    ;�����{ ���߇������������������~ �ǟI�4�m��X�|��  �i  �  
����� ����+��������
����l�.x����"�l�ڲ۰�s�d�������_�GROU��L��� ��	��۠07�K�QUPD  d���PČ�TYg������TTP_AUTH 1M��� <!iPeOndan���<��_�!KARE�L:*�����K�C%�5�G��VI�SION SETZ���|��Ҽߪ� ��������
�W�.��@��d�v���CTRL N��������
�FFF9�E3���FRS�:DEFAULT��FANUC� Web Server�
���� ��q��������������WR_CONFI�G O�� ����IDL_CP�U_PC"��B���= �BH#M�IN.�BGNR_IO��� ���% �NPT_SIM_�DOs}TPM�ODNTOLs >�_PRTY�=�!OLNK 1P���'9K�]o�MASTE�r �����O_CFG��UO����CYCLE���_ASG 1Q���
 q2/D/V/ h/z/�/�/�/�/�/�/��/
??y"NUM����Q�IPC�H��£RTRY�_CN"�u���SGCRN������1 ���R�����?��$J23_�DSP_EN������0OBPROqC�3��JOGV��1S_�@��8G�?�';ZO'??0C�POSREO�KANJI_�ϠuH�A#��3T ���E<�O�ECL_LM B2�e?�@EYLOGG+IN��������LANGUAGE� _�=� ,}Q��LG�2U���+�� �x�����P�C � �'0������MC:\�RSCH\00\�˝LN_DISP V������f�TOC�4Dz\�A�SOGBOOK W+��o���o�o���Xi�o�o�o�o�o~}	x(y��	ne�i�ekEl�G_BUFF 1%X���}2�� ��Ӣ������ '�T�K�]��������� ��ɏۏ���#�P���ËqDCS Z>xm =���%|d�1h`���ʟܟ�g�I�O 1[+ �?'����'�7�I�[� o��������ǯٯ� ���!�3�G�W�i�{�@������ÿ׿�El /TM  ��d��#� 5�G�Y�k�}Ϗϡϳ� ����������1�C߀U�g�yߋߝ߈t�S�EV�0m�TYP�� ��$�}��ARS"�(_�s�2F�L 1\��0� ��������������5�TP<P���>DmNGNAM�4�U��f�UPS`GI�5�A�5s�_LO{AD@G %j{%@_MOV�u�����MAXUALRMB7�P8��y��D�3�0]&q��Ca]s�3�~�� 8@=@]^+ طv	��+V0+�P�A5dƋr���U ������E (iTy���� ���/ /A/,/Q/ w/b/�/~/�/�/�/�/ �/??)?O?:?s?V? �?�?�?�?�?�?�?O 'OOKO.OoOZOlO�O �O�O�O�O�O�O#__ G_2_D_}_`_�_�_�_ �_�_�_�_o
ooUo 8oyodo�o�o�o�o�o��o�o�o-��D_L?DXDISA^��� �MEMO_AP�X�E ?��
 �0y�����������ISCw 1_�� � O����W�i����� Ə�����}��ߏD� /�h�z�a�������� ������@���O� a�5������������ u��ׯ<�'�`�r�Y� �����y�޿�ۿ� ��8Ϲ�G�Y�-ϒ�}� �ϝ�����m�����4���X�j�#�_MST�R `��}�SC/D 1as}�R��� N��������8�#�5� n�Y��}������� �����4��X�C�|� g��������������� 	B-Rxc� ������ >)bM�q�� ���/�(//L/ 7/p/[/m/�/�/�/�/ �/�/?�/"?H?3?l?�W?�?{?�?�?�?n�MKCFG b����?��LTARMu_�2cRuB� �3WpTNBpM�ETPUOp�2�����NDSP_CMNTnE@F�E��' d���N�2A��O�D�EPOSCF��G�NPSTOL� 1e-�4@�<#�
;Q�1;UK_YW 7_Y_[_m_�_�_�_�_ �_�_o�_oQo3oEo��oio{o�o�a�ASI�NG_CHK  y�MAqODAQ2C�fO�7J�eDEV� 	Rz	MC}:'|HSIZEn@�����eTASK �%<z%$123456789 ���u�gTRIG 1]g�� l<u%����3���>svvY�Paq��kEM_I�NF 1h9G� `)AT&FV0E0(����)��E0V1�&A3&B1&D�2&S0&C1S�0=��)ATZ���ڄH������G�ֈAO�w�2�������џ ��������͏ ߏP��t�������]� ί�����(�۟� ^��#�5�����k�ܿ � ϻ�ů6��Z�A� ~ϐ�C���g�y����� ���2�i�C�h�ό� G߰��ߩ��ߙϫ�� ������d�v�)ߚ��� ��y��������<� N��r�%�7�I�[��� ���9�&��J�[�g��>ONIwTOR�@G ?;{�   	EX�EC1�3�2�3��4�5��p�7*�8�9�3�n� R�R�RR RR(R4R@�RLR2Y2e2�q2}2�2�2��2�2�2�3�Y3e3��aR_�GRP_SV 1�it��q(�a�
����fD쿆[��>�\]�w�x@${"}~q_�DCd~�1PL_N�AME !<u�� �!Defa�ult Pers�onality �(from FD�) �4RR2k! �1j)TEX)TsH��!�AX d�? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO@^OpO�O�O�Ox2-? �O�O�O__0_B_T_f_x_�b<�O�_�_�_ �_�_�_o o2oDoVotho&xRj" 1o�)�&0\�b, ��9��b�a @D��  �a?��c�a?x�`�a�aA'�6�e�w;�	l�b	� �xJp��`�`	p� �< ��(p� �.r� K��K ��K=�*�J���J���JV��kq`�q�P�x�|� @j�@T;f�r��f�q�acrs�I�����p����p�r�ph}�3��´  ���>��ph�`z���Ꜭa��3Jm�q� H�N���ac���dw�� ~ �  P� �Q� �� |  �а�m�Əi}	'�� � �I�� �  ��ވ�:�È�È�=���(�ts�a	����I  �n @H�i~�ab�ӋB�b�w��urN0��  'Ж�q�p�@2��@���X�r�q5�C�pC0C�@ C���=�`
�A1q]N� @B�V~�X�
nwB0h�A��p�ӊ�p�`���aDz���֏���Я�	�pv�( �� -��I��0-�=��A�a��e_q��`�p �?�f�f ��m��� ����Ƽuq@tݿ�>1�  P�apv(�`ţ� �=�qxst��?���`�x`�� <
6b<�߈;܍�<��ê<� <G�&P�ό�AO���c1��ƍ�?fff�?O�?&��qt@��.�J<?�`��wi4����dly �e߾g;ߪ�t��p� [ߔ�߸ߣ����� �`���6�wh�F0 %�r�!��߷�1ى�����E�� E�~O�G+� F�!� ��/���?�e�P���t�,��lyBL�cB��E nw4�������+��R ��s�����<����h�Ô�>��I�m0Xj���A�y��weC������Ƀ�#/*/c/N/wi�6����v/C�`� CCHs/`
=$�p�<!��!��ܼ�'�3A��A�AR1A�O�^?�$�?���5p±
=�ç>����3�W
=�#�]�n;e�׬a@�����{����<��>(�B��u��=B�0�������	R��zH�F�G����G��H��U`E���C��+��}I#��I��HD��F��E��R�C�j=�>
�I��@H�!�H�( E<YD0w/O*OONO 9OrO]O�O�O�O�O�O �O�O_�O8_#_\_G_ �_�_}_�_�_�_�_�_ �_"oooXoCo|ogo �o�o�o�o�o�o�o 	B-fQ�u� ������,�� P�b�M���q�����Ώ ���ݏ�(��L�7� p�[������ʟ��� ٟ���6�!�Z�E�W�t��#1($1��9��K���ĥ%�����ƯS�3�8�x��S�4Mgs���,�IB+8�J��a���{�d� d�����ȿ���ڼ%%P8�P�=:G����S�6�h�z���R��Ϯ����������  %�� ��h�Vߌ� z߰�&�g�/9�$�������7����A�8S�e�w�  ��������������2 �F�$�&Gb���������!C���@���8������F� DzN��� F�P D�!������)#B�'�9K]o#?��W�@@v
��8��8��8�.
 v���! 3EWi{�����:� ��ۨ��1��$MSK�CFMAP  ���� ����(.�ONR�EL  ��!9��EXCFE�NBE'
#7%^!F�NCe/W$JOGO/VLIME'dO S"]d�KEYE'�%]�RUN�,�%��SFSPDT�Y0g&P%9#SIG�NE/W$T1MOT��/T!�_CE_�GRP 1p��#\x��?p��?�? �?�?�?O�?OBO �?fOO[O�OSO�O�O �O�O�O_,_�OP__ I_�_=_�_�_�_�_�_�oo�_:o�TC�OM_CFG 1�q	-�vo�o�o
�Va_ARC_b"��p)UAP_CP�L�ot$NOCHE�CK ?	+ �x�%7I [m���������!�.+NO_?WAIT_L 7%6S2NT^ar	+��s�_ERR_129s	)9�� ,ȍޏ��x���&��d�T_MO��t��,� 6�*oq�9�P�ARAM��u	+��a�ß'g{��� =?�345678901��,�� K�]�9�i�������ɯۯ��&g������C��cUM_RSP�ACE/�|����$ODRDSP�c�#6p(OFFSET�_CART�o��D�ISƿ��PEN_FILE尨!�ai���`OPTION_�IO�/��PWOR�K ve7s# ���V�ؤ���p<�p�4�p�	 ����p��<�� C�_DS�BL  ��P#���ϸ�RIENTkTOD ?�C�� �!l�UT_SIM_D$�"����V��LCT w�}�h�iĜa[�1�_P�EXE�j�RAT�vШ&p%� ��2^3j�)TEX)TH�>)�X d3��� ����%�7�I�[�m� ������������ �!�3�E���2��u� ��������������c�<d�ASew ���������Ǎ�^0OUa0o(��(����}u2, ����O H @D�  &[?�aG?��c�c�D][�Z�;��	ls���xJ���������<� ���s��ڐH�(��H3k7H�SM5G�22G���Gp
͜��'f�/-,ڐC%R�>�D!�M#{|Z/��3�����4y H "�c/u/��/0B_���{�jc��t�!�/ �/�"t32�����/6  ���P%�Q%��%�|�T��S62�q?'e	'�� � �2I�� �  �=�+==��ͳ?�;�	�h	�0�I  ?�n @�2�.��Ov;��ٟ?&g9N�]O  ''�uDt@!� C�C�@F#�H!�/�O�O sb
����@�@�H�@�e0@B�QA�0Yv: �13Uwz$oV_�/z_e_�_�_�	��( �� -�2�1�1ta��Ua�c���:A�����.  �?�ff ���[o"o�_U�`oDX�0A8���o�j>�1'  Po�V(���e�F0�f�Y���L�?�����xb0@<�
6b<߈;�܍�<�ê<� <�&�,/aA�;r�@Ov0P�?fff?�0?&�ip�T@�.{r�?J<?�`�u#	 �Bdqt�Yc�a� Mw�Bo��7�"�[� F��j�������ُ� ���3����,����(�E�� E�~�3G+� F��a ��ҟ�����,��PP�;���B�pAZ� >��B��6�<OίD��� P��t�=���a�s���<��6j�h��7o��>�S��O��0���Fϑ�A�a�_���C3Ϙ�/�%?��?���������#	�Ę��P �N||CH���Ŀ�������@I�_�'�3�A�A�AR1�AO�^?�$��?�����±
�=ç>�����3�W
=�#�\ U��e���B��@���{����<����(�B��u��=B�0�������	�b�H�F�G����G��H��U`E���C��+��I#��I��HD��F��E��R�C�j=[�
�I��@H�!�H�( E<YD0߻������ ��� �9�$�]�H�Z� ��~������������� #5 YD}h� ������
 C.gR���� ���	/�-//*/ c/N/�/r/�/�/�/�/ �/?�/)??M?8?q? \?�?�?�?�?�?�?�? O�?7O"O[OmOXO�O |O�O�O�O�O�O�O�Ot3_Q(�������b��gUU���W_i_2�3�8�x�_�_2�4Mgs�_��_�RIB+�_�_�a���{�m iGo5okoYo�o}l��%P'rP�nܡݯ�o�=_�o�_�[R�?Q�u���  �p���o��/� �S��z
uүܠ�������ڱ�������8����  /�M��w�e��������l2 �F�$��Gb���t��a�`�p�S�C�y�@p�5�G�Y�۠�F� Dz��� F�P D�!�]����پ��ʯ�ܯ� ��~�?��W�@@�?�K��K���K���
 �|�������Ŀ ֿ�����0�B�TϸfϽ�V� ���{���1��$PAR�AM_MENU �?3���  DE�FPULSEr��	WAITTMO{UT��RCV��� SHELL�_WRK.$CU�R_STYL���	�OPT��P�TB4�.�C�R_DECSN���e�� ߑߣ���������� �!�3�\�W�i�{�����USE_PRO/G %��%����.��CCR���e�����_HOST �!��!��:���T �`�V��/�X��>��_TIME��^���  ��GDE�BUG\�˴�GI�NP_FLMSKĻ���Tfp����PG�A  ����)CyH����TYPE��������� �� -?hc u������� //@/;/M/_/�/�/ �/�/�/�/�/�/??�%?7?`?��WORD� ?	=	R}Sfu	PNSU�Ԝ2JOK�DR�TEy�]TRACECTL 1x3���� �`X/ &�`�`�>��6DT Qy3��%@�0D � ޱc�a0:@V�@BR�2ODOVOhOzO�B�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo*x`|d�b�h�o �g�m�amj�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�.Iv� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��j� ���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�o�o�o�o ��o0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�L�^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ����������*��$PGTR�ACELEN  �)�  ���(��>�_U�P z���2m�u�Y�n�>�_CFG {m�SW�(�n����PКӂ�DEFSP/D |��'�P���>�IN��TR�L }��(�8�����PE_CON�FI��~m���mњ��ղ�L�ID����=�G�RP 1��W���)�A ����&ff(�A+33�D�� D]� ?CÀ A@1����(�d�Ԭ��0�0�?� 	 1��8�֚��� ´�����B�9����O��9�s�(�>�T?��
5�������� �=��=#�
 ����P;t_�������� G Dz (�
 H�X~i��� ���/�/D///�h/S/�/��
V7�.10beta1���  A��E�"ӻ�A �(�� ?!G��!>����"����!{���!BQ��!�A\� �!���!2p
����Ț/8?J?\?�n?};� ���/� �/�?}/�?�?OO:O %O7OpO[O�OO�O�O �O�O�O_�O6_!_Z_ E_~_i_�_�_�_�_�_ �_'o2o�_VoAoSo �owo�o�o�o�o�o�o .R=v1�/�#F@ �y�}� �{m��y=��1�'� O�a��?�?�?������ ߏʏ��'��K�6� H���l�����ɟ��� ؟�#��G�2�k�V� ��z��������o� �ίC�.�g�R�d��� �������п	���-� ?�*�cώ���Ϯ� �����B�;�f� x�������DϹ��߶� �������7�"�[�F� X��|��������� ��!�3��W�B�{�f� �������� ����� /S>wbt� �����= OzόϾψ����� �� /.�'/R�d�v� �߁/0�/�/�/�/�/ �/�/#??G?2?k?V? h?�?�?�?�?�?�?O �?1OCO.OgORO�OvO �O�O���O�O�O__ ?_*_c_N_�_r_�_�_ �_�_�_o�_)oTf x�to���/�o />/P/b/t/m o�|����� ��3��W�B�{�f� x�����Տ������ �A�S�>�w�b����O ��џ������+�� O�:�s�^�������ͯ ���ܯ�@oRodo�o `��o�o�o��ƿ�o� ��*<N�Y��}� hϡό��ϰ������� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�c�N�ﲟ��� l��������;�&� _�J���n��������� ��,�>�P�:L�� ���������� (�:�3��0iT� x�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?a?s?��?�?X?�? �?�?�?O'OOKO6O oOZO�O~O�O�O�O�O *\&_8_r����_�_��$PLI�D_KNOW_M�  ��� Q�TSV ���P��?o"o4o�OXo�CoUo�o R�SM_?GRP 1��Z'U0{`�@�`uf
�e�`
�5� �gpk 'Pe] o�������X���SMR�c��m1T�EyQ}? yR�� ��������폯���ӏ �G�!��-������� ����韫���ϟ�C� ��)������������寧���QST�a1W 1��)���P;0� A 4��E 2�D�V�h�������߿ ¿Կ���9��.�o� R�d�vψ��ϬϾ�����2�0� Q�	<3��3�/�A�S߂�4l�~ߐߢ��5 ���������6
��.�@��7Y�k�}���8��������M_AD  )���PARNUM  !�}o+��WSCHE� S�
��pf���S��UPDf��x��_CM�P_�`H�� �'��UER_CHK-���ZE*<�RSr��_�Q_MO�G���_�X�_R/ES_G��!��� D�>1bU� y�����/�	/����+/� k�H/g/l/��Ї/�/ �/�	��/�/�/�X� ?$?)?���D?c?h?�����?�?�?�V �1��U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_�INRr�J�b�Ud�2FMASS?O Z�SGMN>OqCMON�_QUEUE a��U�V P~P X�N$ UhN�FV�@�END�A��IEX1E�O�E��BE�@�O>�COPTIO�G���@PROGRAM7 %�J%�@�?����BTASK_I�G�6^OCFG ኤOz��_�PDATuA�c��[@Ц2=�DoVohozo�j2o �o�o�o�o�o)x;M jINFO[��m��D��� �����1�C�U� g�y���������ӏ����	�dwpt�l �)�QE DIT ��_i��^WERF�LX	C�RGADoJ �tZA���¿�?נʕFA��IOORITY�GW���MPDSPNQ�����U�GD��OTO�E@1�X� (/!AF:@E� c�~Ч!tcpn�>��!ud����!icm���?<��XY_�Q�X�=��Q)� *�1�5��P��]�@�L� ��p��������ʿ� �+�=�$�a�Hυϗ�=*��PORT)QH���P�E��_C?ARTREPPX�>�SKSTA�H�
�SSAV�@�tZ	�2500H86A3���_x�
�'��X�@�swPtS��x�ߧ���URGE�@�B��x	WF��DO�F"[W\��������WRUP_DEL�AY �X���RO_HOTqX	B%��c���R_NORM�ALq^R��v�SE�MI�����9�QS�KIP'��tUr�x 	7�1�1�� X�j�|�?�tU������ ��������$J \n4����� ���4FX |j������ �/0/B//R/x/f/�/�/�/tU�$RCgVTM$��D�� �DCR'����ގ!@Y�1�C
�ց>�<>� 7��B:��ZR�Dܠ��c|���H�}?��<
6�b<߈;܍��>u.�?!<�&Y?g?�?�? �A-2�?O!O3OEOWO iO{O�O�O�O�O�O�? �O�O__A_,_Q_w_ Z_�_�_�?�_�_�_o o+o=oOoaoso�o�o �_�_�o�o�o�o  9K.o��_�� �����#�5�G� Y�k�V��z���ŏ�� �ԏ���C��� y���������ӟ��� 	��-�?�*�c�N��� r��������į�� Z�;�M�_�q������� ��˿ݿ�����7� "�[�F��j�|ϵϘ� ����.��!�3�E�W� i�{ߍߟ߱������� �����/��S�>�w� ��l��������� �+�=�O�a�s����� �����������' K]@���� ����#5G�Yk}��!GN_�ATC 1�	;� AT&F�V0E0�A�TDP/6/9/�2/9�ATA��,AT%G1%B960�_+++�,��H/,�!IO_T?YPE  �%�#�t�REFPO�S1 1�V+ 'x�u/�n�/ j�/
=�/�/�/Q?<? u??�?4?�?X?�?�?^�+2 1�V+�/��?�?\O�?�O�?�!3 1�O*O<OvO�O��O_�OS4 1� �O�O�O_�_t_�_+_S5 1�B_T_f_�_o	oBo�_S6 1��_�_�_5o�o�o|�oUoS7 1�lo�~o�o�oH3l�oS8 1�%_����SMAS�K 1�V/  
8?�M��XNOS/�r�������!MOT�E  n��$��_CFG ����q����"PL_RANG������POWER� �����S�M_DRYPRG %o�%�P��TART ���^�UME_PRO�-�?����$_EXE�C_ENB  <���GSPD��Ր8ݘ��TDB��
�sRM�
�MT_'��T����OBO�T_NAME �o����OB_�ORD_NUM �?�b!H863  ��կ���PC�_TIMEOUT��� x�S232�Ă1�� L�TEACH PENDAN��w���-��Ma�intenanc?e Cons����s�"���KCLC/Cm��

���t��ҿ No U�se-��Ϝ�0�N�PO�򁋁z��.�CH_L��3����q	��s�?MAVAIL����糅��SPAC�E1 2��, j�߂�D��s�߂�� �{S�8�?�k�v�k�Z߬��� ���ߚ� �2�D��� hߊ�|��`������ ����� �2�D�� h��|���`�������(��y���2���� 0�B���f�����{ ���3) ;M_����@��/� /44 FXj|*/���/��/�/?(??=?5 Q/c/u/�/�/G?�/�/ �?O�?$OEO,OZO6n?�?�?�?�?dO�? �?_,_�OA_b_I_w_7�O�O�O�O�O�_ �O_(oIoo^oofo�o8�_�_�_�_�_ �oo6oEf){�x��G �o�� ���
M� ���*�<�N�`� r�������w���o�収���d.��%� S�e�w����������� Ǐَ���Θ8�+�=� k�}�������ůׯ͟ ����%�'�X�K�]� ��������ӿ�������#�E�W� `� @�������x�����\�e����� ������R�d߂�8� j߬߾߈ߒߤ���� ������0�r���X� ������������8�����
�ύ�_M?ODE  �{��/S ��{|�2ς0�����3�	�S|)CWORK�_AD��	��^+R  �{�`�� �� _INTV�AL���d���R_�OPTION� ���H VAT_�GRP 2��u;p(N�k|��_� ����/0/B/�� h�u/T� }/�/�/�/ �/�/�/?!?�/E?W? i?{?�?�?5?�?�?�? �?�?O/OAOOeOwO �O�O�O�OUO�O�O_ _�O=_O_a_s_5_�_ �_�_�_�_�_�_o'o 9o�_Iooo�o�oUo�o �o�o�o�o�o5G Yk-���u� ����1�C��g� y���M�����ӏ叧� 	��-�?�Q�c����� ����������ǟ��;�M�_����$SCAN_TIM���_%}�R ��(�#((�<0�4d d 
!D�ʣ���u�/�����U��25���@��d5�P�g��]	 ���������dd�x��  P����; ��  8� ҿx�!���D��$� M�_�qσϕϧϹ���������ƿv���F�X��/� ;G�ob��pm���t�_Di�Q̡  � l �|�̡ĥ������� !�3�E�W�i�{��� ������������/� A�S�e�]�Ӈ����� ��������); M_q����� ��r���j�T fx������ �//,/>/P/b/t/��/�/�/�/�/�%�/  0��6��!?3?E? W?i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O*�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo�O�OJ�o�o �o�o�o�o�o 2 DVhz��������
�7?   ;�>�P�b�t������� ��Ǐُ����!�3� E�W�i�{�������ß �ş3�ܟ�� &�8�J�\�n�������������ɯ�����,� �+�	�1234567�8�� 	� =5���f�x�������������
��.� @�R�d�vψϚ�៾� ��������*�<�N� `�r߄߳Ϩߺ����� ����&�8�J�\�n� �ߒ����������� �"�4�F�u�j�|��� ������������ 0_�Tfx��� ����I> Pbt����� ��!/(/:/L/^/ p/�/�/�/�/�/�/�2�/?�#/9?K?�]?�iCz  B}p˚   ��h�2��*�$SCR�_GRP 1�(��U8(�\x�d�@} � ��'�	 �3�1�2�4(1*�&��I3�F1OOXO}m��D�@�0ʛ�)���HUK�LM�-10iA 89�0?�90;��F;�M61C D�:�CTP��1
\&V�1 	�6F��CW�9)A7Y	(R�_�_�_�_�_�\���0i^�o OUO>oPo#G�/����o'o�o�o�o�oB��0�rtAA�0*  @�Bu&"Xw?��ju�bH0{�UzAF@ F�`�r��o���� �+��O�:�s��mBq�rr����������B� ͏b����7�"�[�F� X���|�����ٟğ�� �N���AO�0�B�CU�
L���E�jqBq>73����$G@�@pϯ7 B���G�I�
E�0EL_DEFAULT  �T���E���MIPOWERFL  
E*���7�WFDO� �*��1ERVENT? 1���`(��� L!DUM�_EIP��>��j�!AF_INEx�¿C�!FT�������!o:� ���a�!RP?C_MAINb�D�q�Pϭ�t�VIS}��Cɻ����!TP&��PU�ϫ�d��E��!
PMON_POROXYF߮�e4ߐ���_ߧ�f����!�RDM_SRV��߫�g��)�!R��Iﰴh�u�!
�v�M�ߨ�id���!RLSYNC���>�8���!R3OS��4��4��Y� (�}���J�\������� ������7��[" 4F�j|�����!�Eio�I�CE_KL ?%�� (%SVCPRG1n>����3��3���4�//�5./3/�6V/[/�7~/�/��D$�/�9�/�+�@� �/��#?��K?� �s?� /�?�H/�? �p/�?��/O��/ ;O��/cO�?�O� 9?�O�a?�O��?_ ��?+_��?S_�O {_�)O�_�QO�_� yO�_��Os��� �>o�o}1�o�o�o�o �o�o�o;M8 q\������ ���7�"�[�F�� j�������ُď��� !��E�0�W�{�f��� ��ß���ҟ��� A�,�e�P���t�����࿯�ί�y_DE�V ���MC:���_.!�OUT��2�~�REC 1�`e��j� �� 	 ������������ѽ��ſۿ��
 ��PSD#6 �r  ��O����  �  `D��>��`e�����E���0�R��+^ͪ3���I3��3�!
3����^Ͽ�_��� h��� ���$��H�6� l�~�`ߢߐ��ߴ��� ���� ���V�D�z� h������������ �
��R�@�v���j� ������������* N<^�r�� ����&J 8Z�b���� ���"/4//X/F/ |/j/�/�/�/�/��2� �/�/�/?:?(?^?L? �?�?v?�?�?�?�?�? �? O6OOFOlOZO�O ~O�O�O�O�O�O_�O 2_ _B_h_V_�_n_�_ �_�_�_�_
o�_.o@o "odoRotovo�o�o�o �o�o�o<*` Np�x���� ���8�J�,�n�\� ��������Ə�Ώ�� ���F�4�j�X���`��p�V 1�}� P亸����� ?n7 1����TYPE\��HE�LL_CFG �.�є��?�r�����RSR������ ӯ�������?�*� <�u�`���������Ῥ���N��%@�3�E��Q�\���1M�o�p������2��d]�K�:�HKw 1�H� u� ������A�<�N�`� �߄ߖߨ������������&�8��=�OM�M �H���9�FTOV_ENB&��1�OW_REG�_UI��8�IMW�AIT��a���O�UT������TI�M�����VA�L����_UNIT���K�1�MON_ALIAS ?ew�? ( he���� ��������ж��) ;M��q���� d��%�I [m�<��� ���!/3/E/W// {/�/�/�/�/n/�/�/ ??/?�/S?e?w?�? �?F?�?�?�?�?�?O +O=OOOaOO�O�O�O �O�OxO�O__'_9_ �O]_o_�_�_>_�_�_ �_�_�_�_#o5oGoYo koo�o�o�o�o�o�o �o1C�ogy ��H����	� �-�?�Q�c�u� ��� ����ϏᏌ���)� ;��L�q�������R� ˟ݟ�����7�I� [�m��*�����ǯٯ 믖��!�3�E��i� {�������\�տ��� ��ȿA�S�e�wω� 4ϭϿ����ώ���� +�=�O���s߅ߗߩ� ��f�������'��� K�]�o���>���� ������#�5�G�Y���}���������n���$SMON_DE�FPRO ������� *SYST�EM*  d=���RECALL �?}�� ( �}��>Pbt�� ,���� �;M_q��( ����//�7/ I/[/m//�/$/�/�/ �/�/�/?�/3?E?W? i?{?�? ?�?�?�?�? �?O�?/OAOSOeOwO �OO�O�O�O�O�O_ _�O=_O_a_s_�_�_ *_�_�_�_�_oo�_ 9oKo]ooo�o�o&o�o �o�o�o�o�o5G�Yk}�"x&co�py mc:di�ocfgsv.i�o md:=>i�nspiron:3648���	��~0�rfrs:o�rderfil.�dat virt:\temp\��`�r�����)q(.�*.dB�T�W������{
xyzrate 61 ��ˏݏn�����%u.�O�H� Z�����"x3.�@�?mpbackN�b��t����� }*�sdb��*C�U�Y����l�!y.x.�:\���8�R�ݯn�����%u/.�a6�H�_�^��� �&�8���ܯm�ϑ� ����ȯZ������"� 4�ǿX�i�{ߍߠ��� C�ֿ������0�B� T�e�w��Ϯ�I��� ������,߿�P�a� s�������;���`��� (�������n�������6044  HZ��"�4�� �as����E� Y��/!�3�F� �n/�/�/��6/H/�  ^/�/??&8�� m??�?���Z?�?��?O!7�$SNP�X_ASG 1�����9A�� P 0 �'%R[1]�@1.1O 9?�#3%dO�OsO�O�O�O �O�O�O __D_'_9_ z_]_�_�_�_�_�_�_ 
o�_o@o#odoGoYo �o}o�o�o�o�o�o�o *4`C�gy �������	� J�-�T���c������� ڏ�����4��)� j�M�t�����ğ���� ��ݟ�0��T�7�I� ��m��������ǯٯ ���$�P�3�t�W�i� �������ÿ���� :��D�p�Sϔ�wω� �ϭ��� ���$��� Z�=�dߐ�sߴߗߩ� ������ ��D�'�9� z�]��������� 
����@�#�d�G�Y� ��}������������� *4`C�gy ������	 J-T�c��� ���/�4//)/ j/M/t/�/�/�/�/�/��/�/?0?4,DPA�RAM �9E}CA �	��:�P�4�0$HOF�T_KB_CFG�  p3?E�4PI�N_SIM  9K�6�?�?�?�0,@�RVQSTP_DSB�>�21On8J0�SR ��;� ?& CAR=O~N��6TOP_O/N_ERl@�F�8~�APTN �5��@A�BRING_PRM�O� J0VDT_G�RP 1�Y9�@  	�7n8_(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2Dkhz �������
� 1�.�@�R�d�v����� ����Џ�����*� <�N�`�r��������� ̟ޟ���&�8�J� \�����������ȯگ ����"�I�F�X�j� |�������Ŀֿ�� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�tߛߘߪ� ����������(�:� a�^�p������� ���� �'�$�6�H�Z� l�~���������������3VPRG_CO7UNT�6��A�5NENB�OM=��4J_UPD 1}��;8  
 p2������  )$6Hql~� ����/�/ / I/D/V/h/�/�/�/�/ �/�/�/�/!??.?@? i?d?v?�?�?�?�?�? �?�?OOAO<ONO`O �O�O�O�O�O�O�O�O __&_8_a_\_n_�_��_�_YSDEBSUG" � �Pdk	��PSP_PASS�"B?�[LOG� ��mr�P�X�_  �g~�Q
MC:\d<�_b_MPCm�H�o�o�Qa�o �~vfSAV �m�:dUb�U\gS�V�\TEM_TI�ME 1�� �(�P��T��o	T1SVGUNS} �#'k�spAS�K_OPTION�" �gospBC?CFG ��|� �b�{�}` ����a&��#�\�G� ��k�����ȏ����� �"��F�1�j�U��� y���ğ���ӟ��� 0��T�f��UR��� S���ƯA������ � �D��nd��t9�l��� ������ڿȿ���� �"�X�F�|�jϠώ� �ϲ���������B� 0�f�T�v�xߊ��ߦ� ��������(��L� :�\��p������ ����� �6�$�F�H� Z���~����������� ��2 VDzh ������� ��4Fdv�� ����//*/� N/</r/`/�/�/�/�/ �/�/�/??8?&?\? J?l?�?�?�?�?�?�? �?�?OO"OXOFO|O 2�O�O�O�O�OfO_ �O_B_0_f_x_�_X_ �_�_�_�_�_�_oo oPo>otobo�o�o�o �o�o�o�o:( ^Lnp���� �O��$�6�H��l� Z�|�����Ə؏ꏸ� ���2� �V�D�f�h� z�����ԟ���� 
�,�R�@�v�d����� ����ίЯ���<� �T�f�������&�̿ ��ܿ��&�8�J�� n�\ϒπ϶Ϥ����� �����4�"�X�F�|� jߌ߲ߠ��������� ��.�0�B�x�f�� R������������,� �<�b�P�������x� ��������&( :p^����� �� 6$ZH ~l������ ��/&/D/V/h/��/�z/�/�/�/�/�&0��$TBCSG_G�RP 2��%�  �1� 
 ?�   /?A?+?e?O?�?s?�?@�?�?�?�;23�<�d, �$A?~1	 HC���6�>��@E�5CL  B�'2^OjH4Jw��B\)LF�Y  A�jO�MB��?�IBl�O�O�@��JG_�@�  DA	�15_ __$YC-P�{_F_`_j\��_�]@ 0�>�X�Uo�_�_6o�Soo0o~o�o�k�h��0	V3.0�0'2	m61c�c	*�`�d2�o&�e>�JC0(�a�i� ,p�m-  �0����omvu1JCFG ��%� 1 #0vz�ʠrBrv�x����z� �%�� I�4�m�X���|����� ���֏���3��W� B�g���x�����՟�� ������S�>�w� b�����'2A ��ʯܯ ������E�0�i�T� ��x���ÿտ翢�� ��/��?�e�1�/�� �/�ϜϮ�������� ,��P�>�`߆�tߪ� ���߼�������� L�:�p�^����� ������� �6�H�>/ `�r������������ ���� 0Vhz 8������
 .�R@vd� ������// </*/L/r/`/�/�/�/ �/�/�/�/�/?8?&? \?J?�?n?�?�?�?�? ���?OO�?FO4OVO XOjO�O�O�O�O�O�O __�OB_0_f_T_v_ �_�_�_z_�_�_�_o o>o,oboPoroto�o �o�o�o�o�o( 8^L�p��� ����$��H�6� l�~�(O����f�d�� ؏���2� �B�D�V� ������n����ԟ
� ��.�@�R�d����v� �������Я���*� �N�<�^�`�r����� ̿���޿��$�J� 8�n�\ϒπ϶Ϥ��� ����ߊ�(�:�L��� |�jߌ߲ߠ������� ���0�B�T��x�f� ������������� ,��P�>�t�b����� ����������: (JL^���� �� �6$Z H~l��^��� dߚ //D/2/h/V/ x/�/�/�/�/�/�/�/ ?
?@?.?d?v?�?�? T?�?�?�?�?�?OO <O*O`ONO�OrO�O�O �O�O�O_�O&__6_ 8_J_�_n_�_�_�_�_ �_�_�_"ooFo�� po�o,oZo�o�o�o�o �o0Tfx� H������� ,�>��b�P���t��� ������Ώ��(�� L�:�p�^�������ʟ ���ܟ� �"�$�6� l�Z���~�����د� �o��&�ЯV�D�z� h�������Կ¿��
� �.��R�@�v�dϚ�΄�  ���� ��������$TB�JOP_GRP �2ǌ��?  ?������������xJBЌ���9� �<� �X���� �@���	 �C��� t�b  C�x���>��͘�̐դ�>̚йѳ33=�CLj��fff?��?�ffBG��ь�����t޽ц�>�(��\)�ߖ�E噙��;��hCYj���  @h��B� � A����f��C�  Dhъ�1����O�4�N�����
:���Bl^��j�i�l�l����?Aə�A�"��sD��֊=qH����нp�h�Q�;�A�j��ٙ�@L��D	�2�������$�6�>BÏ\��T���Q�ts}x�@33@���C���y�1����>��Dh�����������<{�h�@i� �� t��	���K &�j�n|�� �p�/�/:/k/��ԇ���!��	�V3.00J�m761cI�*� I�����/�' Eo��E��E���E�F���F!�F8���FT�Fq�e\F�NaF����F�^lF����F�:
F���)F��3G��G��G���G,I�!C�H`�C�dTD�U�?D��D���DE(!/E�\�E��E��h�E�ME���sF`F�+'\FD��F�`=F}'�F���F�[
F����F��M;^��;Q�T,8�4E` *�ϴ?�2����3\�X/O��ES�TPARS  ظ�	���HR@AB_LE 1����0��
H�7 8��9
G�
H
H����
G	�
H

H
HYE���
H
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_ P_b_t_�^:BS _� �JGoYoko}o�o�o �o�o�o�o�o1 CUgy����` #oRL�y�_�_�_�_�O��O�O�O�OX:B�rN�UM  ��*�P��� V@P�:B_CFG �譋Z�h�@��IMEBF_TT%AU��2@�VERS�q���R 1���
' (�/����b� ����J�\���j�|� ��ǟ��ȟ֟���� �0�B�T���x��������2�_���@�
���MI_CHAN��� � ��DBGLV����������ETHERAD �?��O���ಯ��h�����ROUmT�!��!�������SNMASK�D��U�255.����#�����OOL�OFS_DI%@��u.�ORQCTRL �����}ϛ3 rϧϹ��������� %�7�I�[�:���h�z����APE_DET�AI"�G�PON_�SVOFF=���P_MON �֍��2��STRTC_HK �^������VTCOMPA�T��O�����FPR�OG %^�%�CA�����ISP�LAY&H��_IN�ST_Mް �������US�q��L�CK���QUIC�KME�=���SC�REZ�G�tps� ���u�z�����_��@@n�.�S�R_GRP 1о^� �O� ���
��+O=sa�쀚�
m�� ����L/C 1gU�y��� ��	/�-//Q/?/�a/�/	1234�567�0�/�/@X�t�1���
 �}�ipnl/� g?en.htm�?� ?2?D?V?`P�anel setupZ<}P�?�?�?�?�?�? �??,O >OPObOtO�O�?�O!O �O�O�O__(_�O�O ^_p_�_�_�_�_/_]_ S_ oo$o6oHoZo�_ ~o�_�o�o�o�o�o�o so�o2DVhz� 1'���
�� .��R��v��������ЏG���UALR�M��G ?9� �1�#�5�f�Y��� }�������џן����,��P��SEV � ����E?CFG ������A��   BȽ�
 Q���^� ���	��-�?�Q�c�@u�������������C �����I��?���(%D�6� � $�]�Hρ�lϥϐ��� ��������#��G����� �߿U�I_�Y�HIST 1վ�  ("�� ��(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1����(�f:�'����71�߀�����J���`�ewdit��CARt� 
��.�@�K�=�g�y� ��������P�����	 -?��cu�� ��L^�) ;M�q�������f��f// '/9/K/]/`�/�/�/ �/�/�/j/�/?#?5? G?Y?�/�/�?�?�?�? �?�?x?OO1OCOUO gO�?�O�O�O�O�O�O tO�O_-_?_Q_c_u_ _�_�_�_�_�_�_� �)o;oMo_oqo�o�_ �o�o�o�o�o�o% 7I[m� � ������3�E� W�i�{������ÏՏ �������A�S�e� w�����*���џ��� ��ooO�a�s��� ������ͯ߯��� '���K�]�o������� ��F�ۿ����#�5� ĿY�k�}Ϗϡϳ�B� ��������1�C��� g�yߋߝ߯���P��� ��	��-�?�*�<�u� ������������ �)�;�M�������� ��������l�% 7I[����� ��hz!3E Wi������ �v////A/S/e/�P���$UI_P�ANEDATA �1�����!�  	�}w/�/�/�/�/?? )?>?V�/i?{? �?�?�?�?*?�?�?O OOAO(OeOLO�O�O �O�O�O�O�O�O_&Y� b�>RQ?V_ h_z_�_�_�__�_G? �_
oo.o@oRodo�_ �ooo�o�o�o�o�o �o*<#`G��}�-\�v�#�_� �!�3�E�W��{��_ ����ÏՏ���`�� /��S�:�w���p��� ��џ������+�� O�a���������ͯ ߯�D����9�K�]� o��������ɿ��� Կ�#�
�G�.�k�}� dϡψ����Ͼ���n� ��1�C�U�g�yߋ��� ����4�����	��-� ?��c�J����� �����������;�M� 4�q�X��������� ��%7��[�� �����@� �3WiP� t�����/� //A/����w/�/�/�/ �/�/$/�/h?+?=? O?a?s?�?�/�?�?�? �?�?O�?'OOKO]O DO�OhO�O�O�O�ON/ `/_#_5_G_Y_k_�O �_�_?�_�_�_�_o o�_Co*ogoyo`o�o �o�o�o�o�o�o-�Q8u�O�O}���������) �>��U-�j�|����� ��ď+��Ϗ��� B�)�f�M��������� �����ݟ��XS�K��$UI_PAN�ELINK 1��U  ��  ��}�1234567890s���������ͯ դ�Rq����!�3�E� W��{�������ÿտDm�m�&����Qo�  �0�B�T�f�x� �v�&ϲ��������� ߤ�0�B�T�f�xߊ� "ߘ����������� ��>�P�b�t���0� ������������$� L�^�p�����,�>�������� $�0, &�[�XI�m�� �����>P 3t�i��Ϻ � -n��'/9/K/]/ o/�/t�/�/�/�/�/ �/?�/)?;?M?_?q? �?�UQ�=�2"��? �?�?OO%O7O��OO aOsO�O�O�O�OJO�O �O__'_9_�O]_o_ �_�_�_�_F_�_�_�_ o#o5oGo�_ko}o�o �o�o�oTo�o�o 1C�ogy��� ��B�	��-�� Q�c�F�����|����� ��֏�)��M�� �=�?��?/ȟڟ� ���"�?F�X�j�|� ����/�į֯���� �0��?�?�?x����� ����ҿY����,� >�P�b��ϘϪϼ� ����o���(�:�L� ^��ςߔߦ߸����� ��}��$�6�H�Z�l� �ߐ���������y� � �2�D�V�h�z�� ��-���������
�� .RdG��} ����c���< ��`r����� ���//&/8/J/� n/�/�/�/�/�/7�I� [�	�"?4?F?X?j?|? ��?�?�?�?�?�?�? O0OBOTOfOxO�OO �O�O�O�O�O_�O,_ >_P_b_t_�__�_�_ �_�_�_oo�_:oLo ^opo�o�o#o�o�o�o �o ��6H�l ~a������ ��2��V�h�K��� ����1�U
�� .�@�R�d�W/������ ��П������*�<� N�`�r��/�/?��̯ ޯ���&���J�\� n�������3�ȿڿ� ���"ϱ�F�X�j�|� �Ϡϲ�A�������� �0߿�T�f�xߊߜ� ��=���������,� >���b�t����� +������:�L� /�p���e��������� �� ��6����ۏ��$UI_Q�UICKMEN � ����}��RESTO�RE 1٩��  � 
�8m3\ n���G��� �/�4/F/X/j/|/ '�/�/�//�/�/? ?0?�/T?f?x?�?�? �?Q?�?�?�?OO�/ 'O9OKO�?�O�O�O�O �OqO�O__(_:_�O ^_p_�_�_�_QO[_�_ �_I_�_$o6oHoZolo o�o�o�o�o�o{o�o  2D�_Qcu �o������� .�@�R�d�v�������Џ⏜SCRE�� ?�uw1sc� u2�U3�4�5�6��7�8��USE�R����T���k�s'���4��5��6ʆ�7��8��� ND�O_CFG ڶ�  �  � P�DATE h��None��SEUFRAME�  ϖ��R�TOL_ABRT8����ENB(��?GRP 1��	�Cz  A�~� |�%|�������į֦!��X�� UH�X�~7�MSK  K�4S�7�N�%uT��%�����VISCAND_MAXI��I�3���FAI�L_IMGI�z ��% #S���IMRE/GNUMI�
���gSIZI�� �ϔ�,�ONTMOiU'�K�Ε�&�����a��a���s�FR:�\�� � �MC:\(�\LO�Gh�B@Ԕ !�{��Ϡ�����z? MCV����oUD1 �EX	��z ��PO64�_�Q��n66��PO!�LI�O�䞶e�V�N�f@�`�I�� =	_�S�ZVmޘ��`�W�AImߠ�STAT' �k�% @��4�F�T�$#�x �2�DWP  ���P G��=���͎���_JMPERR 1ޱ�
  �p2345?678901�� �	�:�-�?�]�c��� ��������������$�MLOW�ޘ���Ό�_TI/�˘'���MPHASE � k�ԓ� ��SoHIFT%�1 Ǚ��<z��_ ����F/ |Se����� ��0///?/x/O/ a/�/�/�/�/�/�����k�	VSFT]1[�	V��M+3� �5�Ք p��~��A�  B8[0[0�Πpg3a1Y21�_3Y�7ME��K��͗	6e���&%�J�M���b��	���$��TDINE#ND3�4��4OH�+�G1�OS2OIV I����]LRELE�vI��4.�@��1_ACTIV�IT��B��A �m��/_���BRDBГOZ�YBOX �ǝf_[��b�2�TI190.0.�P�83p\�V25�4p^�Ԓ	 ��S�_�[b���robot84q_ ?  p�9o[�pc�PZoMh��]Hm�_Jk@1�o�ZWABCd��k�,�� �P[�Xo}�o0) ;M�q����@����>��aZ�b��_V