��  ���A��*SYST�EM*��V7.5�0130 3/�19/2015 AM  �����ABSPOS�_GRP_T �   $PA�RAM  �(�ALRM_RECOV1�   $AL]MOENB��]�ONi�APCO�UPLED1 �$[PP_PRO�CES0  ��1�"  |U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $� �� NO�PS_SPI_INDE���$�X�SCR�EEN_NAME� �SIG�N��� PK�_FIL	$T�HKYMPANE��  	$DUMMY12 � �u3|4|�RG�_STR1 � $TITP/$I��1�{������5�6��7�8�9�0 ��z�����U1�1�1 '1
'�2"�SBN_C�FG1  8 �$CNV_JN�T_* |$DATA_CMNT�!$FLAGS��*CHECK�!��AT_CELLS�ETUP  �P $HOMEW_IO,G�%�#�MACRO�"RE�PR�(-DRUNj� D|3SM5�� UTOBACK�U0 $�ENAB��!EV�IC�TI �� D� DX!2S�T� ?0B�#$IN�TERVAL!2D�ISP_UNIT�!20_DOn6ER=R�9FR_F!2{IN,GRES�!�0Q_;3!4C_�WA�471�:OFFu_ N�3DELH�LOGn25Aa2c?i1@N?�� �-M�� W+0�$�Y $DB� 6CkOMW!2MO� x21\D.	 \r;VE�1$F��A{$O��D�B�C�TMP1_F�E2��G1_�3�B�2����AXD�#
 �d $CARD�_EXIST4�$FSSB_TY�PuAHKBD_YS�B�1AGN Gn� $SLOT�_NUMJQPREV,DBU� g1� �;1_EDIT1� � 1G=�� S�0%$EP<�$OP��AETE_OK�RUS�P_CR�Q$;4�V� 0LACIw1�RAP�k �1x@ME@$D�V�Q�Pv�Ah{oQL� OUzR ,mA�0�!� =B� LM_O�^e=R�"CAM_;1� xr$A�TTR4NP� AN�N�@5IMG_H�EIGHQ�cWI7DTH4VT� �U�U0F_ASPE�CQ$M�0EX�P��@AX�f�C�FT X $�GR� � S�!�@B@NFLI�`t� �UIRE 3dTuGI�TCHC�`N� S&�d_L�`�C�"�`�EDlpE� J�4S��0� �zsa�!ip;G�0 � 
$WARNM�0f�!,P�� �s�pNST� C�ORN�"a1FLT�R�uTRAT� Tv�p H0ACCa1����{�ORI�
`"S={RT0_S��B�qHG,I1� [ Tp�"3I�9�TY�D,P*2 ��`w@� �!R*HED�cJ* C��2��U3��4��5��6��U7��8��94�qO�$ <� $p6xK3 1w`O_M�@��C t � E�#6NGP�ABA � �c��ZQ���`���@Bnr��� ��P�0X����x�p�P@zPb26����"J�S_R��BC�J��3�JVP��tBS���}Aw��"�@G CP�_*0OFSzR @� RO_K8���a�IT�3��NOM_��0�1ĥ34 �pPT �� $���AxP��K}EX�� �0�g0I01��p�
$TyFa��C$MD3���TO�3�0U� �� ��Hw2�C1|�EΡg0wE{vF0�vF�40CPp@�a�2 
P$A`PU8�3N)#�dR�*�AX�!sDETAI�3BUFV�p@�1 |�p۶�pP�IdT� PP[�M�Z�Mg�Ͱj�F[�SIMQSI�"0��A�.����Pkx T�p|zM��P�B�F�ACTrbHPEW�7�P1Ӡ��v��MC�d� �$*1JqB�p<�*1DECH��H��a� � �+PNS_EMP���$GP���,P_���3�p�@Pܤ��TC��|r��0�s��b��0�� �B���!
���J�R� ��SEGFRR��Iv �aR�Tkp9N&S,�PVF4��>� &k�Bv �u�cu��aE�� !2��p+�MQ��E�SIZ�3����T��P�����>�aRSINF��� ��kq���������LX�����F�CRCMu�3CClpG��p� ��O}���b�1��������2�V�DxIC��C ���r����P��{� SEV �zF_�եF�pNB0�?�p�����A�! �r �Rx����V�lp�2ݠ�aR�t�,�g"�qR>Tx #�5��5"2��uAR���`CNX�$LG�p��B�1  `s�P�t�aA�0{��У+0R���tME`�`!BupCrRA 3�tAZ�л�pc�OFT�FC�b�`�`FNpp���1��ADI+ �a%��b�{��p$�pSp�c�`S�P��a&,QMP6�`Y�3��IM'�pU��aUw  $>�TITO1��S�S�!��$�"0�?DBPXWO��=!��$SK��F�DB�"�"@�PR8� 
� ����# >�q1$���$��+�L9$�?(�V�%@?R4Cr&_?R4ENE�Ƃ'~?(�� RE|�pY2(H ��OS��#$L�3$�$3R��;3�MVO�k_D@!V�ROS�crr�w�S���CRIoGGER2FPA�S|��7�ETURN0Bn�cMR_��TUː�[��0EWM%�ơ�GN>`��RLAȜ��Eݡ�P�&$P�t�'�@4a��C�DϣV�DXQ��4��1��MVGO_AWAYRMO#�aw!_�DCS_o)  `IS# � �� �s3S�AQ�� 4Rx�ZSW�AQ�p��@1UW��cTNTV)�5RV
a���|c���Wƃ��JB��x0���SAFEۥ�V_S}V�bEXCLUU�:;��ONL��c1Yg�~az�OT�a{�HI_V? ��R, M�_ *�0� ��9_z�2� �"P;SGO  +�rƐ m@�A�c~b���w@���V�i�b�fANNU�Nx0�$�dIDY�UABc�@Sp�i�a+ ��j�fΰAPIx2,���$F�b�$ѐO�T�@A $DUMMY��Ft��Ft�±� 6U- ` !�HE�|s���~bc�B@ SUFFmI��4PCA�UGs5Cw6Cq�!wMSWU. 8!��KEYI��5�TM`�1�s�qoA�vINޱpE��!, / D��oHOST�P!4� ��<���<�°<��p<�cEM'���Z�F��p�L� UL��0 � �	����D�T�01 � �$��9USAMPL�о�/���決�$ I�@갯 $SUB ӄ��w0QS�����#��SAV�����c�S�< 9�`�fP$�0E�!� YN_B�#2� 0�`DI�d�pO�|�m��#$F�R_�IC� �ENC�2_Sd3  ��< 3�9���� cgp����4�"��2�rA��ޖ5�� �`ǻ�@Q@K&D-!<�a�AVER�q�����DSP
���PC_�q��"�|�ܣ�oVALU3�HE��(�M�IP)���OkPPm �THЈ*��S" T�/�Fb�;�d����d D��q��16 H(rLL_DUǀ�a�@��0k���֠OT�"U��/���R_N_OAUTO70�C$}�x�~�@s��*|�C� ��C� 2��!z�L�� 8/H *��L� � ��Բ@sv��`� �� � ����Xq��cq���q��T�q��7��8��9���0���1�1 �1�-�1:�1G�1T�1*a�1n�2|�2��U2 �2-�2:�2G�U2T�2a�2n�3|ʥ3�3� �3-�3�:�3G�3T�3a�3
n�4|������9 <���z�ΓK�I����H硵BaFE8q@{@: ,��&a1?�pP_P?��>�
����E�@���!QQ���;fp$TP~�$VARI�����,�UP2Q`< W�߃TD��g�����`�������_BAC�"= T2����$�)�,+r³�p IF�I��p�� q M�P�"�l@``>t� ;��6����ST����T��M ����0	��i���F����������kRt ����F?ORCEUP�b܂�FLUS
pH(N𒰚 ��6bD_CM�@E�7N� (�v\�P��REM� Fa���@j���
Kr�	N���EFF/�̎�@IN�QOVܣ�OVA�	TR3OV DT)��DTMX:e �P :/��Pq�vXpCLN _�p��@ �2�	_|��_T: �*|�&PA�QDI���1��0�Y0RQm�_+qH���M���CL�d#�R�IV{�ϓN"EAR6/�IO�PCP��2BR��CM�@N �1b 3GCLF��!DY�(��a�#5T�DG���� ��%(�FSS� )�? P(q1�1��`_1"811R�EC13D;5D6O�GRA���@��i���PW�ON2EBUG�S�2��C`gϐ_E Azg`�TERM�5yB�5���ORIw��0C�5���S�M_-`���0D�9T�A�9E�9UP��F�� -QϒA��P�3�@B$SEG�GJ� EL�UUSE.PNFI��pBx���1@��4>DC$UF�P��$���Q�@"C���G�0T������SNSTj�PATxۡg��APTHJ�A�E*�Z%qB\`F�{E��F�q�pARxPY�aSHFT͢qA�AX_SHOR$�>��6% @$GqPE���GOVR���aZPI@P�@$U?r *aAYLO���j�I�"d��A8ؠ��ؠERV��Q i�[Y)��G�@R��i�e��i�R�!P�uA�SYM���uqAWJ�G)��E��Q7i�RD�U[d�@i�U��C��%UP���P���WORڒ@M��k0SM5T��G��GR��3�aPA�@��p5�'�_H � j�A�'TOCjA7pP]Pp$OPd�O��C��%�p�O!��R%E.pR�C�AO�?��Be5pR�EruIx|'QG�e$PWR) 3IMdu�RR_$s��\5��B Iz2H8��=�_ADDRH�H_LENG�B�q�qT:�x�R��So�J.�SS��SK�����0� ��-�SE*��ھrSN�MN1K�	�j�5�@r�֣O�L��\�WpW�Q�>pACRO�p���@H �����Q� ��OUPW3�b_>�I��!q�a1��������|�� ������-���:���ViIOX2S=�D��e��]���L $x��p�!_OFF��^_�PRM_�̱_HTTP_�H��wM (�pOBJ�"l�pG�$H�LE�C���ٰN � \9�*�AB_�T��b
�S�`�S��LV���KRW"duHITC�OU?BGi�LO�q����d� Fp�k�GpSS� ���HQWh�wA��O.��`�INCPUX2VISIO��!��¢.��á<�á-� �IO�LN)�P 87�R�'���$SL�b�d PUT_��$�dp�Pz �� F�_AS2Q/�$ALD���D�aQT U�0�]P�A������PH�YG灱Z�Ͱ5�U9O� 3R `F����H�Yq�Yx�ɱvpP��Sdp���x��ٶ�&�UJ��S����N�E�WJOG�G �DIS��&�KĠ��3T |��AV��`_��CTR1S^�FLA�Gf2&�LG�dU ��n�:��3LG_SIZ��ň��,=���FD��I���� Z �ǳ��0�Ʋ�@s�� -ֈ�-�=�-���-��0<-�ISCH_��DqR��N?���V��EAE!2�C��n�U�����`L�Ӕ�DAU��EA��Ġt�����GHr��I�BOO>)�WL ?`�� �ITV���0\�REC�SCRf 0�a��D^�����MARG ��`!P�)�T�/ty�?I�S�H�WW�I����T�JGM��MNC�H��I�FNKEY���K��PRG��UqF��P��FWD��HL�STP��V`��@�����RSS�H�` �Q�C�T1�ZbT�R ���U����� |R��t�i���G��8PCPO��6�F�1�M���FOCU��RGE]XP�TUI��I���c��n��n�� ��ePf���!p6�eP7�9N���CANAI�jB޾�VAIL��CL�t!;eDCS_HI�4�.��O�|!�S Sn��^I�BUFF1XY�5�PT�$�� ��v��fĘ�1�A�rY�Y��P �����pO+S1�2�3����_�0Z � � ��aiE�*��ID%X�dP�RhrO�+��A&ST��R��Y�z�<! Y$EK&CK+���Z&m&�5�0[ L��o�0 ��]PL�6pwq�t^����t0��7�_ \ �`��瀰�7��#��0C��] ��C�LDP��;eTRQ�LI�jd.�094F�LGz�0r1R3�DM�R7��LDR5<4R5ORG.���e2(`�ŀ�V�8.��T<�4�d^� �q�<4��-4R5SB�`T00m��0DFRCLMC!D�?�?�3I@��MIC��d_� d���RQm��q�DSTB	�  ��Fg�HAX;b ��H�LEXCESHZr�rBMup�a`Z���B;d�!rB`��`a��F_A�J��$[�O�H0K�db \���ӂS�$MB��L�IБ}SREQUI�R�R>q�\Á�XDESBU��oAL� MPŁc�ba��P؃ӂ!BFoAND���`�`d�Ҙ��c�cDC1��I�N�����`@�(h?Npz�@q��o� �SwPST8� e�r7LOC�RI�p�EX�fA�p��AoA�ODAQP�f Xf��ON��(2MF�� ���f)�"I��%�e���T� �FX�@IG}G� g �q�@�"E�0��#���$R�a%;#7y��Gx��Vv<CPi�DATAw�pAE:�y��RFЭ�NV�h t $MD
�qIё)�v+�tń�tH�`�P�u�|��sANSW}��t�?
�uD�)�b�	@Ð�i �@CU��V��T0�eRR2�j� Dɐ�Qނ�Bd$OCALI�@F�G�:s�2�RIN��v��<��NTE���k�E���,��b����_Nl��ڂ��kDׄR�m�DIViFDH��@ـn�$V؀�'c!$��$AZ�����~�[���oH �$B�ELTb��!ACC�EL+��ҡ��ICRC�t����T/!���$PS�@#2LPq�Ɣ83������<� ��PATH����D����3̒Vp�A_� Q�.�4�B�Cᐈ��_MGh�$DDxQ���G�$FWh���p��m�����b�DE���PPABNԗR?OTSPEED����00J�Я8��@��~P$USE_�2�P��s�SY��c�ZA >qYNu@Ag���OFF�q�MO�UN�NGg�K�OL�H�INC*��a���q��Bj�L@�BENCS��q�Bđ���D��IN#"I̒��4�\B�ݠVEO�w�Ͳ23�_UPE�߳LOWL���00����D���BwP��� �1RyCʀƶMOSIV��JRMO���@GPE�RCH  �OV ��^��i�<!�ZD <!�c��d@�P��!V1�#P͑��L���EW��ĸUP�������TRKr�"AYLOA'a�� Q-�̒�<�1Ӣ`0 ��RTI$Qx�0 MO���МB@ R�0J��D��s�H�x���b�DUM2(��S_BCKLSH_C̒��>�=�q�#��U��ԑ���2�t�]ACLALvŲ�1n�PN�CHK00'%SD�RTY4�k��y�1r�q_6#2�_UM$Prj�Cw�_�SCL���ƠLMT_J1_�LO��@���q��E������๕�幘S�PC��7������P	Co���H� �PU�m�C/@�"XT_�c�C�N_��N��e���S	Fu���V�&#�����9�̒��=�C�u�SH6#��c����1�Ѩ��o�0�͑
��_�PALt�h�_Ps�W�_10���4�R�01D�VG�Jb� L�@J�OGW����TORQU��ON*�Mٙ�sRHљ�&�_W��-�_=��PC��I��I�I�%II�F�`�JLA.,�1[�VC��0�D(R�O1U�@i�B\J�RKU��	@DBOL_SMd�BM%`�_DLC�BGRV���C��I��H_p� �*COS+\�(LN�7+X>$ C�9)I�9)u*c,)b�Z2 HƺMY@!̳( "TH&-�)TH�ET0�NK23�I��"=�A CB6CB=�C�A�B(261C�616SBC�T25'GTS QơC��a�S$" �4c#�7r#$DUD�EX�1s�t��(R�6��(QQ|r�f$NE�DpIB U�\B$5��$!��!A�%Ep(G%(!LPH$U�2׵�2SXpCc%pC�r%�2�&�C�J�&!�V�AHV6H3�YLVhJV�uKV�KV�KV�KV
�KV�IHAHZF`RXM���wXuKH�KH�KH��KH�KH�IO2LORAHO�YWNOhJOuKUO�KO�KO�KO�KO�&F�2#1ic%�d�4GSPBALANgCE_�!�cLEk0H_�%SP��T&�b�c&�br&PFULC��hr�grr%Ċ1k�y�UTO_?�jTg1T2Cy��2N&� v�ϰctw�g�p�0Ӓ~���T��O���� �INSEGv�!�R�EV�v!���DIF���1l�w�1m�
�OB�q
����M�Iϰ1��LCHW3AR��
�AB&u�?$MECH,1� X:�@�U�AX:�P��pY�G$�8pn 
Z���|���ROBR�C�R��N� (��MSK_�`f�p WP Np_��R����΄ݡ�1��ҰТ`΀ϳ��΀"�IN�q��MTCOM_�C@j�q  �L��p��$NOR�E³5���$�r� 8� GR�E�S�D�0ABF�$XYZ_DA5A���DEBU�qI��Q��s �`$�COD��� ��k�F��f�$BUFIN�DXР  ��M{OR��t $-��U��)��r�B����͓�Gؒu � $SIMULT ৐~�� ���OBJ�E�` �ADJUS<>�1�AY_Ik���D_����C�_FIF�=�T� ��Ұ ��{��p� �����p�@:��D�FRI��ӥMT��RO� ��E�<���OPWO�ŀ�v0��SYSByU�@ʐ$SOP�ȸ��#�U"��pPR�UN�I�PA�DpH�D����_OU��=��qn�$}�I�MAG��ˀ�0Pf�qIM����IN��q���RGOVRDȡ:���|�P~���Р�0L_6p���i��SRB���0��M���EDѐF� ��N�`M*����'��˱SL�`ŀw x $OVSL�vwSDI��DEXm�@g�e�9w�����V� ~�N���w����Û��ȳ�M���q<�>�� x HˁE�^F�ATUS����C�0àǒ��BTMT����If���4����(�ŀy DˀEz�g���PE�r����8�
���EXE��V���E�Y�$Ժ ŀz �@ˁ��UP{�h�$�p��XN���9x�H� �PG"��{ h $SUB��c�@_��01\�_MPWAI��P��&��LO��-�F�p��$RCVFAI�L_C�-�BWD�"�F���DEFSP>up | Lˀ`��D�� U�UNI��S���R`����_L�pP�����	P�ā}��� B�~�о�|��`ҲN�`KE)T��y���P� $��~���0SIZE��ଠ{���S<�O�R��FORMAT�/p � F���rEM2R��y�UX�����PLI7�ā � $�P_S�WI���͐�_P�L7�AL_ ��ސR�A��B�(0C���Df�$Eh�����C_=�U� ?� � ����~�J3�0����TI�A4��5��6��MOM������ �B�AD��*��l* PU70NR�W��W R����� A$PI�6 ���	��)�4�l�}69��Q���c�S/PEED�PGq�7 �D�>D����>�tMt[��SA�M�`痰>��MOV���$��p�5�H�5�D�1�$2�@������{�Hip�IN?,{�F(b+�=$�H*�(_$�+�+G�AMM�f�1{�$GGET��ĐH�D��z��
^pLIBR�Ѻ�I��$HI��_���Ȑ*B6E��*8A$>G086LW=e6\<�G9�686��R��ٰV���$PDCK�Q�H�_����;"��z�.%�7�4�*�9� �$_IM_SRO�D�s0"���H�"�LE�!O�0\H��6@�@�U�� �ŀ�P�qUR_SCR�ӚAZ���S_SAVE_DX�E��NO��CgA �Ҷ��@�$����I� �	�I� %Z[� �� RX" ��m���"�q� '"�8�Hӱt@�W�UpS��хDM��O㵐.'}q��Cg@���@ʣ����S�M�A�Â� � $P9Y��$WH`'�NGp���H`��Fb��0Fb��Fb��PLM����	� 0h�H�{�X��O���z�Z�eT�M����# pS��C��O@__0_B_�a��_%�� |S����@	�v ��v �@���w�v��EM��% -�cu�B������ftP���PM��QU� ŉU�Q��A-�QT�H=�HOL��QH�YS�ES�,�U�E��B��O#��  -�P0�|�gAQ����ʠu���O��ŀ��ɂv�-�A;ӝROG��a2D�E�Â�v�_�ĀZ�INFOB&��+����b�R�OI킍 ((@SLEQ/�#�������o���S`c0O��0�01EZ0N9Ue�_�AUT�Ab�COPY��Ѓ�{�
�@M��N�����1�4P�
� ��RGI��͏��X_�Pl�$P�����`�W��P���j@�G���EXT/_CYCtbR���p����h�_NAƹ!$�\�<�RO��`]�� � m��POR�ㅣ�.��SRVt�)����DI �T_l���Ѥ@{�ۧ��ۧ �ۧ5٩�6٩7٩8��R�S��B쐒��$�F6���PL�A�A^�TAR��@E `�Z�����<��d� ,�(@FLq`h��@YN�L���M�C���P�WRЍ�쐔e�D�ELAѰ�Y�pA�D#qX� �QSK;IP�� ĕ�x�-O�`NT!� ��P_x�-�ǚ@�b�  1�1�1Ǹ�?� � ?��>��>�&�>�3�z>�9�J2R;n쐖 4��EX� TQ����ށ�Q����[�KFд���RDCNIf� �U`�X}�R�#%M!*�0�)��$�RGEAR_0I9O�TJBFLG�i&gpERa��TC݃��|����2TH2N���� 1� ��Gq T�0 �$���M���`Ib���Q�REF�1��� l�h��ENAB��lcTPE?@��� !(ᭀ����Q�#�@~�+2 H�W���2������"�4�F�X�j�3�қ{��������j�4�Ҝ��
��P.�@�R�j�5�ҝu�@����������j�6�����(:Lj�7�ҟo������ ����8�Ҡ���"4Fj�SwMSK��  ��+@��E�A��REoMOTE�������@ "1��Q�IO��5"%I��P��PO9Wi@쐣  ��� ��X�gpi�쐤��Y"�$DSB_SIG!N4A�Qi�̰C��>%/S232%�Sb�i�DEVICEUS�#�R�RPARIT|�!OPBIT�Q���OWCONT�R��Qⱓ�RCU�� M�SUXTAS�K�3NB��0�$TA[TU�P�S@@R쐦F�6�_�PC}��$FREEFR�OMS]p�ai�GE�TN@S�UPDl�A�RB�#P%0����� !m$USAࢰ�az9�L�ERI��0���pRY�5~"_ľ@��P�1�!�6WR	K��D9�F9Х?FRIEND�Q4b�UF��&�A@TOO�LHFMY5�$L�ENGTH_VT��FIR�pqC�@�yE� IUFIN�R:���RGI�1�OAITI:�xGX�l�I�FG2�7G1a�0���3�B�GPRR�DA���O_� o0e�I1R�ER�đ�3&���TCp���AQJV �G|�.2���F��1�!d� 9Z�8+5K�+5��E�y�|L0�4�X �0*m�LN�T�3Hz��8P9��%�4�3G��W�0�W�RdD�Z��T�ܳ�pK�a3d��$cV 2���1��RI1H�02K2sk3K3Jci�aI�i��a�L��SL��R$Vؠ�BV�EVk�]V*R
��� �,6Lc����9V2F{/P:B��PS_�E��$rr�C��γ$A0��wPR���v�U�cSk�� {��8��� 0���VX`�!�tX`��0P��Ё�
�5SK!�� �-qR��!0�4��z�NJ AX�!h��A�@LlA��A�THIC�1�������1�TFE���q>�IF'_CH�3A�I0�����G1�x������t9�Ɇ_JF҇�PR(���RVA=T�� �-p���7@����DO�E��CsOU(��AXIg��OFFSE+�TRIG�SK��c������e�[�K�Hk���8��IGMAo0�A-���ҙ�ORG_UNsEV��� �S�~쐮d �$��z����GROU���ݓTO2��!ݓDSP��JOG'��#	�_P'�2OR����>P6KEPl�IR��0�PM�RQ�AP��Q��E�0q�e���ScYSG��"��PG��BRK*Rd�r�3�-��������ߒ<pADx��ݓJ�BSOC�� N�DUMMY�14�p\@SV�PD�E_OP3SFS�PD_OVR��bٰCO��"�OR-��N�0.�Fr�.��OV�SFc�2�f��F��!4�S��RA��"LCHDL�R�ECOV��0�Wb�@M�յ�RO3���_�0� @܄ҹ@VERE�$7OFS�@CV� 0BWDG�ѴC��2j��
�TR�!��E�_FDOj�MB_�CM��U�B �BL =r0�w�=q�tVfQ�Ґx0sp��_�Gxǋ�A�M��k�J0������_�M��2{�#�8$�CA�{Й���8$�HBK|1c��IO␅.�:!aPPA "�N�3�^�F���:"�?DVC_DB�C��@d�w"����!��1����ç�3����ATIEO� �q0�UC�&CAB�BS@�PⳍP�Ȗ��_0~c�SUBCPUq��S�Pa aá�}0�S�b��c��r"ơ$HW_C���:c��Ic�A�A-�l$UNI5T��l��ATN�f�����CYCLųN�ECA��[�FLT?R_2_FI���(��}&��LP&�����o_SCT@SF_��aF����G���FS|!�¹�CHAA/���8��2��RSD�x"�ѡb�r�: _T��PcRO��O�� EM��_��8u�q 1u�q��DI�0e�?RAILAC��}RMƐLOԠdC��:a�nq��wq����PRJ��SLQ�pfC��z� 	��FUNCŢ�rRINkP+a�0 ̆�!RA� >R �
Я�ԯWAR��BLFQ��A0�����DA�����LDm0�a�B9��nqBTI�vrbؑ���PRIA,Q1�"AFS�P�!������`%b���Mr�I1U�DF_j@ؖ�y1°LME�FA��@HRDY�4��P�n@RS@Q�0"�MULSEj@f�b�q� �X��ȑ����$.A$�1�$c1Ó���7� x~�EG70ݓ��q!AR����0�9>B�%��AXE.��ROB��W�A4�_�-֣SY���!6���&S�'WR���-1���STR��5�:9�E�� 	5B��=QB90�@6�������OT�0o 	$�ARY8�w20�Ԛ�	%�FI��;�$LINK�H��1%�a_63�5�q�2XYZ"��;�qH�3@��1�2�8{0	B�{D��� CFI��6G��
�{�_J��6��3NaOP_O4Y;5�FQTBmA"�BC
�z�DU"�66CTURN3�vr�E�1�9�ҍGFL�`���~ �@�5<:7�� W1�?0K�Mc��68Cb�vrb�4�ORQ��X�>8�#op ������wq�Uf����N�TOVE�Q��M;����E#�UK#�UQ"�VW �ZQ�W���Tυ� ;� ����QH�!`�ҽ��U��Q�WkeK#kecXE)R��	GE	0��S�dAWaǢ:D���0�7!�!AX�rB !{q��1uy-! y�pz�@z�@z6P z\Pz� z1v� y�y�+y�;y� Ky�[y�ky�{y�x�y�q�yDEBU��$����L�!º2WG`  AB!�,�r�SV���� 
w� ��m���w����1���1 ���A���A��6Q��\Q����!�m@��2CLAB3B�U������S  ÐER|��
0 � $�@ڳ Aؑ!p�PO���Z�q0w�^�_M�RAȑ� d r T�-�ERR�L�TYz�B�I�qV3@�cΑTOQ�d:`L� �d2�p ��|˰[! � p�`qT}0i��_V1�rP�a'�4�2-�2<�����@P�����F��$W��g��V_!�l�$�P����c���q"�	�SFZ�N_CFG_!� 4��?º�|�ų����8@�ȲW ]���\$� �n���Ѵ��09c�Q��(�FA�He�,�XEDM�(���H��!s�Q�g�P{R�V HELLĥ�� 56�B_BAS!�RSR��ԣo E�#S��[��1r�U%��2ݺ3ݺ4ݺU5ݺ6ݺ7ݺ8ݷ��ROOI䰝0�03NLK!�CAB� n��ACK��IN��T:�1�@�@ z�m�7_PU!�CO� ��OU��P� Ҧ) ���޶��TPFWD�_KARӑ��R�E~��P��(�Q�UE�����P
��C�STOPI_AL �����0&���㰑�0GSEMl�b�|�M��6d�TY|�SOK�}�DI�����(����_TM\�MANR�Q�ֿ0E+�|�$�KEYSWITCaH&	���HE
�OBEAT��cE� �LEҒ���U��F�O�����O_HOuM�O�REF�P�PRz��!&0��Cr+�OA�ECO��xB�rIOCM�D8׵�]���8�` G� D�1����U���&�MH�»P�CFO�RC��� �'쾠��OM�  �� @V��|�U,3P�� 1-�`� 3-�4���NPX_AS�Ǣ� 0ȰADD|����$SIZ���$VARݷ TKIP]�\�2�A�������]�_� �"�S꣩!Cΐ��FRIF⢞�S�"�c���NF��V ��` �� x�`SI�TE�S�R6SSGL(T�2P&��AU�� ) OSTMTQZPm �6BW�P*SHO9Wb��SV�\$߽� ���A00P�a�6�@�PJ�T�5�	6�	U7�	8�	9�	A�	 � �!�'��C@�F�0u�	f0u�	 �0u�	�@u[Pu�%121?1L1�Y1f1s2�	2��	2�	2�	2�	2��	2�	222�%222?2L2�Y2f2s3P)3��	3�	3�	3�	3��	3�	333�%323?3L3�Y3f3s4P)4��	4�	4�	4�	4��	4�	444�%424?4L4�Y4f4s5P)5��	5�	5�	5�	5��	5�	555�%525?5L5�Y5f5s6P)6��	6�	6�	6�	6��	6�	666�%626?6L6�Y6f6s7P)7��	7�	7�	7�	7��	7�	777�%727?7,i7�Y7Fi7s�VP��UPD�� � ��|�԰��YS�LOǢ� �  z��и���o�E��`>�8^t��АALUץ�����CU���wFOqIgD_L�ӿuHI�z�I�$FILE_����t��$`�JvS�A��� h���E_BLCK�#�C>,�D_CPU<�{� <�o����tJr���R ��
PWl O� ��LA���S��������RUN F�Ɂ��Ɂ����F�����ꁬ��TBC�u�C� �X ;-$�LENi���v������I��G�L�OW_AXI�F)1��t2X�M����hD�
 ��I�� ���}�TOR����Dh��� L=��⇒�8s���#�_MA`�8ޕ��ޑTCV����T���&��ݡ�����J�����J����MDo���J�Ǜ ����
���2��� v���l��F�JK��VKi�hΡv�Ρ3��J0㤶ңJJڣJJ�A�ALң�ڣ��42�5z�&�N1-�9�(��␅�L~�_Vj�������� ` �GROU�pD��}B�NFLIC�����REQUIREa�EBUA��p����2¯�����c�ޞ� \��APKPR��C���
�;EN�CLOe�ɇS_M v�,ɣ�
����� ���M�C�&���g�_MG�q�C� �{�9����|�BRKz�NOL��|ĉ R��_LI�|��Ǫ�k�J����P 
���ڣ�����&���D/���6��6��8���Y����� ���8�%�W�2�e�PATHa�z�p�z�=�hvӥ�ϰ�x�CN=��CA�����p�INF�UC��bq��CO�UM��YZ������q�E%���2������P�AYLOA��J2=L3pR_AN��<�L��F�B�6�R�{�R_F2LSHR��|�LOG��р��ӎ�>��ACRL_u��Ր����.���H�p��$H{���FLEX�
��J�� :�/����6�2�`����;�M�_�F16� ����n���������ȟ��Eҟ�����,� >�P�b���d�{�������������5�T��X��v���E ťmFѯ����� ��&�/�A�S�e�+p|�x�� � ��0����j�4pAT����6n�EL  �%ø�J���ʰJE��C�TR�Ѭ�TN��F�&��HAND_V�B[
�pK�� $F2{�6� �r�SWi��("U���� $$Mt�h�R ��08��@<b 35��^6�A�p3�k��q{9t�A(�̈p��A��A�ˆ0���U���D��D��P2��G��IST��$A4��$AN��DYˀ� {�g4�5D���v�6�v瀑�5缧�^�@��P �����#�,�5�>�(#�� &0�_��ER!V9�SQASYM$��] �����x�������_SHl����� ��sT�(����(�:�JA���S�cir��_VI�#Oh9�``V_UNI��td�~�J���b�E�b��d ��d�f��n�������H��uN���(!2�H������"Cq3EN� �pDI��>��ObtC�Dpx�� ��2IxQA�q��q ��-��s �� s������ ��OMMEB��rr/�TVpPT�P ���qe�i�A���P�x ��yT�P�j� $DUM�MY9�$PSm_��RFq�  ��:� s���!~q�� X����K�ST�s�ʰSBR��M�21_Vt�8$S/V_ERt�O��z����CLRx�A  O�r?p? Oր �� D $GLOB���#LO��Յ�$�o��P�!SYS�ADR�!?p�pT�CHM0 � ,x����W_NA���/�e���D�SR~��l (: ]8:m�K6�^2m�i7 m�w9m��9���ǳ��� ����ŕߝ�9ŕ�� �i�L���m��_�_��_�TD�XSCRE��ƀ�� ��ST�F���}�pТ6��C�] _v AŁ� 9T����TYP�r�@K��u�!u���-O�@IS�!��uvD�UE{t� �����H�S���!RSM�_�XuUNEXCcEPWv��CpS_�� {ᦵ�ӕ���÷����COU ��� [1�O�UET�փr|���PROGM� {FLn!$CU��cPO*q��c�I_�p}H;� � 8��.N�_HE
p��Q�~�pRY ?����,�J�*��;�OU}S�� � @d�~��$BUTT���R@���COLUMx�íu�SERVc#�=�PANEv Ł�� � �PGEU�!�F��9�)$H�ELP��WRETER��)״���Q� �����@� P�LP �IN��s�PQNߠw v�1���ލ� ���LNN�� ����_���k�$H��M TEqX�#����FLAn ^+RELV��D4p��������M��?�,��ӛ$����P�=�USRVIEWNŁ� <d��pU�p�0NFIn i�F�OCU��i�PRI�LPm+�q��TR�IP)�m�UNjp{t� QP��Xu�WARNWud�SRWTOLS�ݕ�����O|SORN��R�AUư��T��%���VI|�zu� {$�PATHg���CACHLO9G6�O�LIMybM����'��"�HOSTN6�!�r1�R��OBOT5���IMl� ��C� g!��E����L���i�VCPU?_AVAILB�O�+EX7�!BQNL�(����A�� Q��Q ���ƀ�  QpC����@$TOO�L6�$�_JMP�� �I�u$�SS�!$��VSHsIF��|s�P�p��6�s���R���O�SURW�pRA#DIz��2�_�q��h�g! �q)�LU�za$OUTPU�T_BM��IM�L�oR6(`)�@TI�L<SCO�@C e�;��9��F��T ��a��o�>�3�����w�2u�P{t9��%�DJU��|#��WAIT��h�����%ONE���YBOư �� $@p%�C��SBn)TPE��NEC��x"�$t$���*B_T��R��%�q�R� ���sB�%�tM �+��t�.�F�R!݀v��OPm�MAS�W_DOG�OaT	��D����C3S�	�O2D�ELAY���e2JO��n8E��Ss4'#J��aP6%�����Y_ ��O2$��2���5��`�? ��ZAB�CS��  $��2��J�
���$$�CLAS������AB���'@@V�IRT��O.@AB�S�$�1 <E�� < *AtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v�����M@[�AXLր`�&A��dC  ���IN8��ā��PRE������LARM�RECOV �<I䂥�NG�� �\K	 A   �J�\�M@PPLIC��?<E�E��HandlingTool ��� 
V7.50�P/28[�  ��X���
�_�SW�� UP*A� ��F0ڑ�����A���� 2)0��*A���:����(�(B �7DA5�� �'@Y�@<��None������� ��T���*A4I�xl�_��V����g�UTOB�ค�����HGAPON�8@��LA��U��D [1<EfA����������� Q �1שI Ԁ� �Ԑ�:�i�n�����#B)B ���\�HE�Z�r�HTTHKY�� $BI�[�m�����	� c�-�?�Q�o�uχϙ� �Ͻ��������_�)� ;�M�k�q߃ߕߧ߹� �������[�%�7�I� g�m��������� ����W�!�3�E�c�i� {��������������� S/A_ew� ������O +=[as��� ����K//'/9/ W/]/o/�/�/�/�/�/ �/�/G??#?5?S?Y? k?}?�?�?�?�?�?�? COOO1OOOUOgOyO �O�O�O�O�O�O?_	_�_-_K_Q_��(�TO�4�s���DO_CL�EAN��&��SNMw  9� ��9oKo]ooo�o�DS�PDRYR�_%�H	I��m@&o�o�o #5GYk}�����"���p�Ն �ǣ�qXՄ��ߢ��>g�PLUGGҠ�W\ߣ��PRC�`B`E9��o�=�OB���o&�SEGF��K ������o%o����p#�5�m���LAP�o ݎ����������џ� ����+�=�O�a���TOTAL�.���_USENUʀ׫� �X���R(�RG_�STRING 1���
�Mڜ�Sc�
��_I�TEM1 �  n c��.�@�R�d�v��� ������п������*�<�N�`�r�I�/O SIGNA�L��Tryout Mode��Inp��Sim�ulated��Out��OV�ERR�` = 1�00�In c�ycl���Prog Abor������Statu�s�	Heart�beat��MH� FaulB�K�AlerUم�s߅ߗ߀�߻��������� �S���Q��f� x������������ ��,�>�P�b�t���8����,�WOR���� ��V��
.@R dv��������*<N`PO��6ц��o� ����//'/9/ K/]/o/�/�/�/�/�/p�/�/�/�DEV� *0�?Q?c?u?�?�? �?�?�?�?�?OO)O�;OMO_OqO�O�O�OPALTB��A���O �O__,_>_P_b_t_ �_�_�_�_�_�_�_opo(o:o�OGRI�p ��ra�OLo�o�o�o�o �o�o*<N` r������`o��RB���o�>�P� b�t���������Ώ�� ���(�:�L�^�p�<���PREG�N�� .��������*�<� N�`�r���������̯�ޯ���&����$�ARG_��D ?�	���i���  	�$��	[}�]�}���Ǟ�\�SBN�_CONFIG Si��������CII_SAVE  ��۱Ҳ\��TCELLSET�UP i�%HOME_IO��~��%MOV_�2�8�REP���V�UTOBACK
��ƽFRwA:\�� ��,����'` �����<���� �����$�6�c�Z�lߙ��Ĉ������������� !凞��M�_�q��� ��2���������%� 7���[�m�������� @�������!3E$���Jo��������INI�@ꨔε��MESSAG����q��ODE_D$����O,0.��PAU�S�!�i� ((Ol����� ��� /�//$/ Z/H/~/l/�/�'ak?TSK  q��<���UPDT%��d0;WSM_kCF°i�е|U�'1GRP 2h�V93 |�B��A�/�S�XSCRD+11�
1; ��� �/�?�?�? OO$O�� ߳?lO~O�O�O�O�O 1O�OUO_ _2_D_V_�h_�O	_X���GRO�UN0O�SUP_kNAL�h�	��n�V_ED� 11;�
 �%-BCKEDT-�_`�!oEo$���a��oʨ����ߨ����e2no_˔o�o�b����ee�o"�o�oED3�o�o ~[�5GED4�n#��� ~�j���ED5Z��Ǐ6� ~���}���ED6����k��ڏ ~G���!�3�ED7��Z��~� ~�V�şןED8F�&o��Ů}����i�{��ED9ꯢ�W�Ư
`}3�����CRo �����3�տ@ϯ�����P�PNO_DEL��_�RGE_UNU�SE�_�TLAL_?OUT q�c��QWD_ABOR�� �΢Q��ITR_�RTN����NO�NSe���C�AM_PARAM� 1�U3
 8�
SONY X�C-56 234�567890�H �� @����?���( АTV�|[r؀~�X�HR5k�|U�Q�߿��R57����Af�f��KOWA �SC310M|[�r�̀�d @ 6�|V��_�Xϸ��� V��� ���$�6��Z��l��CE_RIA�_I857�FF�1��R|]��_LIO4W=� ���P<~�F<�GP� 1�,����_GYk*C* Y ��C1� 9� �@� G� �CLCU]� d� l� s�QR� ��[�m� �v� � �� ��W C�� �"�|W��7�HEӰONF�I� ��<G_PR/I 1�+P�m� �/���������'CHKPAUS��  1E� , �>/P/:/t/^/�/�/ �/�/�/�/�/?(??�L?6?\?�?"O������H�1_MOR��� �0�5 	 �9 O�?$OO HO6K�2	���=9"��Q?55��C�PK��D3P������a�-4�O__|Z
�OG_�7�PO�� ȕ�6_��,xV�ADB���='�)
mc�:cpmidbgX�_`��S:�(�����Yp�_)o�S`��BBi�P�_mo8j��(�Koo�o9i�(��og�o�o�o�Lnf�oGq:I�ZD�EF f8��)��R6pbuf.t�xtm�]n�@�����# 	`(Ж�A=�L���zMC�21��=��9���4��=�n׾�Cz  �BHBCCo�C�|��CqD���C���C��{iSZE@D����F.��F���E⚵F,�E�ٙ�E@F��N�IU��I?�O�I<#I6?�I�SY��)�vqG���Em�U(�.��(�(�1�<�q�G�x2��eҢ �� a�D�j��E�e��EX��EQ�EJP �F�E�F� �G�ǎ^F �E�� FB� �H,- Ge���H3Y���  �>�33 ����xV  n2xQ@F��5Y��8B� A�A�ST<#�
� ��_'�%��wRSMO�FS���~2�yT}1�0DE �O� c
�(�;�"� � <�6�z�R��X�?�j�C4��SZ�m� W��{�m�CR��B-G�C�`@$��q��T{�FPROG %i�����c�I��� �Ɯ�f�K�EY_TBL  �vM�u� �	
��� !"#�$%&'()*+�,-./01c�:�;<=>?@AB�C�pGHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������p����͓���������������������������������耇��������������������!j�LCK��.�j����STAT���_A�UTO_DO����W/�INDT_ENB߿2R��9�+��T2w�XSTOP�\߿2TRLl�LE�TE����_SCREEN i�kcsc��U���MMENU 1� i  < g\��L�SU+�U��p3 g������������ 2�	��A�z�Q�c��� ������������. d;M�q�� ����N% 7]�m��� /��/J/!/3/�/ W/i/�/�/�/�/�/�/ �/4???j?A?S?y? �?�?�?�?�?�?O�? O-OfO=OOO�OsO�O �O�O�O�O_�O_P_�Sy�_MANUAyL��n�DBCOU��RIG���DBN�UM�p��<���
��QPXWORK 1!R�ү�_oO�.o@oRk�Q_AWA�Y�S��GCP r��=��df_AL�P�db�RY�������X�_�p 1"�� , 
�^���o �xvf`MT�I^�rl@|�:sONTIM�כ����Zv�i
�õ�cMOTNEN�D���dRECOR/D 1(R�a��ua�O��q��sb �.�@�R��xZ���� ���ɏۏ폄���#� ��G���k�}�����<� ş4��X���1�C� ��g�֟��������ӯ �T�	�x�-���Q�c� u����������>�� ��)Ϙ�Mϼ�F�� �ϧϹ���:������� %�s`Pn&�]�o��ϓ� ~ߌ���8�J����� 5� ��k����ߡ�� J�����X��|��C� U����������0������	��dbTOL�ERENCqdB�ܺb`L�͐PCS_CFG )�k�)wdMC:\�O L%04d.C�SV
�Pc�)sA� �CH� z�P�)~���hMRC_OUT *�[��`+P SGN �+�e�r��#��10-MAY-20 10:59*V�17-FEBj9�:0rv PQ�8��)~�`�pa�m��P�JPѬVE�RSION �SV2.0.�8.|EFLOGI�C 1,�[ 	DX�P7)�PF."�PROG_ENB��o�rj ULSew ��T�"_WRST�JNEp�V�r`dEM�O_OPT_SL� ?	�es
 ?	R575)s7)��/??*?<?'�$TO  �-��?&[V_@pEX�Wd�u��3PATH ASA\�?�?O�/{ICT�aFo`�-�gds�egM%&ASTBF_TTS�x�Y^C��SqqF�PMAU�� t/XrMSWR.D�i6.|S/�Z!D_N�O0__T_C_�x_g_�_�tSBL_/FAUL"0�[3w/TDIAU 16M6�p�A12�34567890gFP?BoTofo xo�o�o�o�o�o�o�o ,>Pb�S�p-P�_ ���_s �� 0`����� )�;�M�_�q����������ˏݏ��|)UM�P�!� �^�T�R�B�#+�=�PME�fEI�Y_TEMP9 È�3@�3A �v�UNI�.(YN_BRK 2Y�)EMGDI_S�TA�%WЕNC2_SCR 3��1o"�4�F�X�fv����������#��ޑ14����)�;���t��ݤ5��� ��x�f	u�ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /߭P�b�t�� ��x� �߰���������
�� .�@�R�d�v���� ����������*�<� N���r����������� ����&8J\ n������� �"`�FXj| �������/ /0/B/T/f/x/�/�/ �/�/�/�/�/4?,? >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO ^OpO�O�O�O�O�O? �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �o�O�O�o�o�o
 .@Rdv��� ������*�<� N�`�r����o����̏ ޏ����&�8�J�\� n���������ȟڟ�����H�ETMODoE 16���W ��ƨ
R��d�v�נRROR_PROG %A��%�:߽�  ��TABLE  A�������#�L�RR�SEV_NUM � ��Q���K�S���_AUTO_ENB  ���I�Ϥ_NOh� �7A�{�R�  �*������������^�+��Ŀֿ迄��HISO�͡I�}�_�ALM 18A�� �;�����+ �e�wωϛϭϿ��_H���  A��|��4�TCP_�VER !A�!�����$EXTLO�G_REQ��{�V�SIZ_�Q�T�OL  ͡Dz���A Q�_B�WD����r���n�_�DI�� 9���}�z�͡m���ST�EP����4��OP�_DO���ѠF�ACTORY_T�UN�dG�EAT?URE :�����l�Han�dlingToo�l ��  - C�Englis�h Dictio�nary��ORD�EAA Vi�s�� Masteyr���96 H���nalog I/yO���H551���uto Soft�ware Upd_ate  ��J���matic Ba�ckup��Par�t&�ground Edit���  8\ap�Camera��F���t\j6R�elyl���LOADR�7omm��shq��oTI" ��co��
! o���p�ane�� 
!���tyle s�elect��H5�9��nD���oni7tor��48�����tr��Relia�b���adin�Diagnos�"����2�2 ual� Check S�afety UI�F lg\a��h�anced Ro�b Serv q� ct\��lUs�er FrU��D�IF��Ext. oDIO ��fiAs d��endr �Err L@��I%F�r��  �П��90��FCTN /MenuZ v'���74� TP In���fac  S�U (G=�p���k Excn g��3��High-wSper Ski+�  sO�H9 � m�munic!�on5sg�teur� �����V����c�onn��2��ENމ�Incrst�ru���5.fd�KAREL �Cmd. L?u�aA� O�Runw-Ti� Env��R��K� ��+%�s#�S/W��74��L?icenseT��  (Au* ogBook(Sy���m)��"
MACROs,V�/Offse��a�p��MH� ����p�fa5�MechS�top ProtL��� d�b i��Shif���j545�!xr ��#���,[�b ode Switch��m\e�!o4.�& pro�4���g��Multi�-T7G��net�.Pos RGegi��z�P���t Fun���3s Rz1��Numx ������9m�1�  �Adjuj��1 J7�7�* ����6�tatuq1EIK�RDMtot���scove�� ���@By- }uest1�$Go� � U5�\SNPX �b"���YA�"Li�br����#�� �$~@h�pd]0�J�ts in VCCCM�����0�  �u!��2 R�0�/�I�08��TMI�LIB�M J92:�@P�Acc>�F�{97�TPTX�+6�BRSQelZ0�M�8 Rm��q%��6�92��Unexc�eptr motn>T  CVV�P���KC����+-��~K  II)�VS�P CSXC�&.ac�� e�"�� t�@�Wew�AD� Q�8bvr nm�en�@�iP� a�0y�0�pfGri�dAplay !�� nh�@*�3R�1M-�10iA(B20k1 �`2V"  F����scii�lo{ad��83 M��yl����Guar�dO J85�0�mP'��L`���stuaPa9t�&]$Cyc����|0ori_ x%Da�ta'Pqu���cAh�1��g`� j� RLJam�5���IMI De-B(�\A�cP" #^0C~  etkc^0�asswo%q�)6�50�ApU�Xn�t��Pven�CT�qH�5�0YELLOW BO?Y���� Arc�0vi�s��Ch�Wel=dQcial4Izt�Op� ��gs�`k 2@�a��poG3 yRjT1 NEf�#HT� xyWbF��! �p�`gd`����p\� =P��JP�N ARCP*P�R�A�� OL��pSup̂fil��p��J�� ��cro�670�1C~E�d���SS�pe�tex��$ �P� So7 t^� ssagN5 <Q"�BP:� �9 "0�Q#rtQC��P�l0dpn�笔�rpf�q��e�ppmas�cbin4psy=n�' ptx]08��HELNCL �VIS PKGS9 �Z@MB &���B J8@IPE� GET_VAR� FI?S (Un�i� LU�OOL:� ADD�@29.KFD�TCm���E�@�DVp���`A�ТN�O WTWTEST �� f�!��c��FOR ��ECT� �a!� ALSE� ALA`�CPMO-130��� b �D: HANG FROMg��2���R709 DRA�M AVAILC�HECKS 54�9��m�VPCS �SU֐LIMCH�K��P�0x�FF WPOS� F�� q�8-12 C�HARS�ER6�O�GRA ��Z@AV�EH�AME��.SV��Вאn$��9�wm "y�TRCv�� SHADP�UP�DAT k�0��S�TATI��� M�UCH ���TI�MQ MOTN-�003��@OB�OGUIDE DAUGH���b��@�$tou� �@C� <�0��PATH�_��MOVET�� R�64��VMXPA�CK MAY A�SSERTjS��C�YCL`�TA��B�E COR 71��1-�AN��RC �OPTIONS � �`��APSH-�1�`fix��2�S�O��B��XO򝡞�_�T��	�i��0j��d�u�byz p wa��y�٠HI�������U�pb XSPD �TB/�F� \hcehΤB0���END�[CE�06\Q�p{ }smay n@��pk��L ��tr'aff#�	� ���~1from sy�svar scr��0R� ��d�DJUD���H�!A��/��SET ERR��D�P7����NDA�NT SCREE�N UNREA �VM �PD�D��P�A���R�IO gJNN�0�FI��}B��GROUNנD Y�Т٠�h�SVIP 53 Q�S��DIGIT �VERS��ká�N{EW�� P06�@=C�1IMAG�ͱ4���8� DI`����pSSUE�5��EPLAN JON�� DEL���157�QאD��CALL�I���Q��m���IP�ND}�IMG N�9 PZ�19��MwNT/��ES ���`LocR Hol�߀=��2�Pn� PG�:��=�M��can�����С: 3D� mE2view gd X��ea1 ��0b�pof Ǡ"�HCɰ�ANNO�T ACCESS? M cpie$E�t.Qs a� lo^MdFlex)a:���w$qmo G�sA�9�-'p~0��h0pa���eJ AUTO1-�0��!ipu@Т|<ᡠIABLE+�� 7�a FPLN:9 L�pl m� �MD<�VI�и�W�IT HOC�Jo~1Qui��"���N��USB�@�Pt� & remov����D�vAxis �FT_7�PGɰC�P:�OS-14�4 � h s 2968QՐOST�p � CRASH D�U��$P��WOR�D.$�LOGI�N�P��P:	�0�0�46 issue�E�H�: Slo[w st�c�`�6����໰IF�I�MPR��SPOT�:Wh4���N1STyY��0VMGR�\b�N�CAT��4oR�RE�� � 5�8�1��:%�RTU�!Pe -M a�SE:B�@pp���AGpL��r�m@all���*0a�OCB WA����"3 CNT0� T9DWroO0a�larm�ˀm0d� t�M�"0�2|� 9o�Z@OME<�� ���E%  #1-�S�RE��M�st}0g�     5K�ANJI5no �MNS@�INISITALIZ'�3 E�f�we��6@�� dr�@ fp �"��SCII L��afails w|��SYSTE[��i��  � Mq��1QGro8�m �n�@vA����&��nx�0q��RWRI �OF Lk��� \gref"�
�up� de-rela�Q_d 03.�0SS�chőbetwe�4�IND ex 6ɰTPa�DO� �l� �ɰGigE��soperabi]l`p l,��Hc�B��@]�le�Q0c�flxz�Ð���O�S {����v4pfigi GLA�$�c2z�7H� lap�0�ASB� If��g�2 l\c�0��/�E�� EXCE	 㰁�P���i��� o0��Gd`]Ц�f<q�l lxt��EFal��#0�i�O�Y�n�CLOS��S[RNq1NT^�F��U��FqKP�ANIO' V7/ॠ1�{����DB �0���v��ED��DET|��'� �bF�NLI;NEb�BUG�T�:��C"RLIB��A���ABC JAR�KY@��� rkeMy�`IL���PR���N��ITGAR� D$�R �Er *�T��a�U�0��h�[��ZE V� TASK p.vr��P2" .�XfJ�srqn�S谥dIBP	c����B/��BUS.��UNN� j0-��{��cR'���LO�E�DIVS�CUL`s$cb����BW!���R~�W`P�����I�T(঱tʠ�OF��UNEXڠ+����p�FtE��SVE�MG3`NML 5�05� D*�CC_SAFE�P*� ���� PET��'P�`��F  !���IR(����c i S>� �K��K�H GU�NCHG��S�M�ECH��M��T�*�%p6u��tPOR�Y LEAK�J���SPEgD��2�V 74\GRI���Q�g��CTLN��TRe @�_�p ��6�EN'�IN���`���$���r��T3)�.i�STO�A�s�	L��͐X	���q��1Y� ��TO2�J �m��0F<�K����D)U�S��O��3	 9�J F�&���S?SVGN-1#I�N��RSRwQDAU�C@ޱ� �T6�g��� 3��]���BRKCTR8/"� �q\j5��_��Q�S�qINVJ0D ZO�Pݲ���s���г�Ui ɰ̒�a�D�UAL� J50�e�x�RVO117 AW�TH!Hr%�nN�247%�52��|�&aol ���R��(�at�Sd�cU���P,�LER��iԗQ0�ؖ  ST���M�d�Rǰt� \fosB�A�0Np�c�����{�U��ROP �2�b�pB��ITP�4M��b !AU�t c0< � plet9e�N@� z1^q�R635 (Ac�cuCal2kA���I) "�ǰ�1
a\�Ps��ǐ� b���0P򶲊���ig�\cbacul "A3p_ �1��ն����etaca��AT���PC�`�����;_p�.pc!Ɗ�<�:�circB����5�tl��Bɵ�:�f!m+�Ί�V�b�ɦ�~r�upfrm.����ⴊ�xed��Ί�N~�pedA�D �}b>�ptlibB�� �_�rt��	Ċ�a_\׊ۊ�6�fm�� ��oޢ�e��̆Ϙ���c�Ӳ�5�j>�����#tcȐ��	�r���ʸ�mm 1��T�sl�^0��T�mѡ�#�r�m3��ub Y�q�s3td}��pl;�&�cckv�=�r�vf������9�vi����Cul�`�0fp�q ��.f��� daq�; i Data A�cquisi��nB�
��T`��1��89��22 D�MCM RRS2�Z�75��9 3 �R710�o59�p5\?��T "��1 (D�T� nk@��������E Ƒ�ȵ��Ӹ�etdm�m ��ER����gxE��1�q\mo? ۳�=(G���[0(

�2�` ! �@�JMACRO��S�kip/Offs�e:�a��V�4o9<� &qR662����s�H�
 6Bq8�����9Z�43 �J77� 6�J783�o ��n�"vv�R5IKCBq?2 PTLC�Z�g R�3 (�s�, �������0�3�	зJԷ\sf�mnmc "MN�MC����ҹ�%mnf�FMC"Ѻ0�>� etmcr� ��8���� ,�[�Df� �  874\p'rdq>,jF0�ޢ�axisHPr�ocess Axwes e�rol^�PRA
�Dp� 56o J81j�59� 56o6� ���0w��690 98� [!I#DV�1��2(x2��2ont�0�
�����m2���?C��e�tis "ISD���9�� Fprax�RAM�P� D��d�efB�,�G�is_basicHB�@p޲{6�� 708�6��(�Acw:�������D
�/,��AMOX �� ��DvE��?;T��2>Pi� RAFM';�]�!PAM�V�W�Ee`�U�Q'
bU�75��.�ceNe� nt?erface^�1' 5&!54�K��b(Devam±�/�#����/<�Tane`"�DNEWE���btp_dnui �AI�_�s2�d_rsono���bAsfjN��bdv_arFvf�x0hpz�}w��hkH9x�stc��gApon1lGzv{�ff� �r���z�3{q'�Td>pchamp�r;e�p� ^597@7��	܀�4}0��mɁ��/�����lf�!�pcochmp]aMP&xB�� �mpev��8����pcs��Ye�S�� Macro�OD��16Q!)*��:$�2U"_,��Y�(PC ��$_;�������o��J�gegemQ@GEMSW�~ZG�gesndy��OD��ndda��S��s1yT�Kɓ�su^Ҋ�ĩ�n�m���L��  ���9:p'ѳ޲���spotplusp���`-�W�l�J��s��t[�׷p�key�ɰ�$��s�-Ѩ��m���\featu� 0FEAWD�o;olo�srn'!�2 p���a�As3��t�T.� (N. A.)��!e!�J#
 (j�,��oBIB��oD -�.�n��k9�"K��u[-�_����p� "PSE�qW����wop "sEЅ�&�:�J��� ���y�|��O8��5� �Rɺ���ɰ[��X� ������%�(
ҭ�q HL�0k�
�z�@a!�B�Q�"(g� Q�����]�'�.��� ��&���<�!ҝ_�#��tpJ�H�~Z��j��� ��y������2��e� �����Z����V��! %���=�]�͂��^2�@�iRV� on�Q$Yq͋JF0� 8ހ�`�	(^�dQueue���X\1�ʖ`�+~F1tpvtsn��YN&��ftpJ0v �RDV�	f��J1 iQ���v�en�^�kvstk��mp���btkclrq8���get�����r��`kacqk�XZ�strŬ�%�stl��~Z�np:!�`���q/�ڡ6!l�/Yr�m	c�N+v3�_� �����.v�/\jF��� �`Q�΋�ܒ�N50 (FR�A��+��͢fraparm��Ҁ�} =6�J643p:V��ELSE
#�V�AR $SGSY�SCFG.$�`_UNITS 2�D`G~°@�4Jgfr��4A�@FRL-��0ͅ �3ې���L�0NE�: �=�?@�8�v�9~Q�x304��;�BPR�SM~QA�5TX.�$VNUM_OLp��5��DJ507��~l� Functʂ�"qwAP��琉�3 �H�ƞ�kP9jQ�Q5 ձ� ��@jLJzBJ[ �6N�kAP����S>��"TPPR��\�QA�prnaSV��ZS��AS8Dj510U�-�`cr�`8 ���ʇ�DJR`jYȑH_  �Q �P�J6�a21��48�AAVM 5̕Q�b0 lB�`TU�P xbJ54s5 `b�`616����0VCAM ~9�CLIO b71�5 ���`gMSC8�
rP R`�\sSTYL� MNIN�`J6�28Q  �`NR�Ed�;@�`SCH ���9pDCSU M�ete�`ORSR� Ԃ�a04 kR�EIOC �a5.�`542�b9vpP@<�nP�a�`�R�`7�`��MASK 3Ho�.r7 �2�`OOCO :��r3� �p�b�p���r0X��a��`13\mn�a3?9 HRM"�q�q~��LCHK�u�OPLG B��a0�3 �q.�pHCR� Ob�pCpPosyi�`fP6 is[r�J554�òpDS�W�bM�D�pqR�a337 }Rjr0 �1�s�4 �R6�7��52�r5 �2�r7 1� P6���Regi��@T�uFRD�M�uSaq%�4�`9{30�uSNBA�u�SHLB̀\sf�"pM�NPI�S�PVC�J520v��TC�`"MNрoTMIL�IFV��PAC W�pTP�TXp6.%�TELN N Me��09m3UEC9K�b�`UFR�`���VCOR��VIPuLpq89qSXC�S��`VVF�J�TPy �q��R626l��u S�`Gސ�2�IGUI�C��P�GSt�\ŀH86�3�S�q�����q34:sŁ684���a��@b>�3 :B��1� T��96 .�+�E�51 y�q53̀3�b1 ���b1 �n�jr9 ���`VAsT ߲�q75 s�xF��`�sAWSMӞ�`TOP u�ŀRq52p���a80 
��ށXY q���0 \,b�`885�QXр�OLp}�"pE࠱t�p�`LCMD��EgTSS���6 �>V�CPE oZ1�gVRCd3
�NLH�h��001m2Ep���3 f��p��4 //165C��6l����7PR��008 �tB��9 -200��`U0�pF�1޲1	 ��޲2L"���p���޲4��5 \h�mp޲6 RBCF`�`ళ�fs�8 ������~�J�7 rbcfA�L�8\PC����"�32m0u�n�K��Rٰn�5 5EW�
n�9 z��4�0 kB��3 ��6|ݲ�`00iB/��I6�u��7�u��8 �0�������sU0�`�t� �1 05\rb��2 E���K���dj���5˰��60��a�HУ`:�63�jAF�_���F�7 ڱ݀H�a8�eHЋ��cU0���7�p��1u��8<u��9 73����&��D7� ��5t�W97 ��8U�1���2��1�1:���h���1np�"��8(�U=1��\pyl��,�p��v ��B�854���1V���D�4��im��1�<���>br�3pr�4@pGPr�6C B���цp��1��r��1�`͵155ض�157 �2��62 �S����1b��2$����1Π"�2����B6`�1<c�4� 7B�5 DR��8�_�B/��187 �uJ�8 06�9s0 rBn�1 (���202 0EW,�ѱ2^��2��90�U12�p�2��2 b��u4��2�a"RB����9\�U2�`w�l����4 60Mp��7�������b�s
5 ¿�3����pB"9 �3 ����`ڰR,:7 �2��V�2���5���2^��a^9����qr����n�5 ����5᥁"�8a�Ɂ}�5B���5����`!UA���� ��86 �+6 S�0��5�p�2<�#�529 �2^��b1P�5~�2�`���&P5��8"��5��u�!�5��ٵW544��5��R��P nB^z�c (4�����U5J�V�5��1�1^���%�����5 b2a1��gA��58W[82� rb��5N��E�5890r� 1�95 �"������ c8"a��|�L ���!�J"5|6��^!�6��B�"8�`#��+�58%�6B�AME�"�1 iC��622D�Bu�6V��d� 4��{84�`ANRSP�e/S� C�5 � �6� ��� \� �6�� �V� 3t��� �T20CA�R��8�� Hf� 1DH�� A�OE� �� ,[|�� �0\�� �!64K��ԓrA� ��1 (M-7�!/50T�[PM��P�Th:1�C�#Pe� ��3�0� 5`M75cT"� �D8p� �0�Gc� u�4��i1-7'10i�1� Skd�7�j�?6�:-HS, � �RN�@�UB�f<�X�=m75sA*A�6an���!/CB�B2.6A �0;A�CIB�A��2�QF1�UB2�21� /70�S� �4��A��Aj1�3p���8r#0 B2\m*A@�C��;bi"i1K�u"A�~AAU� imm7c�7��ZA@I�@�Df��A�D5*A�E� 0TkdR1�35Q1�"*�@�Q�1�QC)P�1*A�5�*A�EA�5B�4>\77
B7=Q�D�2�Q$BR�E7�C�D/qAHEE�W7�_|`jz@� 2�0�Ejc7�`�E
"l7�@7�A
1�E�V$~`�W2%Q�R9ї@0L_�#����"Aȉ��b��H3s=rA/2�R5nR4�74rNUpQ1ZU�A�s\m9
1M92L2�!F!^Y�ps� 2ci��-?�qhimQ�t  w043�C��p2�mQ�r�H_ �H2�0�Evr�QHsXBSt62�q`s����� �<�Pxq350_*A3#I)�2�d�u0�@� �'4TX�0�pa3i1A3sQ25�c��st�r�VR1%e�q0
��j1��O2  �A�UEiy�.�‐ �0dCh20$CXB79#A��ᓄM Q1]�~�� 9�Q��?PQ��qA!P vs� 5	15aU����?PŅ���ဝQ9A6�zS*�7�qb5�1p����Q��00P(��V7]u�aitE1���À�p?7� !?�z��r=bUQRB1PM=�Q�a9��H��QQ�25L��������Q��@L���8ܰ��y00\}ry�"R2BL�t�N  ��� �1Df��2�qeR�5���_b�3�X^]1m1lcqP1�a��E�Q� 5F����!5<���@M-16Q��  f���r��Q�e� ��8� PN�LT_�1��i1��9453��@�e�|�b1l>F1u *AY2�
��R8�Q����RJ�J3�D}T� 85
Qg�/0��*A!P@�*A�Ð𫿽�2ǿپ6t�6=Q���P�ȓ��� AQ�  g�*ASt]1^u�ajrI� B����~�|I�b��y&I�\m�Qb�I�uz��A�c3Apa9q� B6�S��S��m���}�8�5`N�N�  �(M���f1���6�����161��5�s`�SC��U��A�����5\set06c�����10�y�h8���a6��6��9r�2HS ���Er���W@}�a��I�lB���Y�ٖ�m�u�C��� �5�B��B��h`�F� ��X0���A:���C�M�B��AZ��@��4�6i� ���� e�O�-	�� �f1��F �ᱦ�1pF�Y	���T6HL3���U66~`���U�dU�9D20Lf0��Qv � ��fjq��N���� ��0v
� ��i	�	.��72lqQ2�������� \chng�move.V��d����@2l_ar f	�f~��6��� ���9C�Z���~���kr41 S���0��V��t�����U�p7nuqQ%�A]�,�V�1\�Qn�BJ�2W�EM!5�0��)�#:�64��F��e50S�\��0� =�PV���e�������E�����m7;shqQSH"U��)@��9�!A��(����� ,[��ॲTR1!��,�60e=�4F�����2��	 R-����� ������Ж��4���LSR�)"�!l�OA��Q�) %!� 16�
U/��2�"2��E�9p���2X� SA�/i��'�
7F�H �@!B�0��D���5V ��@2cVE��p��T�2�pt갖�1L~E�#ȚF�Q��9E�#De/��RT��59���	�A��EiR������9\7m20�20��+�-u�19r4�`�E1�= `O9`�1"ae��O2��_$W}am4�1�4�3�/d1c_std��1)�!�`_T��r�_ 4\jdg�a�q�PJ%! ~`-�r�+bgB��#Nc300�Y�5j�QpQb1�bq��vB��v25�U�����qm43� �Q<W�"Ps A��e���� t�i�P�W.��c�@FX.�e�kE14��44�~6\j4��443sj��r�j4up���\E19�h�PA�T�=:o�APf���coWo!\�2a���2A;_2��QW2��bF�(�V11�23`�`��X5�Ra21�!J*9�a:88J99X�l5�m1a첚��*���(85�&��� ����P6���R,!52&A����,fA9INfI50\u�z�OV
 �v��}E֖J���Y>� 16r�C�Y��;��1��L���Aq�&� �P1��vB)e�m������1p� �1D�f��27�F�KA�REL Use =S��FCTN��� J97�FA+�� (�Q޵�p%�)?�V�j9F?(�j�Rtk?208 "Km�6Q��y�j��iæPr�9��s#��v�krcfp�RCFt3���Q�¿kcctme�!M�E�g����6�mai�n�dV�� ��ru��kDº�c���o��L��J�dt�F ����.vrT�f������E%�!��5�FRj7%3B�K���UER�H�J�O  J�� (ڳF���F�q�Y�&T���p�F�z��19�tk vBr���V�h�9p�E�y�<�k������;�v���"CT��f�� ��)�
І��)�V	� 6���!��qFF��1 q���=�����O�?�$"����$��je��T?CP Aut�r�<�520 H5�J[53E193��9��+96�!8��9��	 n�B574��52�uJe�(�� Se%!�Y�����u��ma�Pqtool�ԕ��������conrel��Ftrol Re?liable�Rmv9CU!��H51���p�� a551e"<�CNRE¹�I�c�&��it�l\�sfutst "�UTա��"X�\u@��g@�i�6Q]V0�B$,Eѝ6A� �Q� )C���X��Yf�I�1�|6s@6i��T6AIU��vR�d�
$e%1��2�C58�E6���8�Pv�iV4OFH58�SOeJ� mvBM6E~O58�I�0�E�#+@ �&�F�0���F�P6a����)/++�</N)0�\tr1�����P �,[�ɶ�rmaski�msk�aA���Iky'd�h	A	�P�s�DisplayI�m�`v����J88G7 ("A��+Heůצprds��IϩǪ��h�0pl�2�R2Ƚ�:�Gt�@��PRD�TɈ�r�C�@Fm�8�D�Q�AscaҦ�� V<Q&��bVvbrl�eې@��^S��&5�Uf�j8710�yAl	��Uq���7�&��p�p��P^@�P�firmQ����Pp�2�=bk�6�r�3��6��otppl��PL���O�p<b�ac�q	��g 1J�U�d�J��gait_9e��Y�&��Qx���	�Shap��eration�0<��R67451j9:(`sGen�ms�42-f��r�p�5����2�rsgl�E��pp�G���qF�205p��5S���Ձ�retsdap�BP�O�\s�� "GCR�ö? ^�qngda�G��V��st2axU��A1a]��bad�_�>btputl/�&�|e���tplibB_��=�2.����5���gcird�v�slp���x�hex��v�rqe?�Ɵx�key��v�pm��x�us$�6�gcr��F���p���[�q27j92��v�ollismqS�k�9O�ݝ� (p#l.���t��p!o��A29$Fo8��cg7no~@�tptcls` �CLS�o�b�\�km�ai_
�s>�v�o�	�t�b���ӿ�E��H��6�1enu�501�[m��ut�ia|$calma�UR��CalMat�eT;R51%�i=1 ]@-��/V� ��Z��� �fq1�9 "K9�E�L����2m�C�LMTq�S#��et �LM3!} �F�c�nspQ�c���Oc_moq��� ��cc_e�����su���ޏ �_ �@�5�G�join�i�j��oX���&cWv	 ���N�sve��C�clm��&Ao# �|$find�e�0STD� ter Fi�LANG���R���
��n3��z0C3en���r,���� ��J����� ���K ��Ú�=���_Ӛ���r� "FNDRК� 3��f��tguid�䙃N�."��J�tq�� �������@������J����_�� ����c��	m�Z�~�\fndr.��n#>
B2p��Z�C�P Ma�����3�8A��� c��6� ( ���N�B�������� 2�$�81��m_���"ex�z5 �.Ӛ��c��bS���efQ��	���RBT;�OPTN �+#Q�*$�r *$��*$r*$%/s#C��d/.,P�/0*ʲDPN��$���$*��Gr�$k Exc��'IF�$MASK��%93 H5�%H�558�$548 H�$4-1�$��#1(�$�0 E�$��$�-b�$���!UPDT �B�4�b�4�2�49��0�4a�3�9j0"Mx�49�4  ��4<�4tpsh���4<�P�4- DQ� �3 �Q�4�R�4�pR%0�2�r�4.b
E\���5�Ax�4��3adq\�5K979":E�ajO? l "DQ^E^�3i�Dq ��4ҲO) ?R�? ��q�5��T��3rAq�O�Lst�5~��7p�5��REJ#�2�@av^Eͱ�F蠠�4��.�5y N|� �2il(in�4��31 JH1�2Q4�251ݠ�4rma	l� �3)�REo�Z_ �æOx����4��^F�?onorTf��7_ja��UZҒ4l�5rms�AU�Kkg���4�$HCd\�fͲ�eڱ�4�RE	M���4yݱ"u@�RE�R5932fO��47|Z��5lity,�Up��e"Dil\�5���o ��7987p�?�25 �3hk910 �3��FE�0=0P_>�Hl\mhm�5 ��qe�=$�^�
E�x�u�IAymptm�U0��BU��vste�y\ �3��me�b�DvI�[� Qu�:F�Ub�*_�
EL,�su��_ �Er��ox���4hGuse�E-�?�sn��������FE��,�box�����c݌,"� ������z��M��<g��pdspw)�	� �9���b���(��1���c��Y�R� � �>�P���W��������'�0ɵ�[���͂���  �� ,[@� ��A�bump�šf��B*�Box%��7Aǰ60�BBw�\��MC� (6�,f��t I�s� ST ��*��}B�����=w��"BBF
�>��`���)��\bb?k968 "�4��ω�bb�9va699����etbŠ��1X�����ed	�F�b�u�f� �sea""������'�\��,� ���b�ѽ�o6�H�
�x�$�f���!y�����Q[�! tpe�rr�fd� TP�l0o� Recov�,��3D��R64�2 � 0��C@}s�� N@��(U�rroč��yu2r��  �
  �����$$CLe� ��������������$z�_DI�GIT��������.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$j���+c:PROD�UCTM�0\PG/STKD��V&oho�zf99��D����$FEAT_�INDEX��xd���  �
�`ILECOM�P ;���#���`�cSETUPo2 <�e�b?�  N �a�c�_AP2BCK �1=�i  �)wh0?{%&c����Q�xe%�I �m���8��\� n����!���ȏW�� {��"���F�Տj��� w���/�ğS������ ���B�T��x���� ��=�үa������,� ��P�߯t������9� ο�o�ϓ�(�:�ɿ ^���Ϗϸ�G��� k� �ߡ�6���Z�l� �ϐ�ߴ���U���y� ���D���h��ߌ� ��-���Q������� ��@�R���v����)� ����_�����*�� N��r��7� �m�&�3\t�i
pP 2#p*.VRc�*��� /�ƗPC/1/F'R6:/].��/+T�`�/�/F%�/�,�`r/?�*.F��8?	H#&?e<x�/�?;STM �2��?�.K �?�=�iPendant? Panel�?;H�?@O�7.O�?y?�O:GIF�O�O�5�OpoO�O_:JPG _�J_�56_�O_�_�	�PANEL1.D	T�_�0�_�_�?O�_2�_So�WAo�_o�o�Z3qo�o�W�o�o�o)�Z4�o[�W�I��
TP�EINS.XML��0\���q�Custom T?oolbar	���PASSWOR�DyFRS:�\L�� %Pa�ssword Config���֏ e�Ϗ�B0���T�f� ���������O��s� �����>�͟b��[� ��'���K��򯁯� ��:�L�ۯp�����#� 5�ʿY��}��$ϳ� H�׿l�~�Ϣ�1��� ��g��ϋ� ߯���V� ��z�	�s߰�?���c� ��
��.��R�d��� ����;�M���q�� ����<���`������ %���I�������� 8����n���!� �W�{"�F �j|�/�S e��/�/T/� x//�/�/=/�/a/�/ ?�/,?�/P?�/�/�? ?�?9?�?�?o?O�? (O:O�?^O�?�O�O#O �OGO�OkO}O_�O6_ �O/_l_�O�__�_�_ U_�_y_o o�_Do�_ ho�_	o�o-o�oQo�o �o�o�o@R�ov ��;�_�� �*��N��G���� ��7�̏ޏm����&� 8�Ǐ\�돀��!��� E�ڟi�ӟ���4�ß X�j��������įS���w������B�#���$FILE_DG�BCK 1=���/���� ( �)
S�UMMARY.DyGL���MD:������Diag� Summary���Ϊ
CONSLOG�������D�ӱ�ConsoleO logE�ͫ���MEMCHECK�:�!ϯ���X�Me�mory Dat�a��ѧ�{)>��HADOW�ϣ����J���Shad�ow Chang�esM�'�-��)	FTP7Ϥ�3������Z�mmen�t TBD��ѧ0�=4)ETHERNET��������T�ӱEther�net \�figurationU��ؠ��DCSVRF��߽߫�����%��� verify� all��'�1P{Y���DIFF��p����[���%��diff]�������1R�9�K��� ����X��CH�GD������c��r����2ZAS�� ��GAD���k��z��FY3bI[�� �/"GAD���s/�����/*&UPDAT�ES.� �/��FORS:\�/�-Ա�Updates �List�/��PS�RBWLD.CM�(?���"<?�/Y�P�S_ROBOWEL��̯�?�?��?&� O-O�?QO�?uOOnO �O:O�O^O�O_�O)_ �OM___�O�__�_�_ H_�_l_o�_�_7o�_ [o�_lo�o o�oDo�o �ozo�o3E�oi �o���R�v ���A��e�w�� ��*���я`������ ���O�ޏs������ 8�͟\�����'��� K�]�쟁����4��� ۯj������5�įY� �}������B�׿� x�Ϝ�1���*�g��� ��Ϝ���P���t�	� ߪ�?���c�u�ߙ� (߽�L߶��߂��� (�M���q� ���6� ��Z������%���I� ��B�����2������h����$FIL�E_� PR� ���������MDONL�Y 1=.�� 
 ���q��� �������~% �I�m�2 ��h��!/�./ W/�{/
/�/�/@/�/ d/�/?�//?�/S?e? �/�??�?<?�?�?r? O�?+O=O�?aO�?�O �O&O�OJO�O�O�O_��O9_�OF_o_
VI�SBCKL6[�*.VDv_�_.POFR:\�_�^.P�Vision VD file�_ �O4oFo\_joT_�oo �o�oSo�owo�o B�of�o�+� ������+�P� �t������9�Ώ]� 򏁏��(���L�^�� �����5���ܟk� � ��$�6�şZ��~������
MR_GR�P 1>.L~��C4  B����	 W������*u����RHB ��2 ���� ��� ���B�����Z�l� ��C���D�������Ŀ���K�bYJ��_�I��Tx��F�5UP��2]���ֿ E���G�7E�&T�;�Kv:]�S@q��@���@�%U�f�@�)��@�*λ� F@ ��������J��NJk��H9�Hu���F!��IP�s��?����(�9��<9�8�96C'6<,6\b��+�&Ϡ(�a�L߅�p�A��A��߲�v���r����� �
�C�.�@�y�d�� ��������������?�Z�lϖ�BH��� �Ζ�������
�0�PS@�P�Waf��ܿ� �B���</ ��@�33:��q.�gN�UUU��U��q	>u.�?!rX��	��-=[z�=��̽=V6<��=�=�=�$q�����@8��i7G��8��D�8@9!�7�:�����D�@ D��g Cϥ��C������'/0-��P/� ���/N��/r��/���/ �??;?&?_?J?\? �?�?�?�?�?�?O�? O7O"O[OFOOjO�O �O�O�O�гߵ��O$_ �OH_3_l_W_�_{_�_ �_�_�_�_o�_2oo VohoSo�owo�o�i�� �o�o�o��);�o _J�j���� ���%��5�[�F� �j�����Ǐ���֏ �!��E�0�i�{�B/ ��f/�/�/�/���/� �/A�\�e�P���t��� �����ί��+�� O�:�s�^�p�����Ϳ ���ܿ� ��OH�� o�
ϓ�~ϷϢ����� �����5� �Y�D�}� hߍ߳ߞ��������o �1�C�U�y��߉� ������������-� �Q�<�u�`������� ��������;& _J\������� ���ڟ�F�j 4�������� �!//1/W/B/{/f/ �/�/�/�/�/�/�/? ?A?,?e?,φ?P�q? �?�?�?�?O�?+OO OO:OLO�OpO�O�O�O �O�O�O_'__K_� o_�_�_�_l��_0_�_ �_�_#o
oGo.okoVo ho�o�o�o�o�o�o �oC.gR�v �����	��� <�`�*<��`�� ���ޏ��)��M� 8�q�\�������˟�� �ڟ���7�"�[�F� X���|���|?֯�?�� ���3��W�B�{�f� ����ÿ�������� �A�,�e�P�uϛ�b_ �����Ϫ_��߀�=� (�a�s�Zߗ�~߻ߦ� ������� �9�$�]� H��l�������� ����#��G�Y� �B� ������z�������
 ԏ:�C.gRd� �����	� ?*cN�r�� ���/̯&/�M/ �q/\/�/�/�/�/�/ �/�/?�/7?"?4?m? X?�?|?�?�?�?�?�� O!O3O��WOiO�?�O xO�O�O�O�O�O_�O /__S_>_P_�_t_�_ �_�_�_�_�_o+oo Oo:oso^o�o�op��o �� ��$�� o�o�~���� ���5� �Y�D�}� h�������׏��� �
�C�.�/v�<��� 8������П���� ?�*�c�N���r����� ���̯��)��?9� _�q���JO�����ݿ ȿ��%�7��[�F� �jϣώ��ϲ����� ��!��E�0�i�T�y� �ߊ��߮��߮o�o� �o>�t�>��b �����������+�� O�:�L���p������� ������'K6 oZ�Z�|�~��� ��5 YDi �z������ /
//U/@/y/@��/ �/�/�/���/^/?? ?Q?8?u?\?�?�?�? �?�?�?�?OO;O&O 8OqO\O�O�O�O�O�O��O�O_�O7_��$�FNO ����VQ��
F0fQ kP oFLAG8�(LR�RM_CHKTY/P  WP��^P��WP�{QOM��P_MIN�P�����P�  X�NPSSB_CFG� ?VU ��_���S o�oIUTP_DEF�_OW  �|�R&hIRCOM�P�8o�$GENOV�RD_DO�V��6�flTHR�V dz�edkd_ENBWo� k`RAVC_?GRP 1@�WCa X"_�o_1 U<y�r�� ���	��-��=� c�J���n�������� ȏ����;�"�_�F��X���ibROU�`F\VX�P�&�|<b&�8�?���埘������� � D?�јs���@@g�B�7�p�)�ԙ\���`SMT�cG�m�M���� �LQHO7STC�R1H���P���at�SM���f�\����	127.0��1��  e��ٿ� ����ǿ@�R�d�v����0�*�	anonymous������������[�� � �����r����� �ߺ�����-���&� 8�[�I�π���� ��1�C��W�y� ��`�r������ߺ��� ����%�c�u�J\ n�������� �M�"4FX��i ������7/ /0/B/T/���m/ ��/�/�/??,? �/P?b?t?�?�/�?� �?�?�?OOe/w/�/ �/�?�O�/�O�O�O�O �O=?_$_6_H_kOY_ �?�_�_�_�_�_'O9O KO]O__Do�Ohozo�o �o�o�O�o�o�o
 ?o}_Rdv���_ �_oo!�Uo*�<� N�`�r��o������̏ ޏ�?Q&�8�J�\����>�ENT 1I��� P!􏪟  ����՟ğ�� �����A��M�(�v� ��^�����㯦��ʯ +�� �a�$���H��� l�Ϳ�����ƿ'�� K��o�2�hϥϔ��� ���ϰ�������F� k�.ߏ�R߳�v��ߚ� �߾���1���U��y��<�QUICC0 ��b�t����1�����%���2&���u��!ROUTER�v�R�d���!PC�JOG����!�192.168.�0.10��w�NA�ME !��!�ROBOTp�S_CFG 1H��� �A�uto-star�ted�tFTP�������  2D��hz� ���U��
// ./�v���/�� �/�/�/�/�/�!?3? E?W?i?�/?�?�?�? �?�?�?���AO�? eO�/�O�O�O�O�?�O �O__+_NO�OJ_s_ �_�_�_�_
OO.Oo B_'ovOKo]ooo�oP_ >o�o�o�o�oo�o 5GYk}�_�_�_ ��8o��1�C� U�$y��������ӏ f���	��-�?��� ��Ə���ϟ�� ���;�M�_�q��� .�(���˯ݯ��P� b�t�����m������� ��ǿٿ�����!�3� E�h��{ύϟϱ��� �$�6�H�J�/�~�S� e�w߉ߛ�jϿ����� ���*߬�=�O�a�s����YT_ERR �J5
���PDU�SIZ  ��^�J����>��WR�D ?t�� � guest}��%�7�I�[��m�$SCDMNG�RP 2Kt������V$��K�� 	P0�1.14 8�� _  y�����B    �;����� ���������
 �������������~����C.�gR|���  �i  �  k
�������� �+�������_
���l .r+���"�l��� m
d������__GROU��L�� �	����0�7EQUPD  �	պ�J�TY�a ����TTP�_AUTH 1M��� <!iP�endany���6�Y!KAR�EL:*��
-�KC///A/ V�ISION SE!TT�/v/�"�/ �/�/#�/�/
??Q?�(?:?�?^?p>�CTRL N����5��
�FFF�9E3�?�FR�S:DEFAUL�T�<FANU�C Web Se/rver�:
��� ��<kO}O�O�O�O�O���WR_CONF�IG O�� ��?��IDL_C_PU_PC@�sB��7P�BHU�MIN(\��<TGNR_IO�������PNPT_SIM�_DOmVw[TPMODNTOLmV} �]_PRTY�X�7RTOLNK 1P����_o!o3o�EoWoio�RMAST�ElP��R�O_C3FG�o�iUO��o>�bCYCLE�o�d�@_ASG 1Q����
 ko,> Pbt����������sk�bNU�M����K@�`IP�CH�o��`RTRY_CN@oR��b�SCRN����Q�b�� �b�`�bR����Տ��$J23_DSP_EN	�����OBPR�OC�U�iJOG�P1SY@��8��?�!�T�!�?>*�POSRE�zV?KANJI_�`��o_�� ��T�L�6x͕����CL_LGP�<�_���EYLOGWGIN�`����LANGUAGgE YF7RDY w���LG��U�?V⧈�x� ���j��=P��'0����$ NMC:�\RSCH\00�\��LN_DISP V��
���������OC�R.RDz�VTA{�OGBOOK W
{��i��ii��X����� ǿٿ�����"��6	h�����e��?�G_BUFF K1X�]��2	� �ϸ���������� �!�N�E�W߄�{ߍ� �߱�����������J���DCS }Zr� =���� ^�+�ZE��������a��IO 1[
{ ُ!� �!�1�C� U�i�y����������� ����	-AQc�u�������E^fPTM  �d�2 /ASew�� �����//+/ =/O/a/s/�/�/���SEV����TYP�/??y͒�RS@"��×��FL 1\
������?�?�?�?�?�?L�?/?TP6��"}>�NGNAM�ե�U`�UPS��G�I}�𑪅mA_L�OAD�G %��%DF_MO�TN���O�@MAXUALRM<��J� �@sA�Q����WS �
�@C �]m�-_���M�P2�7�^
{ �Z��	�!P�+ʠ1�;_/��Rr�W�_�WU�W�_��R	o �_o?o"ocoNoso�o �o�o�o�o�o�o�o ;&Kq\�x� ������#�I� 4�m�P���|���Ǐ�� �֏��!��E�(�i� T�f�����ß��ӟ�� �� �A�,�>�w�Z� ������ѯ����د� ��O�2�s�^����� ��Ϳ���ܿ�'��B�D_LDXDIS�AX@	��MEMO�_APR@E ?�+
 � *�~� �Ϣϴ����������@�ISC 1_�+ ��IߨT��Q�c� Ϝ߇��ߧ�����w� ���>�)�b�t�[�� ��{���������� :���I�[�/������ ������o�����6! ZlS��s� ���2�AS '�w����g���.//R/d/�_MSTR `�-~w%SCD 1am��L/�/H/�/�/?�/ 2??/?h?S?�?w?�? �?�?�?�?
O�?.OO RO=OvOaO�O�O�O�O �O�O�O__<_'_L_ r_]_�_�_�_�_�_�_ o�_�_8o#o\oGo�o ko�o�o�o�o�o�o�o "F1jUg� �������� B�-�f�Q���u������ҏh/MKCFG �b�-㏕"LT�ARM_��cL�;� σQ�|N�<�METPUI��ǂ���)NDS?P_CMNTh��8�|�  d�.���ς�ҟܔ|�PO�SCF����PS�TOL 1e'�4=@�<#�
5�́ 5�E�S�1�S�U�g��� ����߯��ӯ���	� K�-�?���c�u������|�SING_CH�K  ��;�ODAQ,�f��Ç��DEV 	L�	�MC:!�HSI�ZEh��-��TA�SK %6�%$�12345678�9 �Ϡ��TRI�G 1g�+ l6�%���ǃ����ό8�p�YP[� ��E�M_INF 1h�3� `�)AT&FV0�E0"ߙ�)��E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ������H�� ���A���AI�q� ,��|���� ��� �ߵ�����J���n��� ����W����������� "����X��/�� ��e������0 �T;x�=�a s��/�,/c=/ b/�/A/�/�/�/�/ ��?���^?p? #/�?�/�?s?}/�?�? O�?6OHO�/lO?1? C?U?�Oy?�O�O3O _ �?D_�OU_z_a_�_玿ONITOR��G� ?5�   	?EXEC1Ƀ�RU2�X3�X4�X5�XT���V7�X8�X9Ƀ�RhBLd�RLd�RLd �RLd
bLdbLd"bLd@.bLd:bLdFbLc2ShU2_h2kh2wh2�hU2�h2�h2�h2�hU2�h3Sh3_h3�R��R_GRP_SOV 1in���(�����C?BPP��A4�>%���gY�>rﳌ�x�_D=R^��P�L_NAME �!6��p�!D�efault P�ersonali�ty (from� FD) �RR�2eq 1j)TU�X)TX��q��X dϏ8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|������2'�П�����@*�<�N�`�r��<�� ������ү������,�>�P�b� �Rdr �1o�y �\�,� �3���� �@D�  ��?�ĸ���?䰺��A'�6����;�	�lʲ	 ��xJ������ �<w �"�� �(���pK�K ���K=*�J����J���JV�`��Z�����r���́p@j�@T;;f���f��ұ�]�l��I���������������b��3��´  ��`�>����b����z��ꜞ����Jm��
� B�H�˱]���q��	� p�  �P�pQ�p��p|  Ъ�g���c�	'� � ���I� �  �����:�È~
�È=���"��nÿ�	�ВI  ?�n @B�c���\��ۤ��q�y��o�N���  '������@2��@Ǔ����/�C���C�C�@ C�������
��A�W�@<�P�JR�
h�B�b�A�Єj�����:��Dz۩��߹������j��( �� -��C���'�7�����q�Y������ �?�ff� ��gy ����o�:a�:�
>+�  PƱj�(����7	�ü�|�?����x�Z�p<
6b<�߈;܍�<��ê<� <�#&Jσ�AI�ɳ�+���?fff?�I�?&�k�@�.���J<?�`�q�.�˴fɺ� /��5/����j/U/ �/y/�/�/�/�/�/?0�/0?q��F�? l??�?/�?+)�?�?~�E�� E�I�?G+� F��? )O�?9O_OJO�OnO�Of�BL޳B�?_h� .��O�O��%_�OL_�? m_�?�__�_�_�_�_��
�h�Îg>��_Co�_goRodo�o�GA�ds�q��C�o�o�o|���A�$]Hq���D���pC���pC!HmZZ7t���6q�q���ܶN'�3A��A�AR1AO��^?�$�?��K/�±
=���>����3�?W
=�#�W���e��9������{����<�����(�B�u���=B0������	L���H�F�G����G��H�U�`E���C�+����I#�I���HD�F���E��RC��j=��
I���@H�!H��( E<YD0q�$��H�3�l� W���{��������՟ ���2��V�A�z��� w�����ԯ������ ��R�=�v�a����� �������߿��<� '�`�Kτ�oρϺϥ� �������&��J�\� G߀�kߤߏ��߳��� ����"��F�1�j�U� ��y���������� ��0��T�?�Q�����(���3/E�y���u����<��q3�8�����q4Mgs&�IB+2D�a���{�^^	�@�����uP2	P7Q4_A��M00bt��R��`����/   �/�b/P/�/t/�/  *a)_3/�/�/�%1a?�/?;?M?_?q?  �?�/�?�?��?�?O 2 F;�$�vGb�/�Aa��@�a�`�qC��C�@�o�Ot���KF�� DzH@�� F�P D���O�O�ys<O!_3_E_�W_i_s?���@U@pZ�422�!2~
  p_�_�_�_	oo-o?o Qocouo�o�o�o�o��Q ��+��1���$MSKCF�MAP  �5?� �6�Q��Q"~�cONREL7  
q3��bEXCFENB�?w
s1uXqFNC�_QtJOGOVLKIM?wdIpMrd�bWKEY?w�u�bWRUN�|�u�bSFSPDTY�xavJu3sSIGN?>QtT1MOT�Nq��b_CE_GRoP 1p�5s\r���j�����T�� ⏙������<��`� �U���M���̟��� ���&�ݟJ��C��� 7�������گ��������4�V�`TCOM_CFG 1q}��Vp�����
P�_/ARC_\r
jyUAP_CPL���ntNOCHECK� ?{  	r��1�C�U�g� yϋϝϯ����������	��({NO_WA�IT_L�	uM�NMTX�r{�[m�o_ERRY�2sy3� &��������r�c� ��T_�MO��t��,  �$�k�3�PAR�AM��u{��	�[���u?�� =�9@345678901��&���E�W� 3�c�����{������������=��UM_RSPAC�E �Vv��$ODRDSP���jx�OFFSET_C�ARTܿ�DIS���PEN_FI�LE� �q��c֮�O�PTION_IO���PWORK kv_�ms � P(�R�Q
�j.j�	 ��Hj&6$�� RG_DSBL'  �5Js�\���RIENTTO>p9!C��PqfA�� UT_SIM_ED
r�b� V� ?LCT ww�b�c��U)+$_PEX9E�d&RATp �v�ju�p��2X�j)T�UX)TX�##X d-�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO-O?O�H2�/oO�O�O �O�O�O�O�O�O_]�<^O;_M___q_�_�_ �_�_�_�_�_o����X�OU[�o(��_�(���$o�, ��IpB`� @D�  Ua?��[cAa?p]a]�D�WcUa쪋l;�	�lmb�`�x7J�`�p����a�< ���`� ��b��H(���H3k7HS�M5G�22G�?��Gp
��
�ƨ��'|��CR�>�>q�GsuaT��3���  �4spBpyr  ]o��*SB_����=j]��t�q� ��rna �,��~�6  ��UPQ�|N��M�,k���	'�� � ��I�� �  ��%�=��ͭ����ba	���I  �n @��~����p�������N	 W�  '!o�:q:�pC	 C�@@sBq��|��� m�
�T!�h@ߐ�n��$��*�B	 �A����p� �-�qbz ��P��t�_�������( �� -��恊�n�ڥD[A]Ѻ�b4�'!5�~(p �?�ff� ��
����OZ�R�*�85�z���>΁  Pia��(5���@����ک�a�c�dF#?˙�5�x��*�<
�6b<߈;����<�ê<�? <�&�o&ς)�A�lcΐI�*�?offf?�?&c�ޒ�@�.uJ<?�`��Yђ ^�nd��]e��[g��G� �d<����1��U�@� y�dߝ߯ߚ����߼� 	���-������&��~"�E�� E��?G+� Fþ��� ��������&��J�(5��bB��AT�8� ђ��0�6���>���J� n�7��[m��0��h��1��>�M�I
�@��A�[���C-�)��?Ƀ��� /�Y���Jp��vav`CH�/������}!@�I�Y�'�3A��A�AR1A�O�^?�$�?�����±
=�ç>����3�W
=�#�����+e��ܒ������{����<���.(�B��u��=B0�������	��*H�F�G����G��H��U`E���C��+�-I#�I���HD�F���E��RC��j=U>
I���@H�!H��( E<YD0/�?�?�?�?�? O�?3OOWOBOTO�O xO�O�O�O�O�O�O_ /__S_>_w_b_�_�_ �_�_�_�_�_oo=o (oaoLo�o�o�o�o�o �o�o�o'$] H�l����� ��#��G�2�k�V� ��z���ŏ���ԏ� ��1��U�g�R���v� ����ӟ�������-�:�(���������a����xQ�c�,!3�8�}�<��,!4Mgs�����ɢIB+կ篴a?���{����A�/�e�S���w��P!�P�������7�`�ӯ�ϑ�R9��Kτ�oχϓϥ�  ���χ����)�� M������z���{߉�����ߒߤ�������  )�G�q��_���2 wF�$�&Gb����n�[ZjM!C��s�@j/�A�S�=�F�� Dz���� F�P D��W����)������������x?��ͫ@@
9�=��=��=��
 v����� ��*<N`ܷ*P ���˨��1��$PARA�M_MENU ?�-�� � DEF�PULSEl	�WAITTMOU�T�RCV� �SHELL_�WRK.$CUR�_STYL��,OPT�/PT�B./("C�R_DECSN���,y/ �/�/�/�/�/�/?	? ?-?V?Q?c?u?�?��USE_PROG %�%�?�?�3CCR�����7�_HOST !F�!�44O�:T̰�?PCO)ARC�O�;_TIME�XB��  �GDEB�UGV@��3GINP_FLMSK�O��IT`��O�EPGA�P �L��#[CH��O�HTYPE����?�?�_�_�_�_ �_oo'o9obo]ooo �o�o�o�o�o�o�o�o :5GY�}� ���������1�Z��EWORD �?	7]	RS�`�	PNS��$��JOE!>�T�Es@WVTRACE�CTL 1x-�]� ������ɆDT Q�y-���D 7� ��,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�T�(� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ j��_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�_����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v��������//"#�$PGT�RACELEN � #!  ���" �8&_�UP z��e�g!o S!h �8!_CFG {Fg%Q#"!x!�$�J �#|"DEFSP/D |�,!!J ��8 IN TR�L }�-" 8��%�!PE_CON�FI� ~g%��g!�$�%�$L�ID�#�-74G�RP 1�7Q!��#!A ����&ff"!A+33�D�� D]� ?CÀ A@+6�!�" d�$�9�9*1*0?� 	 +9�(8�&�"�? ´	C�?�;B@3AO�?OIO�3OmO"!>�T?��
5�O�O�N�O �=��=#�
 �O_�O_J_5_n_Y_��O}_�_y_�_�_�_ G Dzco" 
o Bo�_Roxoco�o�o�o �o�o�o�o>)�bM��;
V7�.10beta1��$  A��E�rӻ�A �" �p?!G��q>����r��0�q{�ͻqBQ��q�A\�p�q�4�q�p
�"�BȔ2�D�V��h�w��p�?�?)2 {ȏw�׏���4� �1�j�U���y����� ֟������0��T� ?�x�c�������ү�� ��!o�,�ۯP�;�M� ��q�����ο���ݿ �(��L�7�p�+9��sF@ �ɣͷ� ��g%������+�!6 I�[߆������ߵߠ� ��������!��E�0� B�{�f�������� �����A�,�e�P� ��t���������� ��=(aL^� ������' 9$]�Ϛ��ϖ� ������/<�5/`� r߄ߖߏ/>�/�/�/ �/�/?�/1??U?@? R?�?v?�?�?�?�?�? �?O-OOQO<OuO`O �O�O�O�O���O_�O )__M_8_q_\_n_�_ �_�_�_�_�_o�_7o Iot���o�o�� �o�o�o(/!L/^/p/ �/{*o����� ����A�,�e�P� b����������Ώ� �+�=�(�a�L���p� �����Oߟ񟠟� � 9�$�]�H���l�~��� ��ۯƯ���#�No`o ro�on��o�o�o�oԿ ���8J\ng� ���vϯϚ������� 	���-��Q�<�u�`� r߫ߖ��ߺ������ �;�M�8�q�\���� ����z������%�� I�4�m�X���|����� ������:�L�^��� Z���������� �$�6�H�Sw b������� //=/(/a/L/�/p/ �/�/�/�/�/?�/'? ?K?]?H?�?��?�? f?�?�?�?O�?5O O YODO}OhO�O�O�O�O �O�O&8J4_F_� ���_�_��_�_ "4-o�O*ocoNo�o ro�o�o�o�o�o�o )M8q\�� �������7� "�[�m��?����R�Ǐ ���֏�!��E�0� i�T���x�������� _$_V_ �2�l_~_�_������R�$PLI�D_KNOW_M�  �T������SV ��U͠�U��
��.�ǟR��=�O�����mӣM_?GRP 1��!`U0u��T@ٰo�
ҵ�
���Pзj� �`���!�J�_�W� i�{ύϟϱ�������X��߱�MR�����1T��s�w� s��� �޴߯߅��ߩ߻��� ��A���'���� �����������=� ��#���������}�������S��ST��1W 1��U# ���;0�_ A .�� ,>Pb���� ����3(i L^p������2*���	<-/3/)/;/M/�4f/x/�/�/5 �/�/�/�/6??(?:?7S?e?w?�?�8�?�?�?�?M_AD  d#�`PARNUM  w�%OWSCH?J ME
�Gp`A�Iͣ�EUPD`O�rE
a�OT_CM�P_��B@�P@'�˥TER_CHK'U��˪?R$_6[�RSl�¯��_MO�A@�_�U_�_RE_R/ES_G �� >�oo8o+o\oOo�o so�o�o�o�o�o�o�o�W �\�_%�U e Baf�S� �� ��S0����SR0 ��#��S�0>�]�b���S�0}������RV �1�����rB@c]���t�(@c\�����D@c[��$���RTHR_�INRl�DA��˥d�,�MASS9� Z�M�MN8�k�MON�_QUEUE a���˦��x� RDNPUbQN{�P[���END���_ڙEX1E�ڕ�@BE�ʟ>��OPTIOǗ�[���PROGRAM7 %��%��ۏ��O��TASK_I�AD0�OCFG ኞ�tO��ŠDATuA���Ϋ@��27�>�P�b�t���,� ����ɿۿ�����#�x5�G���INFOU���������ϭϿ� ��������+�=�O� a�s߅ߗߩ߻���������^�jč� �yġ?PDIT �ίc���WERF�L
��
RGADoJ �n�A��¹�?����@���IOORITY{�QV���MPDSPH������Uz����OTO�Ey�1�R� (/!AF4�E�P]�~��!tcph�>��!ud��!icm��ݏ6�XY_ȡ�R�=�ۡ)� *+/ ۠�W:F �j����� �%7[B�=*��PORT#�BC�۠����_C?ARTREP
�R�> SKSTAz��Z�SSAV���n�	�2500H86A3���r�$!�R����q�n�}/x�/�'� URGE��B��rYWF� DO{�rUVWV��$�A��WRUP_DEL�AY �R��$RO_HOTk��%O�]?�$R_NORM�ALk�L?�?p6SE�MI?�?�?3AQS�KIP!�n�l#x 	1/+O+ O ROdOvO9Hn��O�G�O �O�O�O�O_�O_D_ V_h_._�_z_�_�_�_ �_�_
o�_.o@oRoo vodo�o�o�o�o�o�o �o*<Lr`���n��$RCgVTM�����p�DCR!�L���qB��C*J��C$�>�$� >5>�;���04M¹�O���ǃ��������~��9On�Y�<
�6b<߈;����>u.�??!<�&{�b� ˏݏ��8�����,� >�P�b�t��������� Ο���ݟ��:�%� 7�p�S������ʯܯ � ��$�6�H�Z�l� ~�������ƿ���տ ���2�D�'�h�zϽ� �ϰ���������
�� .�@�R�d�Oψߚ߅� �ߩ���������<� N��r������� ������&�8�#�\� G�����}��������� ��S�4FXj| ������� ��0T?x�u ����'//,/ >/P/b/t/�/�/�/�/ �/�/�?�/(??L? 7?p?�?e?�?�?��? �? OO$O6OHOZOlO ~O�O�O�?�?�O�O�O �O __D_V_9_z_�_ �?�_�_�_�_�_
oo�.o@oRodovo�X�qG�N_ATC 1��� AT�&FV0E/� �ATDP/6/�9/2/9�hA�TA�n,A�T%G1%B96}0/�+++�o�,�aH,�qIO�_TYPE  �u�sn_�oREFPOS1 1�P{� x�o�X h_�d_����� K�6�o�
���.���R�x���{{2 1�P{���؏V�ԏz����q3 1��$�6��p��ٟ���S4 1�����˟���n�|��%�S5 1�<��N�`�����<���S6 1�ѯ���/�𭿘�ѿO�S7 1�f�x���ĿB�-�f�>�S8 1������Y�������y�SM�ASK 1�P � 
9�G��XNO�M���a~߈ӁqMOTE  h�~t��_CFG �������рrPL_RA�NG�ћQ��POW_ER ��e����SM_DRYP_RG %i�%���J��TART ��
�X�UME_P�RO'�9��~t_E�XEC_ENB � �e��GSPD�������c��TDB����RM��MT�_!�T���`O�BOT_NAME� i���iO�B_ORD_NU�M ?
�\q�H863  a�T��������b�PC_TIMEO�UT�� x�`S2�32��1��k �LTEACH PENDAN ��ǅ�}���`�Maintena�nce ConsțR}�m
"{�dKCL/Cg��Z ���n� No Use}�	���*NPO��х����(CH_�L�������	��mMAVAILȰ�{��ՙ�SPACE1 2��| d��(>���&���p��M,8�?�ep/eT/ �/�/�/�/�W//,/ >/�/b/�/v?�?Z?�/ �?�9�e�a�=??,? >?�?b?�?vO�OZO�?��O�O�Os�2� /O*O<O�O`O�O�_��_u_�_�_�_�_[3 _#_5_G_Y_o}_�_ �o�o�o�o�o[4.o@oRodovo$�o �o����"�	�7�[5K]o��A� ���	�̏�?�&�T�[6h�z������� ^�ԏ���&��;�\�C�q�[7�������� ͟{���"�C��X�y�`���[8����Ư دꯘ��0�?�`�#��uϖ�}ϫ�[G ��i� �ϋ
G� ����$�6� H�Z�l�~ߐ��8 ǳ�@����߈��d(� ��M�_�q���� ��������?���2� %�7�e�w��������� �����������!�R E�W�����������?Q; `�� @0�@�ߖrz	�V_ �����
/L/^/ |/2/d/�/�/�/�/�/ �/?�/�/�/*?l?~? �?R?�?�?�?�?�?�?�?2O�?
��O[�_MODE  ��˝IS ���vO,*ϲ�O-_���	M_v_#dCWO�RK_AD�Mx{q�%aR  ���ϰ�P{_�P_INOTVAL�@����J�R_OPTION��V �EBpVA�T_GRP 2�����(y_Ho �e_vo�o�o Yo�o�o�o�o�o* <�bOoNDpw� �����	��� ?�Q�c�u�����/��� ϏᏣ����)�;��� _�q���������O�ɟ ���՟7�I�[�m� /�������ǯٯ믁� �!�3���C�i�{��� O���ÿտ���ϡ� /�A�S�e�'ωϛϭ� oρ�������+�=� ��a�s߅�Gߕ߻��� �ߡ���'�9�K�]� �߁����y����������5�G�Y��E��$SCAN_TI�M�AYuew�R ��(�#((��<0.aJaPaP
Tq>��Q��o����V�OO2/$��:	d/JaR��WY��^���^R�^	r  P��� �  8��P�	�D��GYk}�� ������Qp/@/R//)P;�o\T��Q�pg-�t�_�DiKT��[  � lv%������/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OWW�#�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_olO~O d+No`oro�o�o�o�o �o�o�o&8J \n������u�  0�"0g�/� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q�����$o��˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�����Do ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������w
�  58�J�\�n߀� �ߜկ���������	� �-�?�Q�c�u������ ��-�� ��� �2�D�V�h�z���������������v���& ���%	12345�678�" 	�
�/� `r�������� (:L^p�� ����� //$/ 6/H/Z/l/~/��/�/ �/�/�/�/? ?2?D? V?h?�/�?�?�?�?�? �?�?
OO.O@Oo?dO vO�O�O�O�O�O�O�O __*_YON_`_r_�_ �_�_�_�_�_�_oo C_8oJo\ono�o�o�o �o�o�o�oo"4 FXj|���������	��s�3�E�W�{�Cz � Bp��   ��2���z�$S�CR_GRP 1��(�U8(�\�x^ @�  �	!�	 ׃���"� $� ��-��+��R�nw����D~������#����O����M-10iA 78909905 Ŗ~5 M61C >P4��Jׁ
� ���0�����#�1�	"�z�������4¯Ҭ ���c� ��O�8�J��� ����!�����ֿ��B�y�������r��A��$�  @���<� �R�?��d���H�y�u�O���F@ F�`�§�ʿ�϶� ������%��I�4�m� �<�l߃ߕߧ߹�B���\����1�� U�@�R��v����� �������;���*<=�
F���?�d�<��>7�����@��:��� B����ЗЙ���EL_D�EFAULT  ������B�MIPOWERFL  �x$1 WFDO� $��ERVE�NT 1������"�pL!D?UM_EIP��8���j!AF_I�NE �=�!FIT���!���4 ��[!�RPC_MAIN�\>�J�nVI�Sw=���!�TP�PU��	d��?/!
PMON?_PROXY@/�Ae./�/"Y/�fz/��/!RDM_S�RV�/�	g�/#?!#R C?�h?o?K!
pM�/�i^?��?!RLSYN�C�?8�8�?O!�ROS�.L�4 �?SO"wO�#DOVO�O �O�O�O�O_�O1_�O U__._@_�_d_v_�_ �_�_�_o�_?ooco�iICE_KL �?%y (%SVCPRG1ho 8��e���o�m3�o�o"�`4 �`5(-"�`6PU�`7x}��`���l9��{ �d:?��a�o��a�o E��a�om��a���a B���aj叟a�� �a�5��a�]��a� ���a3����a[�՟�a �����a��%��aӏM� �a��u��a#����aK� ů�as���a��mob �`�o�`8�}�w����� ��ɿ���ؿ���5� G�2�k�VϏ�zϳϞ� ���������1��U� @�y�dߝ߯ߚ��߾� ������?�*�Q�u� `���������� ��;�&�_�J���n������������sj_�DEV y	��MC:�ջ_OUT"�,REC 1q�Z� d   w 	�    ��@��� ���A�����
 �PSD#O6 r��O� ��� �� `�� ��Z�{� �� �*�  +X- � I- �- !- �� �X�YZ�PS�J;4 �?j  (�  Q� ��R ���� E- � b�/e/�l4H�/��� X� (�,/>/P/�/�/�""J4� =�!� � ؀  ?"S1��Z'!�/���("- ��\?�?$=�=�?�? �?"OOFO4OjO|O^O �O�O�O�O�O�O�O_  __T_B_x_f_�_�_ �_�_�_�_�_ooo Po>oto�oho�o�o�o �o�o�o(
L:�\�p���w ,����4�"�X� F�|���p�����֏ď ����0��@�f�T� ��x�����ҟ�Ɵ� ��,��<�b�P���h� z������ί��(� :��^�L�n�p����� ��ܿ�п� �6�$� Z�H�jϐ�rϴϢ��� �������2�D�&�h� Vߌ�z߰ߞ������� ����
�@�.�d�R��ZjV 1�w �P����x 
?� ����
�TYPEVFZ�N_CFG ��5d�4�?GRP 1�A�c/ ,B� A� �D;� B����  B4R�B21HELL":�(
��?���<%RS'!�� H3lW�{� �����2XVh������%w����#!0�1�����7��2�0d����HKw 1��� � k/f/x/�/�/�/�/�/ �/�/??C?>?P?b?��?�?�?�?��OMM� ����?��FT?OV_ENB ����+�HOW_REG�_UIO��IMW�AITB�JKO�UT;F��LITI�M;E���OVA�L[OMC_UNIT�C�F+�MON_ALIAS ?e�9? ( he��_ &_8_J_\_B_�_�_ �_�_j_�_�_oo+o �_Ooaoso�o�oBo�o �o�o�o�o'9K ]n����t ���#�5��Y�k� }�����L�ŏ׏��� ���1�C�U�g���� ������ӟ~���	�� -�?��c�u������� V�ϯ������;� M�_�q��������˿ ݿ����%�7�I��� m�ϑϣϵ�`����� ��ߺ�3�E�W�i�{� &ߟ߱������ߒ�� �/�A�S���w��� ��X���������� =�O�a�s���0����� ��������'9K ]����b� ��#�GYk }�:����� �/1/C/U/ /f/�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_O
O�O�O�O�O�O�vO�O__%_7_�C��$SMON_DE�FPRO ����`Q� *SYST�EM*  d=�OURECALL �?}`Y ( ��}9copy f�rs:order�fil.dat �virt:\tm�pback\=>�192.168.�4�P46:224a4>_�_�_l}0�Rmdb:*.*�_��_ �_boto�oc4x�T:\)o�`;oVapUo�o�o
 }5�ea�o�o�g�ohz�
xyzrate 61 +=O����e�w�~5288 ��c�u��� b�_�_:o;�ُ��� o"o��5�яb�t���r�6����emp:�1660 W����:��.��*.d��ƞ`ϟ`�r����1 +� =�O�����)�Ң ��үc�u�������5� ͗ٿ����"���̘ ѿb�tφϙo��K� V����������>� ��h�z�ߟ���:��� ����
�ϸ�A���d� v���.�;������� �ߪ��O�`�r��� �ߩ�2�������� '���K�\n���� 8�������#�� G�j|���3E�W��� ��V472 ��b/t/�/8����*/< �/�/�// �/3)�/a?s?�?3��/-T? �?�?	O�	(�?6&�? fOxO�O�/OAOSO�O0�O_�>�54>��O a_s_�_���/3?4Y�_ �_�_"?�_5X�_bo@to�o���_��8!5=� Wo�o�o�o��o�j�o as��O��<N� ��_(_�s��c� u����_�_5o�gُ� ��o"o���hяb�t�������$SNPX�_ASG 1��������� P 0 '�%R[1]@g1.1����?���%֟��&�	��\� ?�f���u�������� ϯ��"��F�)�;�|� _�������ֿ��˿� ��B�%�f�I�[Ϝ� Ϧ��ϵ�������,� �6�b�E߆�i�{߼� ������������L� /�V��e������ �������6��+�l� O�v������������� ��2V9K� o������ �&R5vYk� ����/��</ /F/r/U/�/y/�/�/ �/�/?�/&?	??\? ??f?�?u?�?�?�?�? �?�?"OOFO)O;O|O _O�O�O�O�O�O�O_ �O_B_%_f_I_[_�_ _�_�_�_�_�_�_,o o6oboEo�oio{o�o �o�o�o�o�oL /V�e���� ����6��+�l��O�v�������PAR�AM ������ �	��P�����OFT�_KB_CFG � ⃱���PIN_SIM  ����C�U�g�����R�VQSTP_DS�B,�򂣟����S�R �/�� &�  AR������TOP_ON_+ERސ����PTN /��@�A	�RI�NG_PRM� ���VDT_GR�P 1�ˉ�  	������������ Я�����*�Q�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߣ� �߲����������� 0�B�i�f�x���� ���������/�,�>� P�b�t����������� ����(:L^ p�������  $6HZ�~ �������/  /G/D/V/h/z/�/�/ �/�/�/�/?
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8___\_���VPRG_COUNT��@���R'ENBU��UM�S���__UPD 1�>/�8  
s_� oo*oSoNo`oro�o �o�o�o�o�o�o+ &8Jsn��� ������"�K� F�X�j���������ۏ ֏���#��0�B�k� f�x���������ҟ�� ����C�>�P�b��� ������ӯί������UYSDEBU)G�P�P�)�d�YH�SP_PASS�U�B?Z�LOG [��U�S)�9#�0�  ��Q)�?
MC:\��6���_MPC���U�$��Qñ8� �Q趿SAV ���ج�ǲ%�ηSV�;�TEM_TIM�E 1��[ (��P'�T&y�ؿT1?SVGUNS�P�U�'�U���ASK_OPTION�P��U�Q�Q��BCC�FG ��[u� 1n�X�G�`a�gZ o��߃ߕ��߹����� ��:�%�^�p�[�� ������� ����� 6�!�Z�E�~�i���������%�������& 8��nY�}� ?��ԫ ��( L:p^��� ����/ /6/$/ F/l/Z/�/~/�/�/�/ �/�/�/�/2?8 F? X?v?�?�??�?�?�? �?�?O*O<O
O`ONO �OrO�O�O�O�O�O_ �O&__J_8_n_\_~_ �_�_�_�_�_�_o�_  o"o4ojoXo�oD?�o �o�o�o�oxo. TBx��j�� ������,�b� P���t�����Ώ��ޏ ��(��L�:�p�^� ������ʟ��o� �6�H�Z�؟~�l��� ����د���ʯ �� D�2�h�V�x�z���¿ ���Կ
���.��>� d�Rψ�vϬϚ��Ͼ� ������*��N��f� xߖߨߺ�8������� ��8�J�\�*��n� ������������"� �F�4�j�X���|��� ����������0 @BT�x�d�� ���>,N tb������ /�(//8/:/L/�/ p/�/�/�/�/�/�/�/ $??H?6?l?Z?�?~? �?�?�?�?�?O�&O 8OVOhOzO�?�O�O�O �O�O�O
__�O@_._ d_R_�_v_�_�_�_�_ �_o�_*ooNo<o^o �oro�o�o�o�o�o�o  J8n$O� ����X����4�"�X�B�v��$T�BCSG_GRP� 2�B���  �v� 
? ?�  ���� ��׏�������1���U�g�z���ƈ�d�, ���?v�	� HC��d�>󙚲�e�CL  �B���Пܘ��ݸ��\)��Y g A�ܟ$�B�g�FB�Bl�i�X�ɼ�|��X��  D	J���r�����C����$үܬ���D�@v�=� W�j�}�H�Z���ſ���������v�	V3.00���	m61c�	�*X�P�u�g�p�>ə��v�(:�� ���p͟�  O�����p�����z�JC�FG �B���� ������8���=��=�c� q�K�qߗ߂߻ߦ��� �����'��$�]�H� ��l���������� ��#��G�2�k�V��� z����������� ���p*<N���l �������# 5GY}h�� ��v�b��>�//  /V/D/z/h/�/�/�/ �/�/�/�/?
?@?.? d?R?t?v?�?�?�?�? �?O�?*OO:O`ONO �OrO�O�O��O�O�O _&__J_8_n_\_�_ �_�_�_�_�_�_�_�_ oFo4ojo|o�o�oZo �o�o�o�o�o�oB 0fT�x��� ����,��P�>� `�b�t�����Ώ��� ����&�L��Od�v� ��2�����ȟʟܟ�  �6�$�Z�l�~���N� ����دƯ�� �2� �B�h�V���z����� Կ¿����.��R� @�v�dϚψϪ��Ͼ� ������<�*�L�N� `ߖ߄ߺߨ����ߚ� ������\�J��n� ����������"� ��2�X�F�|�j����� ����������. TBxf���� ���>,b P�t����� /�(//8/:/L/�/ �ߚ/�/�/h/�/�/�/ $??H?6?l?Z?�?�? �?�?�?�?�?O�?O DOVOhO"O4O�O�O�O �O�O�O
_�O_@_._ d_R_�_v_�_�_�_�_ �_o�_*ooNo<oro `o�o�o�o�o�o�o�o &�/>P�/� �������� 4�F�X��(���|��� ��֏����Ə0�� @�B�T���x�����ҟ ������,��P�>� t�b������������ ���:�(�^�L�n� ������2d����� ̿�$�Z�H�~�lϢ� ���������Ϻ� �� 0�2�D�zߌߞ߰�j� ���������
�,�.� @�v�d������� ������<�*�`�N� ��r����������� ��&J\�t� �B������ F4j|��^�����/�  92 6# 6&J/�6"�$TBJOP_GRP 2����  �?�X,i#�p,�� �x�J� �6$�  �< �� =�6$ @2 �"	 �C�� �&b  Cق'�!�!�>���
559>��0+1�33=�CL� fff}?+0?�ffB� �J1�%Y?d7�.��/>w��2\)?�0�5���;���hCY� �  @�� �!B�  A��P?�?�3EC�  �D�!�,�0*BO�ߦ?�3JB��
:_���Bl�0��0��$�1�?O6!Aəg�AДC�1D�G�6�=q�E6O0��p��B�Q�;��A�� ٙ�@L3D	�@�@_x_�O�O>B�\JU��OHH�1ts�A@�33@?1� C��� �@�_�_&_8_>�#�D�UV_0�LP�Q�30<{�zR� @ �0�V�P!o3o�_<oRi foPo^o�o�o�oRo�o �o�o�oM(�ol@�p~��p4�6&��q5	V3.�00�#m61c�$*(��$1!6�A�� Eo�E���E��E��F��F�!�F8��F�T�Fqe\F��NaF���F��^lF���F��:
F�)F���3G�G���G��G�,IR�CH`��C�dTDU�?�D��D��D�E(!/E\��E��E�h��E�ME��s�F`F+'\�FD��F`=�F}'�F���F�[
F����F��M;S@;Q���|8�`rz(@/&�8�6&<��1��w�^$ESTPARS  *({ _#�HR��ABLE K1�p+Z�6#|��Q� � 1�|�|�P|�5'=!|�	|�
|�Q|�˕6!|�|�u|���RDI��z!ʟܟ� ��$���O������¯ԯ�$����S��x# V��� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����U-����ĜP� 9�K�]�o��-�?�Q��c�u���6�NUM [ �z!� �>  Ȑ����_CFG �����!�@b IMEBF_�TT����x#��a�V�ER��b�w�a�R� 1�p+
 ($3�6"1 ��  6! ���������� �9�$� :�H�Z�l�~����������������^$��_���@x�
b MI__CHANm� x�} kDBGLV;0�o�x�a!n ETHERAD ?�� �y�$"��\&n ROUT���!p*!*�SNMASK�x#�255.h�f�x^$OOLOFS�_DI��[ՠ	O�RQCTRL �p+;/���/+/ =/O/a/s/�/�/�/�/��/��/�/�/!?��PE_DETAI���PON_SVO�FF�33P_MOON �H�v�2-9�STRTCHK ����42VT?COMPATa8��24:0FPROG {%�%CA)�&O�3ISPLAY���L:_INST_�MP GL7YDUqS���?�2LCK�L�PKQUICKMExt �O�2SCRE�@��
tps���2�A�@�I��@_�Y���9�	SR_G�RP 1�� ���\�l_zZ�g_�_�_�_�_�_�^� ^�oj�Q'ODo/oho Se��oo�o�o�o�o �o�o!WE{�i������	�1234567���!���X�E1��V[
 �}ip�nl/a�gen.htmno���������ȏ~�Panel setup̌}�?��0�B�T�f� ��񏞟��ԟ ���o����@�R�d� v������#�Я��� ��*���ϯůr��� ������̿C��g�� &�8�J�\�n������ ����������uϣϙ� F�X�j�|ߎߠ���� ;�������0�B�߾*NUALRMb@G7 ?�� [�� ����������� �� %�C�I�z�m�������~v�SEV  �����t�ECFG� Ձ=]/BaA�$   B�/D
 ��/C�Wi{ �������h PRց; �(To\o�I�6?K0(%����0��� ��//;/&/L/q/�\/�/�/�/l�D ؅Q�/I_�@HI�ST 1ׁ9  �(  ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1?v?�?�?�?�� >?P=71c?�?	O�O-O�?�:edit[2CAR�?|O�O�Op�OAO�?]0962kO� __$_6_�O�O�A36�O�_�_�_�_IR�_ �_�_oo+o=o�_ao so�o�o�o�oJo�o�o '9I|��a81 �ou������o ���)�;�M��q� ��������ˏZ�l�� �%�7�I�[����� ����ǟٟh����!� 3�E�W���������� ïկ�v���/�A� S�e�Pb������ѿ ������+�=�O�a� s�ϗϩϻ������� ߒ�'�9�K�]�o߁� ߥ߷��������ߎ� #�5�G�Y�k�}��� �������������1� C�U�g�y���v����� ������	�?Q cu��(��� �)�M_q ���6���/ /%/�I/[/m//�/ �/�/D/�/�/�/?!? 3?�/W?i?{?�?�?�? �����?�?OO/OAO D?eOwO�O�O�O�ONO `O�O__+_=_O_�O s_�_�_�_�_�_\_�_ oo'o9oKo�_�_�o �o�o�o�o�ojo�o #5GY�o}������?��$U�I_PANEDA�TA 1������  	�}�0�B�T�f�x��� )����mt �ۏ����#�5��� Y�@�}���v�����ן �������1��U�g��N������ �1 ��Ïȯگ����"� u�F���X�|������� Ŀֿ=������0� T�;�x�_ϜϮϕ���@�������,ߟ�M� �j�o߁ߓߥ߷��� ���`��#�5�G�Y� k��ߏ�������� ������C�*�g�y� `���������F�X�	 -?Qc����� �����~ ;"_F��|� ����/�7/I/ 0/m/�����/�/�/�/ �/�/P/!?3?�W?i? {?�?�?�??�?�?�? O�?/OOSOeOLO�O pO�O�O�O�O�O_z/ �/J?O_a_s_�_�_�_ �O�_@?�_oo'o9o Ko�_oo�oho�o�o�o �o�o�o�o#
GY @}d��&_8_� ���1�C��g��_ ��������ӏ���^� ��?�&�c�u�\��� ����ϟ���ڟ�)� �M����������� ˯ݯ0�����7�I� [�m����������ٿ �ҿ���3�E�,�i� Pύϟφ��Ϫ���Z�l�}���1�C�U�g�yߋ�)߰�#����� �� ��$�6��Z�A� ~�e�w�������� ���2��V�h�O������v�p��$UI_�PANELINK� 1�v��  �  ���}1234567890����	 -?G ���o� ����a�� #5G�	����p&���  R�� ���Z��$/6/ H/Z/l/~//�/�/�/ �/�/�/�/
?2?D?V? h?z??$?�?�?�?�? �?
O�?.O@OROdOvO �O O�O�O�O�O�O_ �O�O<_N_`_r_�_�_�0,���_�X�_�_ �_ o2ooVohoKo�o oo�o�o�o�o�o�o ��,>r}���� �������� /�A�S�e�w������ ��я���tv�z�� ��=�O�a�s����� ��0S��ӟ���	�� -���Q�c�u������� :�ϯ����)��� M�_�q���������H� ݿ���%�7�ƿ[� m�ϑϣϵ�D����� ���!�3�Eߴ_i�{� 
�߂����߸���� ��/��S�e�H��� ~��R~'�'�a�� :�L�^�p��������� ������ ��6H Zl~���#�5� �� 2D��h z�����c� 
//./@/R/�v/�/ �/�/�/�/_/�/?? *?<?N?`?�/�?�?�? �?�?�?m?OO&O8O JO\O�?�O�O�O�O�O �O�O[�_��4_F_)_ j_|___�_�_�_�_�_ �_o�_0ooTofo�� �o��o��o�o�o ,>1bt�� ��K����(� :����{O������ ʏ܏�uO�$�6�H� Z�l���������Ɵ؟ ����� �2�D�V�h� z�	�����¯ԯ��� ���.�@�R�d�v��� �����п���ϕ� *�<�N�`�rτ��O�� ��Io���������8� J�-�n߀�cߤ߇��� �߽����o1�oX� �o|��������� ����0�B�T�f��� ������������S�e� w�,>Pbt�� '����� :L^p��#� ��� //$/�H/ Z/l/~/�/�/1/�/�/ �/�/? ?�/D?V?h? z?�?�?�???�?�?�? 
OO.O��ROdO�߈O kO�O�O�O�O�O�O_ �O<_N_1_r_�_g_�_�7OM�m�$U�I_QUICKM�EN  ���_AobRE�STORE 1��  �|��Rto�o�im�o�o�o�o�o :L^p�%�� ����o���� Z�l�~�����E�Ə؏ ���� �ÏD�V�h� z���7�������/��� 
��.�@��d�v��� ����O�Я����� ßͯ7�I���m����� ��̿޿����&�8� J��nπϒϤ϶�a� ������Y�"�4�F�X� j�ߎߠ߲������߀����0�B�T�gS�CRE`?#m�u1sco`�u2��3��4��5*��6��7��8��b�USERq�v��TLp���ks����4��U5��6��7��8���`NDO_CFG� �#k  n` �`PDATE ����No�nebSEUFR�AME  �T�A�n�RTOL_A�BRTy�l��EN�B����GRP 1��ci/aCz  A�����Q�� $6HRd��`�U�����MSK � �����Nv��%�U�%���bV�ISCAND_M;AX�I���FAIL_IMG�� �PݗP#��IMREGNUM�9
,[SIZ�n`��A�,VONOTMOU��@����2��a���a�����FR:\ � MC:\��\LOG�B@F� !�'/!+/O/��Uz MCyV�8#UD1r&�EX{+�S�PPOO64_��0'f�n6PO��L!Ib�*�#V���,�f@�'�/� =�	�(SZV�.�����'WAI�/S?TAT ����P!@/�?�?�:$�?�?���2DWP  ?��P G@+b=��� H�O�_JMPERR �1�#k
  �2�345678901dF�ψO{O�O�O�O �O�O_�O*__N_A_�S_�_
� MLOWpc>
 �_TI��=�'MPHA�SE  ��F�|�PSHIFT�k1 9�]@<�\ �Do�U#oIo�oYoko �o�o�o�o�o�o�o6 lCU�y� ���� ��	�V��-�e2����	V�SFT1�2	V:M�� �5�1G�� ���%A�  �B8̀̀�@ p�كӁ˂�у��z�ME@�?�{��!c>W&%�aM1��k��0�{ �$`0TDINEND��\�AO� �z����S���w��P���ϜRELE�Q��Y���~\�_ACTIV�x�:�R�A ��0e���e�:�RD� ����YBOX �X9�د�6��02����190.�0.�83�N�254��QF�	 �X�j��1��robot����   �p�૿�5pc ��̿�����7������-�f�ZABC�����,]@U��2ʿ�e� �ωϛϭϿ����� � ��V�=�z�a�s߰�E�Z��1�Ѧ