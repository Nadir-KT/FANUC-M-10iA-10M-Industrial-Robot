��   �A��*SYST�EM*��V7.5�0130 3/�19/2015 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP � ��$8 A~O  ���z�����o VIR�TUALw�'D�EF\ � � �����ENOABLE� ������LIST 1� ��  @�!������ 
[.@�d�� ���/�3//W/ */</�/`/�/�/�/�/ �/�/�/??S?&?8? J?�?n?�?�?�?�?�? O�?�?OO"OsOFO�O jO|O�O�O�O�O_�O �O7__\_B_�_f_x_ �_�_�_�W