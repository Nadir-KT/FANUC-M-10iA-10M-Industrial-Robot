��  �}�A��*SYST�EM*��V7.5�0122 8/�1/2   A�K  ����A�BSPOS_GR�P_T   � $PARAM�  ����ALRM_REC�OV1   �$ALMOENB���]ONi�A�PCOUPLED�1 $[PP_�PROCES0 � �1�!~H PCUREQ1� � $SO{FT; T_ID��TOTAL_EQf� $� � NO��PS_SPI_I�NDE��$�X��SCREEN_�NAME ^�SIGN���� PK_FIL~	$THKYM�PANE�  	$DUMMY )� u3|4|G�RG_STR1� � $TIT�P$I��1��{�����5��6�7�8�9�0��z���T��1�1�1 '�1
'2"��ASBN_CFG1 � 8 $CNV_JNT_* �|$DATA_�CMNT�!$F�LAGS�*CH�ECK�!�AT_�CELLSETU�P  P �$HOME_IO�,G�%�#MAC{RO�"REPR�(^-DRUN� D|�3SM5H UT�OBACKU0� � $ENAyB��!EVIC��TI � D6� DX!2ST� ?0�B�#$INTER�VAL!2DISP�_UNIT!20_�DOn6ERR�9FgR_F!2IN,�GRES�!0Qy_;3!4C_WA�4H71�8GW+0�$Y �$DB� 6CO5MW!2MO� H�.	 \rVE��1$F�RA{�$O�UDcB]CTM�P1_FtE2}G1�_�3�B�2I'��AXD�#
 �d $CARD�_EXIST4�$FSSB_TY�P!AHKBD_YSNB�1AGN Gn� $SLOT�_NUM�APR{EV4DEBU� �g1G ;1_EDIT�1 � 1G�=� S�0%$�EP�$OP��U0LETE�_OK�BUS�P7_CR�A$;4AV�� 0LACIw�1�R�@k �1$@ME=N�@$D�V�Q@`PvVA{QL� ;OU&R ,A�0��!� B� LM_�O�
eR�"CAM9_;1 xr?$ATTR4�@�� ANNN@5IMG_HEIGH�A�XcWIDTH4V�T� �UU0F_A�SPEC�A$M��0EXP�.@AX�f�CF�D X� $GR� � S��!.@B�PNFLIx�`�d� UIRE 3<T!GITCH+C�`5N� S�d_LZ`AC��"�`EDp�dL
� J�4S�0� <za�4 q;G0 �� 
$WARNM��0f�!�@� -s�pN{ST� CORN�"�a1FLTR{uTR�AT� T}p  $ACCa1�p�8�|{�rORI�P�C6�kRT0_S~B\q�HG,I1 �[ T�`�"3I�pT�YD�@*2 3``#@� �!�B*HDDcQJ* Cd�2_�3_�U4_�5_�6_�7_�U8_�94"\qO�$ <� �o�o�hK3� 1#`O_Mc@AC/ t � E#63NGPvABA� �c�1�Q8��`,��@nr1�� d�P�0e���axnpUP&Pb2�6���p�"J�p_R�rPBC��J�rĘߜJV�@U� B��s}�g�1�"YtP_*0OF�S&R @� RO1_K8T��aIT�3T�ONOM_�0�1p�p34 >��D �� �Ќ@��hPV��mEX�p� �0g0ۤ�p�r�
$TF�2C$M�D3i�TO�3�0U�� F� ��H�w2tC1(�Ez�g0�#E{"F�"F�40C�P@�a2 �@$��PPU�3N1)ύRևAX�!D�U��AI�3BU�F�FODt�1 �|pp���pPITV� PP�M�M��y��F�SIMQ�SI�"ܢVAڤT�3�=�w T�`(zM��P�B�qFACTb�@EW�P1��BTv?�MC�5 �$*1JB`p脎*1DEC��F���%�=�� �H0CHNS_EMP1�G$G��8��@_4��3�p|@P��3�TC c�(r/�0-sx��ܐ�� MBi��!����JR|� i�SEGFR���Iv �aR�TpN�C��PVF4>�bx &��f{u Jc!�Ja��� !28�ץ8�AJ���SIZ�3S�c�B�TM���g��JaRSINFȑb��Ӏq�۽�н����Lp�3�B���CRC�e�3CCp����c� �mcҞb�1J�cѿ�.�T���D$ICb�Cq��5r�ե��@v�'���E�V���zF��_��FR,pN��ܫ�?�84�0A�! �r�� �h�Ϩ��p�2�͕a��� �د]pR>�Dx ϏᏐ�o"27�!ARV�O`CN�$LG�pV�B�1 �P��@�t�aA�0'��|�+0Ro�� ME`p`"1 CRA 3� AZV�g6p�OF �FCCb�`�`F�`pK������ADI� �a�A�bA'�.p��p�`�c�`S4PƑ�a&�AMP��-`Y�3P�IM�]pUR��QUA1w  $@TITO1�/S@S�!����"0�?DBPXWO��B0=!5�$SK���2&�DBq�!"�"�;PR�� 
� =�����!# S q1M$2�$z���L�)!$�/���� %�/�$�C�!&?�$ENE��q.'*?�Ú R�E�p2(H z��O�0#$L|3$$�#�B[�;���F�O_D��RO�Sr�#������3R�IGGER�6PA�pS����ETURN��2�cMR_8�TUrw��0EWM�ҍM�GN�P���BL�AH�<E���P��'&$P� �'P@�Q"3�CkD{��DQ���4�11��FGO_A7WAY�BMO�ѱQ�#!� CS_�)7  �PIS� I  gb {s�C��A��[ �B$�S��AbP�@r�EW-�TNTVճ�BV�Q[C�(c`�UW�r�P�J��P�$0��S�AFE���V_SV>�bEXCLU�砝nONL2��SY��*a&�OT�a'�HI_V�'��!�A���_ *P0� 9�y_z��p #\pv�ASG�� +nr r�@6Acc*b��G�#@�E�V.iHb?fANNcUN$0.$fdID�	U�2�SC@�`�i�a���j�fa�pOGuI$2,O�$Fib�W$}�OT9@�1 $DUMMYk��da��dn�� � �E�- ` ͑HE�4(sg�*b�SAB��SoUFFIW��@�CA=�c5�g6�raMSW�E. =8Q�KEYI5��ӃTM�10s�qA�vI�N����a��/ �D��HOST_P!�rk��ta��tn��tsp�pEMӰV��� �SBLc ULI�0  8	=ȳ#����DTk0�!1� � $S��ESAMPL��j�۰f爒�f���I�0��[ $SUB�k�#0�Cp��T�r#a�SAVʅ ��c���C��P�f�P$n0E�w YN�_B#2 0Q�D�I{dlpO(��9#�$�R_I�� �ENC2_S� 3  5�C߰�f�- �SpU����!!4�"g�޲�1T���5X�j`ȷg��0��0K�4�AaŔAV�ER�qĕ9g�DSP�v��PC��r"�(���ƓVALU�ߗHE�ԕM+�I�Pճ��OPP ���TH��֤��P�SH� �۰F��df��J� ���C1+�6 H�bLL_DUs�~a3@{��3:���OTX"���s�"~�0NOAUTO�!7�p$)�$�*��c�4�(�Cy�8�C�, �"a&�L�� �8H *8�L H <6����c"�`,  `Ĭ�kª�q��q��Psq��~q��7��8���9��0����1��1�̺1ٺ1�1�1� �1�1�2(�2T����2̺2ٺ2�U2�2 �2�2ʕ3(�3��3��̺3�ٺ3�3�3 �3
�3�4(�ɢT�?��!9 <�9�&�z���I��1���M��QFqE@'@� : ,6���Q? �@P?Q9��5�9�E�@�A�a�A� ;p�$TP�$VA�RI:�Z���UP2f�P< ���TDe� ��K`Q����q��wBAC�"= T�p��e$)_,�bn�kp+ IFIG�kp�H  j��P��p�F@|`�!>t ;E�4�sC�ST�D� D���c�<� 	 C��{��_���l����R  ���FORC�EUP?b��FLUS�`H�N>�F ��^�RD_CM�@E������� ��@vMP��REMr F�Q��1��P���7Q
K4	NJ��5EFFۓ:�@I�N2Q��OVO�O{VA�	TROV���DTՀ�DTMX� ��@�
ے_P`H"p��CL��A_TpE�@�pK	_(�FY_T��v(��@%A;QD� �����`�!0tܑ�0RQ��"�_�a����M�7�sCL�dρRIV'��{��EARۑIOFHPC�@����B�Bƅ�CM9@���R ��GCLF�e!DaYk(M�ap#5Tu�DG��� �%6'��FSSD �s?C P�a�!�1���PQ_�!�(�!1��E�3�!3�+5�&�GR)A��7�@��;�P�W��ONn��EBUG_SD2H`{�_E A �p|뀦`�TERM`5yBi5�p�ORI#�e0Ci5$Z �S#M_�P��e0D�6`�TA�9Ei5{���UP\�F� -�A{�AdPw3S@�B$SEG�:� E�L{UUSE�@NFIJ�B$�;1�p�4��4C$UFlP=�C$,�|QR@���_G90Tk�D�~SNST�PAT����AOPTHJ3Q�E�p %B`�'EC����AR$P�I�aSHF�Ty�A�A�H_SH�ORР꣦6 �0$��7PE��E�OVRH=��aPI�@�U�b= �QAYLOW���IE"�r�A��?���ERV��XQ�Y�� mG>@�BN��U����R2!P.uASYMH�.uAWJ0G�ѡAEq�A�Y�R�Ud@>@��EC���EP;�XuP;�6WOR>@M`�0SMT6�G�3�GR��13�aPA�L@���`�q�uH �� ���TOC�A�`P	P�`$O�P����p�ѡ�`�0O��RE�`R�4C�AO�p낎Be��`R�Eu�h�A��eo$PWR�IMu��RR_�c�q�b=B �I&2H���p_A�DDR��H_LE�NG�B�q�q�q$�Rj��S�JڢSS��SKN��u���u̳�u�ٳSE�A� D��HS��MN�!K�����b����OLX��p����`ACRO3pJ�@���X�+��Q��6�OU)P3�b_�IX��a�a1��}򚃳���( ��H��D��ٰ��氬��IO2S�D�������`�7�L� $d��`Y!_OFyFr�PRM_���#�HTTP_�+�H:�M (|pOcBJ]"/���$���LE~Cd���N � ��֑AB_�TqᶔS�`H�LVh�KR"uH�ITCOU��BG�LO�q���h�`����`��`SS� ����HW��#A:�O�ڠ<`INCPU>2VISIOW�͑���n��to��to�ٲ ��IOLN��P �8��R��p$S�Lob PUT_&n�$p��P& ¢���Y F_AS�"Q��$L������Q"  U�0	P4A��^���ZPHY��-������UOI �#R ` �K����$�u�"pPpk���$���Z����UJ5�S-�v��NE6WJOGKGN̲DIS����Kp�L��#T (�uAVF��+`�CTR�C
�FgLAG2��LG�d�U ���؜�13LG_SIZ����bŰ4�a��a�FDl�I `�w� m�_�{0a�^� �cg���4�����Ǝ����{0��� SCH_<���a�LN�d�VW���E�"����D4��UM�Aљ`LJ�n@�DAUf�EAU��p��d|�r�GH�b�6�OGBOO��W�L ?�6 ITp��y0�REC��GSCR ܓ�D
�<\���MARGm�!���զ ��d%�����S�����W���U� �J{GM[�MNCHJ���FNKEY\�Kn��PRG��UF���7P��FWD��HL.��STP��V��=@X��А�RS��HO`����C9T��b ��7�[�UL���6�(RD�� ����Gt��@POЛ�������MD�FO{CU��RGEX���TUI��I��4� @�L�����P@����`��P��NE���CANA��Bj�V7AILI�CL !�U?DCS_HII4�D�s�O�(!�S����S����_�BUFF�!X�?PTH$m���vP`�ěԃ�AtrY��?P��j�3��`OS1Z2Z3Z����|� � Z � ���[aEȤ��ȤIDX�dPSRrO���zAV�STL�R}�Y&�~� Y$E�C���K�&&����![ LQ��+00� 	P���`#qdt
�U�dw�<���_ \ �?�4Г�\��Ѩ#\0C�4�] ��CLD�PL��UTRQLI��dڰ�)�$FLG &�� 1�#�D���'�q0LD�%�$�%ORGڰ5�2�PVŇVY8��s�T�r�$}d^ ����$6��$�%S�`T�� �B0�4�6RCLMC�4]?o?�9�渰MI�p}d_ d�=њRQ��DgSTB�p� ;Fl�HHAX�R JH>dLEXCESrD�RBM!p�a`ip/BP�T�F��`a�p=F�_A7Ji��KbOtHw�MK�db \Q����v$MBC�LI�|�)SREQUIR�R�a.\o�AXDEB�UZ�ALt M��c@�b�{P����2A#NDRѧ`�`d;�2��ȺSDC��N�IN@l�K�x`��X� N&���aZ���UPST�� ezrLOCf�RIrp�EX<f�A�p�9AAODA�Q��f XY�OND�rMF,Łf�@s"��}%�e/� �b��FX3@IGG�� g ��t"��ܓhs#N�s$R�a%���iL��hL�v�@�D'ATA#?pE�%��tR��Y�Nh t_ $MD`qI}�A)nv� ytq�ytHP`��Pxu��(�zsANSAW)�yt@��yuD+��)\b���0o�i �@CUw�V�p 0XewRR2��j Du��{Q��7Bd$CALIIA@��G��2���RIN��"�<E�NTE��Ck�r^�آXXb]���_N�qlk�@��9��b����Bm��7DIVFDH�@��:�qnI$V,��Sv�$��$Z��X�o�*����o�H �$BEL�T�u!ACCEL��.�~�=�IRC��� ���D�T�8��$PS�@�"L�@ �r��#^�S�Eы T�PATH3���I���3x�p�A_W��ڐ����2nC��4�_M=G�$DD��T���$FW�Rp9���I�4��DE7�P�PABN��ROTSPEE�[g�� �J��[�C@4��@�$USE_+�VP�i��SYY���1 ��aYN!@A�ǦOsFF�qǡMOU��3NG���OL����INC�tMa6��HBx��0HBENCS+��8q9Bp�4�FDm�IN��IԒ]��B��V�E��#�y�23_UyP񕋳LOWL�A��p� B���Du�@9B#P`�x ���BCv��r�MOSI��BM�OU��@�7PERC7H  ȳOV��â 
ǝ����D�Sc@F�@MP����� Vݡ�@y�j�LUk��GjĆp�UP=ó���ĶT�RK��AYLOA�Qe��A��Ԓ����8N`�F�RTI�A$��MOUІ�HB�BS0�p7D5���ë�Z��DUM2ԓS_�BCKLSH_C Ԓk����ϣ����=���ޡ �	ACLA�L"q��1Л��C�HK� �S�RT�Y��^�%E1Qq_��޴_UM�@�C�#��SCL0�r�LMT_J1_L��"9@H�qU�EO�p��b�_�e�k�e�SPC`��u���N�PC�BN�Hz \P��C�0�~"XT��CN_b:�N9��I�SF!�?�V���U�/���ԒdT���CB!�SH� :��E�E1T�T����0y���T��PA ��_P��_� =��Ơ���!����J6 L��@��OG�G�ToORQU��ONֹ���E�R��H�E�g_	W2���_郅T���I�I�I��	Ff`xJ�1�~1��VC3�0BD:B�1��@SBJRK�F9�0DBL_�SM��2M�P_D9L2GRV��0��fH_��d���COS���LNH���������!*,�aZ���fMY�_(��TH��)THET=0��NK23���"l��CB�&CB�CAA�B�"��!��!Ư&SB� 2�%GT	S�Ar�CIMa������,4#97#$DU���H\1� �:Bk6�2�:AQ(rSf$NE�D�`I��B+5��	$̀�!A�%�5�7���LPH�E�2���2SC%C%�2�-&FC0JM&̀V�8V��8߀LVJV!KV�/KV=KVKKVYKVgIH�8FRM��#X�!KH/KH=KHKKH�YKHgIO�<O�8OT�YNOJO!KO/KUO=KOKKOYKOM&�F�2�!+i%0d�7S�PBALANCE�_o![cLE0H_�%SPc� &�b&�b>&PFULC�h�b��g�b%p�1k%�U�TO_��T1T2�i/�2N��"�{� t#�Ѱ`�0�*�.��T��OÀ<�v IN�SEG"�ͱREV84vͰl�DIF�ŕ��1lzw��1m��OaBpq�я?�MI{����nLCHWAR�Y�_�AB��!�$MECH�!o ��q�AX��P����7Ђ�`n 
�d(�nU�ROB��CRr��H���ʀMSK_|f`�p P �`_��R/�k�z�����1S�~�|�z�{���z���qINUq�MT�COM_C� �q�  ���pO��$NOREn�����pЂr 8p G�Re�uSD�0AB��$XYZ_D�A�1����DEBU�Uq������s z`$COD�� �L���p�$B�UFINDX|��c�=�MORm�t $فUA��֐�Р�r�<��rG��u� � $SIMUL  S�*�Y�̑a��OBJE�`̖AD�JUS�ݐAY_	IS�D�3���_FI�=��T u 7�~�6�'��p} =��C�}p�@b�D��FRiIr��T��RO@ �\�E}��c�OPsWOYq�v0Y��SYSBU/@v�$�SOPġd���ϪU<Ϋ}pPRUN����PA��D���rɡL�_OUo顢q�{$)�IMAG��iw��0P_qIM���L�INv�K�RGOVRDt��X�(�aP*�J�|��0L_�`0]��0�RB1�0e��M��ED}�*�p ��N�PMֲ��o('�w�SL�`�q�w x $OwVSL4vSDI��DEX����#�$��-�V} *�N4�\@#�B�2�G�B�_�M� �q�E� x Hw��p�ЯATUSW���Cp�0o�s���BTM��*��I�k�4��x�\԰q�y Dw�E&���@E�r��7����З�EXE��ἱ������f q�z @�w���UP'��$�pQ�XN������ļ��� �PG΅{� h $SUB�����0_���!�M/PWAIv�P7ãՓLOR�٠F\p˕�$RCVFAILs_C��٠BWD΁|�v�DEFSP!p | Lw����p��\���UNI+������H�R�+�}_L\pP��x�t���p�}H�> �*�j�(�s`:~�N�`KETB�%��J�PE Ѓ~��J0SIZE����X��'���S�OR��FORMAT�`��c X��WrEM�t���%�UX��G��PL�I��p�  }$ˀP_SWI�p�q�J_PL��ALO_ �����A���B��� C��D��$E��.�C_��U�� � �c ���*�J3K0�����TIA4��5:��6��MOM��������ˀB��A�D����������PU� NR����������m��� A$PI�6q��	�� ���K4�)6�U���w`��SPEEDgPG��������� ��4T�� � @��SAMr`��\8�]��MOV_�_$��npt5��5���1���2��������d'�S�Hp�IN� '�@�+����4(x$4+T+GAMMWf|�1'�$GET`��p���Da���

pL�IBR>�II2�$HI=�_g�t��2�&�E;��(A�.� �&LW�-6<�)56�&]���v�p��V��$PDCK���q��_?�����q�&���7��4���9+� ��$IM_SR�pD�s�rF��r�rLE���Om0H]���0�-�pq���PJqUR_SCR�N�FA���S_SA�VE_D��dE@�NOa�CAA�b�d@�$ q�Z�Iǡs	�I� �J �K� ����H�L�� >�"hq������ ɢ�� bW^US�(A�u��M4���a� �)q`��3�WW�I@v��_�q�.MUAo�� ?� $PY+�g$W�P�vNG� {��P:��RA��RH��RO�PL�����q� ��s'�X;�OI�&�Zpxe ���m�� p��ˀ�3s�O�O�O�O��O�aa�_т� | ��q�d@��.v��.v�� d@��[wFv��E���%(s�t;B�w�|�t�P���PMA�QU.a ��Q8��1�٠QTH�HOL�G�QHYS��ES���qUE�pZB��O.τ�  ـPܐ(��A����v�!�t�O`�q��u�"���FA�ÎIROG�����Q2����o�"��p��INFOҁ�׃V�����R�H�OI��� =(�0SLEQ������Y�N����Á���P0Ow0����!E0NU��A�UT�A�COPY��=�/�'��@Mg�N@��=�}1������ ���RG��Á���X_�P�$;ख�`��W��P��@��������EXT_CYC  b�R��RpÁ�r��7_NAe!А����ROv`	�� � ���PORp_�1�E2�SRV ��)_�I�DI��T_ �k�}�'���dЇ������5��6��7��8�i�H�SdB���2��$��F�p��GPL8eAdA
�TAR�Б@ ���P�2�裔d7� ,�0FL`Ѧo@YN��K�M��Ck��PWR+�9ᘐ=��DELA}�d�Y�pAD�aMF�QSKIP4�� �A�$�OB`NeT�} ��P_$� M�ƷF@\bIpݷ�ݷ �ݷd����빸��@Š�Ҡ�ߠ�9���J2R� ��� m4V�EX� TQQ� ����TQ������ ��~`�$�RDC�V�� �`��X)�R��p�����r��m$R�GEAR_� IOBT�2FLG��fipER�DTC���Ԍ�>��2TH2NS}� 1� ��uG T\0 ���u�M\Ѫ`I�d��REF�1Á� yl�h��ENAB��cTPE�04�]�� ���]��ъQn#��*�X�"���� ��2����߼���������3�қ'�9�K�]�o����4�Ҝ�����P�������5�ҝ!�@3�E�W�i�{��6����������������7�ҟ-?Qc(u���8�Ҡ�������SMSKÁ� �p�0���EkA�REM�OTE6����`�@�݂TQ�IO}5��ISTP�PO9W@��� �pJ�"�������E�"�$DSB_SIG!N�1UQ�x�C\�TP~���RS232����R�iDEVIC�EUS�XRSRPA�RIT��4!OPB�IT�QI�OWCONTR+�TQ��?�SRCU� MpSUX/TASK�3N�p�0�p$TATU�PHE#�0�����p_XP�C)�$FREEFROMS	pna��GET�0��UPD2�A�2��SP� :�ߧ� !$USAN�na&�����ERI�0�RpRY$q5*"_j@�Pm1�!N�6WRK9KD����6��QFRIEND�Q�RUFg�҃�0oTOOL�6MY�t�$LENGTHw_VT\�FIR�p�C�@ˀE> +IUF�IN-RM��RGyI�1ÐAITI�b$GXñ3IvFG2v7�G1���p3�B�GP1R�p�1F�O_n 0��!RE��p�53҅�U�TC��3A�A�F ��G(��":��� e1n!��J�8�%���%�]� �%�� 74�OX O0�L��T�3H&��8���%b4J53GE�W�0�WsR�TD����T��M�����Q�T]�$V C2����1�а91�8��02�;2k3�;3 �:ifa�9-i�aQ���NS��ZR$V��2BVBwEV�	V�B;�����&�S�`��F�"�kX�@�2a�PS�E���$r1C��_$Aܠ6wPR��7vMU��cS�t '�/89��# 0G�aV`��p�d�`���50�@��-�
z25S�� ��a�RW����B�&�N��AX�!�A:@LxAh��rTHIC�1�I���X�d1TFE�j��q�uIF_CH��3�qI܇7�Q�pG�1RxV��]��:�nu�_JF~�PRԀ�Ʊ�RVAT��� ��`���0RҦ�sDOfE��COUԱ���AXI���OF�FSE׆TRIG NS���c����h������H�Y��IGM�A0PA�pJ�E�ORG_UNEV��J� �S�����Od �$CА�J��GROU����TO�ށ�!��DSP��JcOGӐ�#��_Pӱ��"O�q����@�&KEP�IR��ܔ�@�M}R��AP�Q^�Eph0��K�SYS��q"K�PG2�BRK �B��߄�pY�=�d����`AD_�����OBSOC���N��DUMMY14�p�@SV�PDE_O�P�#SFSPD_WOVR-���C��LˢΓOR٧3N]0bڦF�ڦ��OV��CSF��p���F+��r!���CC��1q"LC�HDL��RECOQVʤ�0��Wq@M�������RO�#��Ȑ_�+��� @0�e@V�ER�$OFSfe@CV/ �2WD��}��Z2���TR�!���E_FD}O�MB_CM���B��BL�bܒ#��adtVQR�$0p��2�G$�7�AM5��0� eŤ��_M;��"x'����8$CA���'�E�8�8$HBKX(1���IO<�����QPPA�������
��Ŋ����DVC_DBhC;��#"<Ј��r!S�1[ڤ�S�3�[֪�ATIOq �1q� ʡU�3���CABŐ�2�CvP��9P�^�B���_� �SUOBCPU�ƐS�P  �M�)0NS�cM��"r�$HW_C ��U��S@��SA�A�p�l$UNITm�l�_�AT���e�ƐC�YCLq�NECA����FLTR_2_FIO�7(��)&B��LPқ/�.�_SC-T�CF_`�Fb�l���|�FS(!E�e�CHA�1��4�D°"3�RSD��$"}���v�_Tb�PRO��,��� EMi_��a�98!�a !�a��DIR0�RAI�LACI�)RMr�L!O��C���Qq��X#q�դ�PR=�S�AI�pC/�c 	���FUNCq�0rRI�NP�Q�0��2�!RAC �B ��[����[WARn���BL�Aq�A����DAk�\���LD0���Q��qeq�TI"r���K�hPRIA�!r"AF��Pz!=�;��?P,`�RK���MǀI�!�DF_@B�%1n��LM�FAq@HR�DY�4_�P@RS��A�0� �MULS�E@���a ���ưt��m�$�O�$�1$1�o����� x�*�EG� ����!A1R���Ӧ�09�2,%ܲ 7�AXE��RO%B��WpA��_l-��CSY[�W!‎&S�'�WRU�/-1��@�SCTR������Eb� 	�%��J��AB�� ���&9�����OT�o0 	$��ARAY�s#2��Ԓ�	ё�FI@��$LI�NK|�qC1�a_��#���%kqj2XYZ��t;rq�3�C1)j2^8'0B��'��4����+ �3FI����7�q����'��_�Jˑ���O3�QOP�_�$;5���ATB�A�QBC��&�DU�β�&6��TURN ߁"r�E11:�p��9GFL�`_���* �@�5��*7��Ʊ 1�J� KŐM��&8��p�"r��ORQ�� a�(@#p=�j�g��#qXU�����mTOV	EtQ:�M��i���U��U��VW�Z�A�W b��T{�, ��@;�uQ ���P\�i��UuQ�We0�e�SERʑe�	��E� O���UdA as��4S�/7����AX��B�'q�� E1�e��i��irp�j J@�j�@�j�@�jP�j @ �j�!�f��i��i ��i��i��i�y �y�'y�7yTqHyoDEBU8�$3 2���qͲf2G + CAB����رnSVS�7� 
#�d��L� #�L��1W��1W�JAW� �AW��AW�QW�@!Ep@?D2�3LAB�2�9U4�Aӏ��C � o�ERf�5� O� $�@_ A��!�PO��à�x0#�
�_MRAt�_� d � T���ٔERR����;T)Y&���I��V�0�cNz�TOQ�d�PL[ ��d�"�� ?�w�! /� pp`T)0���_V1Vr�aӔ��
��2ٛ2�E����@q�H�E���$W������V!��$��P��o�cI��aΣ	� HELL_CF}G!� 5���B_BASq�SR�3��� a#S�b���1�%��2���3��4��5��6ʯ�7��8���RO0����I0�0NL�\C�AB+�����ACK 4�����,�\@2@�&�n?�_PU�CO. U�OUG�P~ ����m�������TPհ_�KAR��_�RE�*��P���7QU�E���uP����CSTOPI_AL7��l�k0��h��]�l0S#EM�4�(�M4�6��TYN�SO���D�IZ�~�A�����m_�TM�MANRQ��k0E����$K�EYSWITCH����m���HE��B�EAT��E- LQE~�����U��F!������B�O_HOM�=OGREFUPPAR&��y!� [�C��9O��-ECOC���>�0_IOCMWD
ǆa�	�m��� �# Dh1���UX����M�βgPgCFORyC��� j��OM.  � @��5(�U�#P, 1���, 3��45~	�NPX_ASt�w� 0��ADD�о�$SIZ���$VAR���TI�P/�.��A�ҹ�M�ǐ��/�1�+ U"S��U!Cz���FRI	F��J�S���5Ԓ��NF�� �� � mxp`SI��TE�C\���CSGL��TQ2��@&����� ��S'TMT��,�P �&�BWuP��SHOW�4���SV�$��� �Q�A00 �@Ma}���� ��ਅ�&���5��6��7*��8��9��A��O ����Ѕ�Ӂ���0��F ��� G��0G���0 G���@G��PG��U1	1	1	1+	U18	1E	2��2��U2��2��2��2��U2��2��2��2��U2	2	2	2+	U28	2E	3��3��U3��3��3��3��U3��3��3��3��U3	3	3	3+	U38	3E	4�4��U4��4��4��4��U4��4��4��4��U4	4	4	4+	U48	4E	5�5��U5��5��5��5��U5��5��5��5��U5	5	5	5+	U58	5E	6�6��U6��6��6��6��U6��6��6��6��U6	6	6	6+	U68	6E	7�7��U7��7��7��7��U7��7��7��7��U7	7	7	7+	e78	7E��VP���UPDs�  ��`NЦ�
�S�YSLOt�� � L��d���A�a�TA�0d��|�AL1U:ed�~�CUѰjg=F!aID_L�Ñe�HI�jI��$FI�LE_���d��$�2�
�cSA>�� �hO��`E_BLC�K��b$��hD_CPUyM�yA��c�o��db����R ��Đ
PW��!� oqLA��S=�ts�q~tRUN�qst�q�~t���qst�q~t ��T��ACCs���X -$�qLEN;��tH��ph�_��I��ǀLOW_A�XI�F1�q�d2�*�MZ���ă��W�Ipm�ւ�aR�TOR���pg�D�Y���LACEk�ւ�pV�ւ~�_MA2�v�������GTCV��؁��T�� ي�����t�V�����V�Jj�R�MA�i�JH��m�u�b����q�2j�#�U�{�t�K�JK��VK;���H����3��J0����JJv��JJ��AAL��Pڐ��ڐԖ4Օ5���N1���ʋƀW�%LP�_(�g����p�r�� `�`GR�OUw`��B��N�FLIC��f�RE�QUIRE3�EB�U��qB���w�2�����p���q5�p��{ \��APPR��iC}�Y�
ްEN٨�CLO7��S_M���H���u�
�qu�7� ���MC������9�_MG��C�C�o��`M�в�N�BRKL�NOL|�N�[�R��_LINђ�|�=�J����Pܔ������������������6ɵ�̲8k����q���� ��
��q�)��7�PATH 3�L�B�L��H�wࡠm�J�CN�CA��ؒ�ڢB�IN�rUChV�4a��C!�UM��!Y,���aE�p�����ʴ���PAYL�OA��J2L`R'_AN�q�Lpp����$�M�R_F2�LSHR��N�LO�ԡ�Rׯ�`ׯ�ACRL_G�ŒЛ� �r�Hj`߂$HM�^��FLEXܣ�q}J�u� :� ������������1�F1�V�j�@�@R�d�v�������E�� ��ȏڏ����"�4� q���6�M���~��U��g�y�ယT��o�X ��H������藕?� ����ǟِݕ�ԕ�����%�7��JJ�� � V�h�z����`AT�採@�EL��� S��J|��v��JEy�CTR���~�TN��FQ��H�AND_VB-����v`�� $��Fa2M����ebSW���q'��� $$	MF�:�Rg�(x�,4�%��0&A�`�=���aM)F�AW�Z`i�A�w�A��X X�'pi�D*w�D��Pf�G�p�)CSTk��!x��!N��DY�pנM�9$`%� ��H��H�c�׎���0� ��Pѵڵ��0������$���� ���1��R�6<��QASYMvř�	��v��J���cі�_SH>��ǺĤ�ED@����������J��İ%��C�IDِ�_V�I�!X�2PV_�UNIX�FThP�J ��_R�5_Rc�cTz�pT �V��@���İ�߷��U� ����'�eT��Hqpˢ��faEN�3�DI�����O4d�`J��) x g"IJAAȱz� aabp�coc�`a�pdq��a� ��OMM�E��� �b�RqAT(`PT�@� S��a7��;�Ƞ�@�h�a�iT��@<� $DU�MMY9Q�$P�S_��RFC�  S�v �p����Pa� XƠ���SuTE���SBRY��M21_VF�8$_SV_ERF�O��\LsdsCLRJtA���Odb`O�p �� D $GL3OBj�_LO���u��q�cAp�r�@aSYS�qADR``�`�TCH  � �,��ɩb�W_NA����7�AD�S�R���l  ���
*?�&Q�0"?� ;'?�I)?�Y)��X��� h���x������)��Ռ �Ӷ�;��Ív�?��O�O�O�DD�XSCR�E栘p����ST��s}y`���S� /_HA�q�� TơgpTYP �b���G�aG�蕵�Od0IS_�䓀d�UEMd� �����ppS�qaR�SM_�q*eUNE�XCEP)fW�`S_}pM�x���g�z�����ӑCOU��S�Ԕo 1�!�UE&���Ubwr��PROG�M�FL@$C�UgpPO�Q��� U�I_�`H� �s 8�� �_HE�P�S�#��`RY �?�qp�b��dp�5��OUS�� �� @6p�v$B�UTTp�RpR�C�OLUMq�e��S�ERV5�PAN�EH�q� � N�@GEU���Fy�~�)$HELPõ^)BETERv�)� ����A � ���0��0��0ҰIN簪c�@N��IH��1��_� �֪�LN�r� ��qpձ_ò=�$H��TEXl�����FLA@��REL�V��D`��������M��?,�ű�m�����"�USR�VIEW�q� <�6p�`U�`�NFyI@;�FOCU��n;�PRI� m�`��QY�TRIP�q�m�UN<`Md� �#@p�*eWARN|)e6�SRTOL%���g��ᴰONCO;RN��RAU����9T���w�VIN�Le�� $גP�ATH9�גCAC�H��LOG�!�LIMKR����v����HOST�!��b�R��OBOT,�d�IM>� �� ���Zq�Zq;��VCPU_AVA�IL�!�EX	�!AN���q��1r��1�r��1 �ѡ�p��  #`C����@_$TOOL�$���_JMP� �<��e$SS�����SHIF��Nc߃P�`ג�E�ȐR�����OSUR��Wk`RADILѮ��_�a��:�9a��`a�r���LULQ$OUTPUT_BM����IM�AB �@�r�TILSCO��C7����� ��&��3��A��@�q���m�I�2G��n�y@Md�}��yDJ�U��N�WAIET֖�}��{�%! {NE�u�YBO��� �� $�`�t�SB@TPE��NECp�J^�FY�nB_T��R��І�a$�[YĭcB��dM���F� �p��$�pb�OP?�M�AS�_DO�
!QT�pD��ˑ#%�|�p!"DELAY�:`7"JOY�@(�nC E$��3@ �xm��d�pY_[�!"g�"��x[���P? Ea�ZABC%�� G $�"R��
ϐ�$$CLAS������!pE`<� � VIRT]��/� 0ABS����1 �5� ?< �!F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6�HZi{0-�AXL�p��"�63  ��{tIN��qztPR�E�����v�p�uL�ARMRECOV� 9�rwtNG��� .;	 A�   �.�0PP7LIC��?5�p��Han�dlingToo�l o� 
V7.50P/23-��  �Pf���
��_SWt� U�P�!� x�F0Ȭ�t���A0v�� 864�� ��it��y� r�2 7DA�5�� �� �Qf@��o�No�neisͅ˰ ���T���!L_Aex>�_l��V�uT��s9�UT�O�"�Њt�y��HGAPON
0g�1���Uh�D 1581����̟ޟry�����Q 1�� �p�,�蘦��ր�;�@��q_��"�2 �c�.��H���D�HTTHKYX��"�-�?� Q���ɯۯ5����#� A�G�Y�k�}������� ſ׿1�����=�C� U�g�yϋϝϯ����� -���	��9�?�Q�c� u߇ߙ߽߫���)��� ��5�;�M�_�q�� ������%����� 1�7�I�[�m������ ����!����-3 EWi{���� ��)/AS ew����/� �/%/+/=/O/a/s/ �/�/�/�/?�/�/? !?'?9?K?]?o?�?�? �?�?O�?�?�?O#O�]���TO�E�W�DO_CLEAN��|7��CNM  � �__/_A_�S_�DSPDRY�R�O��HIc��M@ �O�_�_�_�_oo+o =oOoaoso�o�o���p�B��v �u���aX�t������9�PLU�GG���G��U�PRUCvPB�@��_ĠorOr_7�SEGF}�K[mwxq�O �O�����?rqLAP�_�~q�[�m� �������Ǐُ�����!�3�x�TOTA�L�f yx�USENU�p�� �H���B���RG_STRI�NG 1u�
��Mn�S5��
ȑ_ITEM1Җ  n5�� �� $�6�H�Z�l�~����� ��Ưد���� �2��D�I/O S�IGNAL̕�Tryout M�odeӕInp���Simulat{edבOut��OVERR�P� = 100֒In cycl���בProg A�bor��ב��S�tatusՓ	H�eartbeat�їMH Fauyl��Aler'� W�E�W�i�{ύϟϱ�8������ �CΛ �A����8�J�\�n߀� �ߤ߶����������"�4�F�X�j�|���WOR{pΛ��(ߎ��� �� ��$�6�H�Z�l� ~���������������8 2PƠ� X ��A{���� ���/AS ew�����SDEV[�o�#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C?�U?g?y?PALT ݠ1��z?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O_�?GRI�`ΛDQ�?_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�o2_l�R��a \_�o"4FXj |����������0�B�T��oPREG�>�� f���Ə ؏���� �2�D�V� h�z�������ԟ����Z��$ARG_���D ?	����;�� � 	$Z�	+[O�]O��Z�p��.�SBN_CON?FIG ;��������CII_SAVE  Z������.�TCEL�LSETUP �;�%HOME�_IOZ�Z�%M�OV_��
�RE�P�lU�(�UTOB�ACKܠ��FRA:\z�� \�z�Ǡ'`��z���ǡi�INUI�0z���n�?MESSAG����ǡC���ODE_D������%�O�4�n�oPAUSX!�;�? ((O>��� �ˈϾϬ�������� ��*�`�N߄�rߨ����g�l TSK  �wͥ�_�q�UPD�T+��d!�A�W_SM_CF��;����'�-�GRP� 2:�?� N�B�ŰA��%�XSCR�D1�1
7� �ĥĢ��������� �*�������r����� ������7���[�& 8J\n��*�t�GROUN�Uϩ_UP_NA�:�s	t��_ED��17�
 �%�-BCKEDT-`�2�'K�`����-t�z�q�,q�z���2t1�����q�k�(/��ED3/��/��.a/�/;/M/ED4�/t/)?�/.?p?�/�/ED5`??�?�<?.�?O�?�?ED6O�?qO�?.MO�O'O9OED7�O`O_��O.�O\_�O�OEDa8L_,�_�^-p�_ oo_�_ED9�_�_]o�_	-9o�oo%oCR_ 9]��oF�o�k� � NO�_DEL��GE?_UNUSE���LAL_OUT �����WD_ABORﰨ~��pITR_RTN�=��|NONSk����˥CAM_PARAM 1;��!�
 8
SO�NY XC-56� 2345678�90 ਡ@����?��( �А\�
���{��:��^�HR5q�̹���ŏR57ڏ�A�ff��KOW�A SC310M�
�x�̆�d @<�
���e�^ ��П\����*�<���`�r�g�CE_R�IA_I�!��=�F��}�z� ]��_LIU�]�V����<��FB��GP 1���Ǯ�M�_�q�0�Cg*  ����C1���9��@��G���CVR�C]��d��l��Es��R�����[ԴUm��v�������_�� C����(������=�HE�`O�NFIǰ�B�G_�PRI 1�{ V���ߖϨϺ�����������CHKPA�US�� 1K� ,!uD�V�@�z�d� �߈ߚ��߾������.��R�<�b���OƯ�������_MkOR�� ����<������ 	 �����*�� N�`�������?Ғ�q?;�;����K���9�P���ça�-:���	�

��M���pU�ðț�<��,~��DB��튒)
mc�:cpmidbg��f�:�  %#$¥�p�/��  �I

I� �s>�0�0�)�X��?��p��p�bUg�/� ҋ��Uf�M/w�O/�
?DEF l��s�)�< buf.txts/�t/��ާY�)�	`�����o=L���*MC��1����?43���1��t�īCz�  BHH�CPU�eB�^&B����;��>C����CnY
K�E�?{hDS�D����?r��D���D��^�=�Fǁ,F�M\�F���Cm	fF��F���:X���'w�1����s���.�p���b���BDw�M@x8�̊1( C���( D��p@�0EY�1X��EQ�EJP� F�E�F�� G��>^F� E�� FB�� H,- Ge�߀H3Y��:� � >�33 9���~  n8�~�@��5Y�E>�ðA���Y<#�
"Q ����+_�'RSMOFS�p�.8��)�T1��DE ���F 
Q��;��(P  B_<_��Rb����	op6C4P)�Y
s@ ]AQ�2Js@C�0B3�MaC{@�@*cw��UT�pFPROG %�z�o�oigI�q���v���ldKEY_TBL�  �&S�#� �	�
�� !�"#$%&'()�*+,-./01�i�:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������vq��͓���������������������������������耇���������������������9��p`LCK�l4�<p`�`STAT ��S�_AUTO_DO��5�INDTO_ENB!���R�Q�?�1�T2}�^�STsOPb���TRLr`�LETE��Ċ_�SCREEN ��Zkcsc���U��MMENU� 1 �Y  <�l�oR�Y1�[� ��v�m���̟����� ٟ�8��!�G���W� i��������ïկ�� 4���j�A�S���w� ����迿�ѿ���� T�+�=�cϜ�sυ��� �ϻ�������P�'� 9߆�]�o߼ߓߥ��� �����:��#�p�G� Y����������� $����3�l�C�U��� y����������� ���	VY)�_MAN�UAL��t�DBC�O[�RIGڇ
�DOBNUM� ��B1� e
�PXWOR/K 1!�[�_�U/4FX�_A�WAY�i�GC�P  b=�Pj_A!L� #�j�Y��܅t `�_�  1"�[_ , 
�o�d�&/~&lMZ�I�dPx@P@#ONT�IMه� d��`&�
�e�MOT�NEND�o�RECORD 1(�[qg2�/{�O��! �/ky"?4?F?X?�( `?�?�/�??�?�?�? �?�?)O�?MO�?qO�O �O�OBO�O:O�O^O_ %_7_I_�Om_�O�_ _ �_�_�_�_Z_o~_3o �_Woio{o�o�_�o o �oDo�o/�oS �oL�o����@ ���+�yV,�c� u��������Ϗ>�P� ����;�&���q��� 򏧟��P�ȟ�^�� ����I�[����� � ��$�6�������j�TOLERENC�wB���L���� CS_CFG �)�/'dM�C:\U�L%04�d.CSV�� cl��/#A ��CH��z� //.ɿ��(�S�RC_OUT �*���SG�N +��"���#�09-FEB�-20 18:4�4015-JAN�p�0:51+ P/Vt�ɞ�/.���f�pa�m�?�PJPѲ���VERSION �Y�V2.�0.84,EFLO�GIC 1,� 	:ޠ=�ޠ�L��PROG_E�NB��"p�ULS�k' ����_WRSTJNK ��"f�EMO_OPT_�SL ?	�#
� 	R575 /#=�����0�B��>��TO  �ݵ�l���V_F EX��d�%��PATHw AY�A\�����5+ICT�F�u-�j�#�egS�,�ST?BF_TTS�(�	�d���l#!w�� M�AU��z�^"MSWX�.��4,#�Y�/�
!J�6%�ZI~m��$SB�L_FAUL(�0��9'TDIA[�1�<�� ����12345678#90
��P��H Zl~����� ��/ /2/D/V/h/��� P� ѩ �yƽ/��6�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?�,/�gUMP���� ��ATR���1OC@P�MEl�OOY_TE{MP?�È�3F�8��G�|DUNI��.��YN_BRK �2_�/�EMGDI_STA��]�'�@�NC2_SCR 3�K7(_:_L_ ^_l&_�_�_�_�_)��C�A14_�/oo�/oAoԢ�B�T5�K�ϋo~ol�{_�o �o�o'9K] o������� ��#�5��/V�h�z� �л`~�����ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T���x����� ����ү�����,� >�P�b�t��������� ο����(�f�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� :� �2�D�V�h�z�� �����������
�� .�@�R�d�v������� �������*< N`r����� ��&8J\ n��������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?� �?�?�?�?�?OO,O >OPObOtO�O�O�O�O��O�O�O__NoETMODE 16�5��Q �d��X
X_j_|Q�PRR�OR_PROG �%GZ%�@��_ � �UTABLE  G[�?oo)o�RjRRSEV_N�UM  �`WP��QQY`�Q_A�UTO_ENB � �eOS�T_NONna 7G[�QXb_  *��`��`%��`��`d`+�`�o8�o�o�dHISUc�Q�OP�k_ALM 1]8G[ �A��l�P+�ok}��ȳ��o_Nb�`  �G[�a�R
�:PT�CP_VER �!GZ!�_�$EX�TLOG_REQ�v�i\�SIZ�e�W�TOL  ��QDzr�A W�_BWD�p��xf�́t�_DI�� 9�5�d�T�QsRֆSTEP��:P��OP_DOv��f�PFACTOR_Y_TUNwdM��EATURE �:�5̀rQ�Handling�Tool �� \�sfmEng�lish Dictionary���roduAA� Vis�� Ma�ster����
�EN̐nalog� I/O����g.�fd̐uto S�oftware �Update  �F OR�mat�ic Backu�p��H596�,�ground �Editޒ  1� H5Cam�era�F��OP;LGX�ell𜩐�II) X�omm�Րshw���com揭co���\tp����pane�� � opl��tyl�e select^��al C��nJ�~Ցonitor��gRDE��tr��?Reliab𠧒�6U�Diagno�s(�푥�552�8�u��heck �Safety U�IF��Enhan�ced Rob �Serv%�q )� "S�r�UserG Fr[�����a���xt. DIO 6�fiG� sŢ��wendx�Err�MLF� pȐĳr�r�� ����  !���FCTN Men�u`�v-�ݡ���T�P Inېfac��  ER J�GC�pבk E�xct�g��H55�8��igh-Sp�ex�Ski1�  �2
P��?���m�munic'�on1s��&�l�ur�ې���ST Ǡ��c�onn��2��TX�PL��ncr�s�tru����"FA�TKAREL Cmd. LE�{uaG�545\�ſRun-Ti��E{nv��d
!����ؠ++�s)�S/�W��[�Lic�enseZ��� 4�T�0�ogBook�(Syڐm)��H�54O�MACRO�s,\�/Offs�e��Loa�MH�������r, k�M�echStop �Prot���� l�ic/�MiвSh�if����ɒMixpx��)���xStS��Mode Swiwtch�� R5W��Mo�:�.�� 7#4 ���g��K��2h�ulti-T�=�M���LN (�Pos�Reg�iڑ������d�ݐtO Fun�ǩ�.�����Num~����Ï lne��ᝰ Adjup������  - W��ta�tuw᧒T��RDMz�ot��s�cove U�9����3Ѓ�uesOt 492�*�o������62;�SNP�X b ���8 Jy7`���Libr��FJ�48���ӗ� ����
�6O�� Pa�rts in VCCMt�32���x	�{Ѥ�J990��{/I� 2 P���TMILIB��Ht���P�AccD��L�
TE$TX܍ۨ�ap1S�Te<����pkey���wգ�d��Un�exceptx�motnZ��������3є�� O��΄� 90J�єSP CSXC<�f�l�Ҟ� Py�We}�Β�PRI�>vr\�t�men�� ��/iPɰa������vGrid�play��v��0�)��H1�M-10iA(B201 ��2\� 0\k/�A/scii�l�Т��ɐ/�Col��ԑG7uar� 
�� /�P-�ޠ"K��stN{Pat ��!S��Cyc�҂�or�ie��IF8�ata- quҐ�� ƶ���mH574��RML��am���Pb�HMI De3�(�b����PCϺ�P�asswo+!��"PE? Sp$�[���stp��� ven���Tw�N�p�YEL?LOW BOE	k$wArc��vis���3*�n0WeldW�cial�7�V#Mt�Op����1y�֠ 2F�a�pocrtN�(�p�T1�`T� �� ��xy]ֹ&TX��tw�ig�j�1� b� ct\��JPN ARC?PSU PR��ovݲOL� Sup�2fil� &PAɰא�cro�� "PM�(����O$SS� enвtex�� r����=�t�ssag$T��P��P@�Ȱ�锱�rtW��H'�>r�dpn��n1#
t�!� z ���ascbin4p�syn��+Aj�M� HEL�NCL� VIS PKG�S PLOA`�McB �,�4VW��RIPE GET_VAR FIEo 3\t��FL[��OOL: ADD� R729.FD/ \j8'�CsQ�Q�E��DVvQ�sQNO WTWTE��>}PD  �^��b�iRFOR ��EC�Tn�`��ALSE� ALAfPCPM�O-130  M�" #h�D: H�ANG FROM�mP�AQfr��R7�09 DRAM �AVAILCHE�CKSO!��sQVP�CS SU�@LIMCHK Q +P~d�FF POS��F��Q R593�8-12 CHA�RY�0�PROGR�A W�SAVE�N`AME�P.SV2��7��$En*��p�?FU�{�TRC|� �SHADV0UPD�AT KCJўRS�TATI�`�P M�UCH y�1��I�MQ MOTN-�003��}�ROB�OGUIDE DAUGH�a���*�Gtou����I� Š�hd�ATH�PepM�OVET�ǔVM�XPACK MA�Y ASSERT��D��YCLfqTA��rBE COR �vr*Q3rAN�pR�C OPTION�SJ1vr̐PSH�-171Z@x�tcǠSU1�1Hp^9R!�Q�`_T�P��'��j�d{tby app wa 5IҌ~d�PHI���p�aT�EL�MXSPD' TB5bLu 1��U�B6@�qENJ`CEV2�61��p��s	�may n�0� �R6{�R� �Rtr�aff)�� 40�*�p��fr��sy�svar scr� J7��cj`DJ�U��bH V��Q/��PSET ERR�`J` 68��PN�DANT SCR�EEN UNRE�A��'�J`D�pPA��pR`IO 1����PFI�pB�pG/ROUN�PD��G���R�P�QnRSVIP� !p�a�PDIGI?T VERS�r}B�Lo�UEWϕ P�06  �!��MA�Gp�abZV�DIx�`� SSUE��ܰ�EPLAN {JOT` DEL�p�ݡ#Z�@D͐CAsLLOb�Q ph���R�QIPND��I{MG�R719���MNT/�PES ��pVL�c��Holp�0Cq���tPG:�`:C�M�canΠ���pg.v�S: 3�D mK�view� d�` �p��eat7У�b� of �P�y���ANNOT �ACCESS M���Ɓ*�t4s a��lok��Fle�x/:�Rw!mo?�PA?�-�����`~n�pa SNBPJ AUTO-�0�6f����TB��PIA�BLE1q 636>��PLN: RG$��pl;pNWFMD�B�VI���tWIT� 9x�0@o��Qu�i#0�ҺPN RR�S?pUSB�� t� & removb�@ )�_��&AxEP7FT_=� 7<`�p�P:�OS-14;4 ��h s�g���@OST� � C�RASH DU �9��$P�pW�� .$��LOGI�N��8&�J��6b0�46 issue� 6 Jg��: �Slow �st~��c (Hos`��c���`IL`IMP�RWtSPOT:Wqh:0�T�STYW =./�VMGR�h��T0CAT��hosB��E�q��� �uO�S:+pRTU' �k�-S� ����E:���pv@�2�� t\�hߐ��m ��al�l��0�  $�H� �WA͐��3 CN�T0 T�� Wr}oU�alarm���0s�d � �0SE1����r R{�OMEpBp���K� 55��REàSEst��g�     �KoANJI�no����INISITA�LIZ-p�dn1we�ρ<��dr�� l�x`�SCII L��fails w��� ��`�YSTE�a���o��Pv� IItH���1W�Gro>P�m ol\wpSh�@�P��Ϡn cfslxL@АWRI ЏOF Lq��p?�F��up��de-r�ela�d "A�Po SY�ch�Ab�etwe:0INDc t0$gbDO����r� `�Gig�E�#operab[ilf  PAbHi�xH`��c�lead�\etf�Ps�r��OS 030�&: f{ig��GLA )P� ��i��7Np t�pswx�B��If��g������5aE>�a EXCE#dU��_�tPCLOS��"�rob�NTdpF�aU�c�!���PNIO V750�Q�1��Qa��DB Ė�P M�+P�QED��DET��-� \�rk��ONLINEhSBUGIQ ߔXĠi`Z�IB�S a�pABC JAR�KYFq� ���0MSIL�`� R�pNД� �p0GAR��D�*pR��P�"! jK�0cT�P�Hl#n��a�ZE V�� TwASK�$VP2(��4`
�!�$�P�`WI[BPK05�!FȐ�B/��BUSY oRUNN�� "��ȁ����R-p�LO��N�DIVY�CU9L��fsfoaBW�p���30	�V��ˠIT`�a5�05.�@OF�UGNEX�P1b�af�@��E��SVEMGN� NMLq� D0pCC_SAFEX �0c�08"qD �PE�T�`N@�#J87�����RsP�A'�M��K�`K�H G�UNCHG۔MEKCH�pMc� T� � y, g@�$ ORY LEAKA8�;�ޢSPEm�Ja:��V�tGRIܱ��@�CTLN�T�Rk�FpepR�j506�EN-`IN������p �`�Ǒk!��Tq3/dqo�STO�0)A�#�L�p �0�@�Q�АY�&�;pb1CTO8pP�s���FB�0@Yp`�`DU��a!O�supk�t4 � PЙF� Bnf�Q�PSVGN-1��V�S'RSR)J�UP��a2�Q�#D�q l �O��QBRKCTR5Ұ�|"-�r�<p�c�j!INVP�D ZO� ��T`h#�Q�cHset,|D��"DUAL� w�2*B�RVO117 A�]�TNѫt�+bTa2�473��q.?��sA�Uz�i�B�comp�lete��604�.� -�`haknc�U� F�Нe8��  ��npJ�tPd!q��`��� 5Nh596p�!5d��� "p�P�P�Q�0�P2@�p�A� xP��R(}\*xPe� aʰI����E��1��p� j � � xSt�^t ��A�AxP�q 5 siug��a��"AC;a���
�bCexPb_p��.pc]l<bHbcb_circ~h<n�`tl1�~`xP`o`�dxP�b]o2�� �c�b�c�ixP�jupf�rm�dxP�o�`ex�e�a�oFdxPtpe�d}o��u`�cptlcibxzxP�lcr�xrxP\�blsazEdxP_fm�}gcxP�x@���o|sp�o�mc(�N�ob_jzop�uD6�wf��t��wms�1q��sld�)��jCmc�o\�n��nuhЌ���|st�e��>�p1l�qp�iwck����uvf0uߒ��lv�isn�Cgacu�lwQ
E F  ;! Fc.fd�Qv��� qw���Dat�a Acquis�i��nF�|1�RR6�31`��TR�QDM�CM �2�P75�H�1�P583xP1���71��59`�5�P57<PxP�Q����¨�(���Q��o p�xP!daq\�o�A��@�� ge/�e�tdms�"DMEsR"؟,�pgdD����.�m���-��qacq.<᡾xPmo��Dh���f{�u�`13���MACROs, Sksaff�@z�����03�SR�Q(��Q6���1�Q9ӡ�R�ZSxh��PxPJ643�@�7ؠ6�P�@�PRS��@���e �Q�UС �PIK�Q52 P�TLC�W��xP3 (��p/O��!�P�n �xP5��03�\sfmnmc "MNMCq�<��Qj��\$AcX�FM�� �ci,Ҥ�X����cd�pq+�
�sk�SKx�xP�SH560�,P��,�y�refp "REFp�d�A��jxP	�of�OF�c�<gy�to�TO�_����ٺ����+je�u��caxi�s2�xPE�\�e�q"�ISDTc��]�porax ��MN�x�u�b�isde܃�h�\�w�xP! is_basic��B�� P]��QAxes��R6������.�(sBa�Q�ess� �xP���2�D�@�z�atis���(�{������~��m��F�Mc�u�{�
ѩ�MNIS��ݝ����x�����ٺ��x� j7}5��Devic��� Interfa�c�RȔQJ7540��� xP�Ne`� �xP�ϐ2�б�����dn� "DNE����
tpdnu�i5UI��ݝ	b�d�bP�q_rs�ofOb
dv_aro��u����>�stchkc���z	 �(}onl��G!ffL+H�@J(��"l"/�n�bx��z�hamp���T�C�!i�a"�59`��S�q��0 (�+�P�o�u�!2��xpc�_2pcchm��C�HMP_�|8бpe�vws��2쳌pc�sF��#C SenxPacro�U·�-�R6�Pd�xPk������p��gT�L��1d M�2`��8�1c4ԡ��3 qem��GE�M,\i(��Dgesnd�5���H{�}Ha��@sy���c�Isu�xD��Fmd��I��7��4���u���AccuCal�P�4� ��Rɢ7ޠB0��6+56f�6��99\aFF q�S(�U��2�
X�ap�!Bd��cb_��SaUL��  ��� ?�ܖto��ot�plus\tsr�nغ�qb�Wp��t����1��Tool (N. A.)�[K�7�Z�(P�m�����bfcls� k94�"K4p��qt�pap� "PS�9H�stpswo`��p�L7��t\�q ����D�yt5�4�q��@w�q��� �M�uk��rkey����s���}t�sfeatu�6�EA��� cf)t\�Xq�����d�h5���LRC0�md�!�C587���aR�(�����2V��8c?u3l\�pa3}H�&r-��Xu���t,�� �q "�q�Ot��~,���{@�/��1c�}����y�p �r��5���S�XAg��-�y���Wj874��- iRVis<���Queu�� �Ƒ�-�6�1���(����u���tӑ�����
�tpvtsn? "VTSN�3C�t+�� v\pRDV����*�prdq\�Q<�&�vstk=P�������nm&_�դ��clrqν���get�TX��Bd����aoQϿ�0qstr�D[� ��t�p'Z��Ɵ�npv��@�enlIP0��D!x�'�|����sc ߸��tv�o/��2�q���v b����q���!���h�]��(� Con�trol�PRAuX�P5��556�A�@59�P56.@5�6@5A�J69�$@982 J55?2 IDVR7�hq A���16�H���La��� ��Xe�f�rlparm.fn�FRL�am��C9�@(F������w6{���A��QJ6�43�� 50�0L�SE
_pVAR� $SGSYSC���RS_UNIT�S �P�2�4tA�T�X.$VNUM_OLD 5�1�xP�{�50+�"�` Funct���5tA�� }��`#@�`3�a0��cڂ��9���@HA5נ� �P���(�A ����۶}����ֻ}��bPRb�߶~p{pr4�TPSPI0�3�}�r�10�#;A � t�
`���1���96�����%C�� A�ف��J�bIncr �	����\���1o�5qni4�MNINp	xP�`���!���Hour  �� 2�21� �AAVM����0 ��T�UP ��J5�45 ��616�2�VCAM � (�CLI{O ��R6�<N2�MSC "�P �STY�L�C�28~ 13�\�NRE "FwHRM SCH^��DCSU%O�RSR {b�04� �EIOC��1 j 542 �� os| � eg�ist�����7��1�MASmK�934"7 ���OCO ��"3�8��2���� C0 HB��� 4�";39N� Re�� ��LCHK
%OP�LG%��3"%MH�CR.%MC  ; 4l? ��6 dPI�s54�s� DSW%�MD� pQ�K!63!7�0�0p"�1�Р"�4 �6<27 CgTN K � 5 ��%�"7��<25�%/�=T�%FRDM� ��Sg!��930 FB( NBA�P� ( �HLB  Men��SM$@jB( PV3C ��20v��2�HTC�CT�MIL��\@PAC� 16U�hAJ`SA�I \@ELN��<29�s�UECK <�b�@FRM �b�sOR���IPL��}Rk0CSXC ���VVFnaTg@H�TTP �!26� ��G�@ob�IGUI"%IPG�S�r� H863 �qb�!�07r�!34 |�r�84 \so`0! Qx`CC3 Fb�291�!96 rb!g51 ���!53R%� 1!s3!��~�.rp"9js VATFU�J775"��pLR6�^RP�WSMjUCTO�@xT58 F!s80���1XY ta�3!770 ��8�85�UOL  GTS�o
�{` LCM ��r| TSS�EfP6� W�\@CPE �`��0VR� l�QN�L"��@001 i7mrb�c3 =�b0�0���0�`6 w�b^-P- R-�b8n@75EW�b9 �Ґa�� ���b�`ׁ�b2 O2000��`3��`4*5�`5!�c��#$�`7.%�`8 h�605? U0�@B�6E"aRp7� !Pr8 t�a@�tr�2 iB/�1vp3L�vp5 Ȃtr9Σʐa4@-p�r3 	F��r5&�re`u�&�r7 ��r8�U�p9 \h738�a��R2D7"�1�f��2&�7� �3� 7iC��4>w58Ip�Or60 C�L��1bEN�4 I�py�L�uP��@N�-PJ8d�N�8NeN�9 H�(r`�E�b7]�|�⠂8�Вࠂ9 2H��a`0�qЂ5�%?U097 0��@q1�0���1 (�q�3 5R���0 ���mpU��0�0��7*�H@(q�\P"wRB6�q124�b`;��@���@06� 6x�3 pB/x�u ���x�6 H606�a1� ��7 6� ���p�b15�5 ����7jUU1g62 �3 g���4*�65 2ec "_��P�4U1`����B1���`0'�1�74 �q��P�E1�86 R ��P�7� ��P�8&�3 (��90 B/�s1q91����@202��6 3���A�R�U2� d��2 bI2h`��4�᪂2�L4���19v Q�2�*�u2d�Tpt2� ��EH�a2hP�$�5��F�!U2�p�p
�2�p���@5�0-@��84 @�9��TX@�� :�e5�`rb26Af�2^R�a�2Kp��1y�b5Hp�`
�5�0`@�gqGA���a52ѐ��Ḳ6�60ہ5�� ׁ2��8�E��9��EU5@ٰ\�q5�hQ`S�2ޖ5�p\�w�۲�pJ �-P��5��p1\t�H�4��PeCH�7j��phiw��@��P�x��559 ldu� P�D���Q �@������� �`.���P>��8�581l�"�q58�!AM۲�T�A iC�a58�9��@�x����5 �a��12׀0.�1����,�2����,�!P\�h8��Lp ��,�7z��6�0840\� ANRS 0C}A`��p��{��ran���FRA��Д�� ����A%���ѹ�� ������(����Ќ� ��З���������������$�G��1���⨂��������� xS�`q� � �����`64��M���iC/50T-�H������*��)p46��� C��N�����m75s֐� Sp��b46��v��༌ГM-71?�70�З����42�������C��-�а�70H�r�E��/h����O$��rD���c7c7C�q���ą���L��/��2\?imm7c7�g� ������`���(� ��e�����"��������a r��c�T,�Ѿ�"��,�� ��xx�Ex�m77t����k���5�����v)�iC��-HS -� B
_�>���+�Т�7U�]���M*h7�s��7������-9?�/260L_������QB�������]�9p�A/@���q�S��х���h6k21��c��92�������.�)92c 0�g$�@�����)$p��5$���pylH"O"
�21���t?�350����p���$�
�� �350!���0��9�U/�0\m9��M9AA3��4%� s��3M$��X%u���"him98J3����� �i d�"m4~�103�p�� ����h794̂�&R���H�0���� \���g�5AU��՜� �0���*2��00��#06�АՃ���!07{r ����� ���kЙ@����EP�#������?�p�#!�;&07\;!�B1P�߀A��/��CBׂ2�!�:/��?8�ҽCD25L�����0�"l�2BAL
#��B��\20�2 _�r�re���X��1@��N����A@��z��`C�pU��`��#04��DyA�\�`fQ��sU���\��5  ���� p�^t��<$8�5���+P=�ab1l��1LT��lA�8�!uDnE(�20�T��J�1 e�bH8�5���b�Ռ�5[�16Bs��������d�2��x��m6t !`Q����bˀ���b#�(�6iB;S�p�! ��3� ��b�s��-`�_�W8�_���&�6I	$�X5�1�Uc85��R�p6S� ���/�/+q�!�q��`񈓃6o��5m[o)�m�6sW��Q�?��set06p ��3%H�5��10p$����g�/�JrH�� � ��A�856�����F�� ���p/2��h�܅�✐)�5��̑v��(��m6��Y�H�ѝ̑�m�6�Ҝ��a6�DM�����-S�+��H 2�����Ҽ�� �r ̑��✐��l����p1���F���2�\wt6h T6H�� ��Ҝ�'Vl���� ���V7ᜐ/����;3A7��p~S��������4�`圐�V�T��!3��2�PM[�p�%ܖO�chn��vel5����Vq���_arp#��̑�.�~��2l_hemq$8�.�'�6415��� 5���?����F������5g�L�ј[���1���𙋹1����M7NU�М��eʾ����uq$D;��-�!4��3&H�f�c�Ĝ� h������u�� �㜐��ZS�!ܑ4�&��M-����S�$̑�ք �� 0��<������07shJ�H �v�À�sF��S*� ����̑���vl�3�A�T�#��QȚ�Te���q�pr����T@75j�5�dd�̑1�(UL� &�(�,���0�\�?����̑�a�� xS�t���a�e�w�2ȫ�(�	�2�C��A/����\�+p�����2�1 (ܱ�CL S ����B̺��7F��h�?�<�lơ1L� ���c� ���u9�0����e/q��O���98�K��r9 (��,��Rs�ז�5�G�m20c��i��w�A2��:�0`�$��2�2 l�0�k�X�S� ,�ι�2��O���1!4�1w���2T@� _std��G�y� �ң�<H� jdgm���� w0\� �1L���	�P��~�W*�b��t 5P������3�,����E{������LL��5\L��3��L�|#~���~!���4��#��O����h�L6 A�������2璥���44�����[6\j4s��·��@�#��ol�E"w�8P k�����?0xj�H1�1`Rr�>��]�2a�#2Aw�P ��2��|41�8��ˡ��{� �%�A<��� +�?�l��0`�&�"��|�`Am1�2@��ػ��3�HqB ��K�R��ˑb�W� ��Fs���)�ѐ�!����a�1����5��16�16C��C<����0\imBQ���d����b��\B5�-���DiL���O�_�<ѠPEtL�E�RH��ZǠPgω�am1l ��u���̑�b�<����<�$�T�̑�F�����Ȋ�Dpb��X"x�ᒢ��p� ����^t��9�0\� �j971\kckrcfJ�F�s������c��e "CTM�E�r�����!�a�`main.[��g�`Grun}�_vc�# 0�w�1Oܕ_u����bctme��Ӧ�`�ܑ�j735�-� KAREL U�se {�U���J���1���p� U ̑�9�B@��L�9����7j[�atk208 "K��Kя��\��9��a��̹�����cKRC�a�o ��kc�qJ�&s��� ��Grſ�fsD��:y�0�s��A1X\j|хr�dtB�, ��`.	v�q�� �sǑIf��Wfj52�TKQu�to Set��J�� H5K536�(�932���91�5�8(�9�BA�1(�7�4O,A$�(TCP Ak���/�)Y�� �\tpqtool.v��v���! conre;a�#�Controlw Re�ble��CNRE(�T�<�4��2���D�)���S�55i2��q(g�� (����4X�cOux�\s�futs�UTS `�i�栜���t�棈���? 6�T�!�S#A OO+D6����������,!��6�c+� igt�t6iB��I0�TW8 �0��la��vo58�o�b@Få򬡯i�Xh���!Xk�0Y!8\m6e�!6EC���v��6���������<1!6�A���A�6s��ƀ�U�g�T|ώ���rE1�qR��˔Z4�T������,#�eZp)g ����<ONO0���uJ���tCR;��F�a� �xSt�f��prdsuchk �1���2&&?���t��*D %$�r(�✑�娟:r���'�s�qO��<s�crc�C�\At�trldJ"o�\�V�|���Paylo�nfirm�l�!�87��7��A�3ad�! �?ވI�?hplQ��3��3"�q��x pl�`���d87��l�calC�u�Du���;��movx�����initX�:s8O��a�r4 ���r67A4|�e GeneratiڲĐ��7g2q$��g =R� (Sh��c ,|�bE��$ԒA\�:�"��4���4�4�. sg��5��F$d6"e�!p? "SHAP�T�Q ngcr pGC��a(�&"� ��"G3DA¶��r6�"�aW�/�$dataxX:s�"tpad��<[q�%tput;a__�O7;a�o8�1�yl+s��r�?�:�#�?�5x$�?�:c O�:y O�:H�IO�s`O%g�q�ǒ�?�@0\��"o�j�92;!�Ppl.C�ollis�QSkip#��@5��@J��D ��@\ވ�C@X��7��7�|s2��potcls�LS��DU�k?�\_ et1s�`�< \�Q䜐�@���`dcKqQ�F�C;��J,�n��` (��4eN����T�{���'j(�c�q����/IӸaȁ��̠GH�����зa��e\mcclmt "CLM�/��� �mate\��lmpALM�?>p7qCmc?����2vm�qp��%�3s��_sv90<�_x_msu�2L�^v_� K�o�{in��8(3r<�c_lo�gr��rtrcW� �v_3�~yac��d�<�ten��der$cCe�' Fiρ�R��Q��?�l�enteAr߄|��(Sd��V1�TX�+fK�r�a�99sQ9+�5�r�\tq\� "FN�DR���S�TDn$LAN]G�Pgui��D�`���S������sp�!ğ֙uf�ҝ�s����$�����e+�=�� �������������w�H�r\fn_�ϣ��|$`x�tcpma��- TCP�����?R638 R�Ҭ���38��M7p, ���Ӡ�$Ӡ�8p0Р��VS,�>�tk��99 �a��B3���PզԠ��0D�2�����UI��t� ��hqB���8��������p���re�ȿ��exe@4φ�B���pe38�ԡG�rmpWXφ�var@�φ�@3N�����vx�!ҡ���q�RBT �$cOPTN ask E0��1��R MAS0�H5�93/�96 H5�0�i�480�5�H0��m�Q�K��7�0�g�Pl�h0ԧ�2�ORDP��@"��_t\mas��0�a@��"�ԧ�����k�� �R����ӹ`m��bL��7�.f��u�d���r��splay�D�E���1w�UPD�T Ub��887 M(��Di{���v�� ��Ԛ⧔��#�B���|����o  ��� �a�䣣��60q��B�����qscan0��B���ad@�������q`�䗣��#��К�`2�� vl v��Ù�$�>�b����! S��Easyy/К�Util��|룙�511 J������R7 ��Nor|֠��inc),<6Q�� �`c��"4�[���986FVRx� So����q�nd 6����P��4�a\ (�@�
  �������d���K�bdZ���men�7���- Me`t!yFњ�Fb�0�T�Ua�577?i 3R��\�5�u?��!� n���f���<���l\mh�Ц�pűE|hmn�	���<\O���eD�1�� l!��y��Ù�\|p����B���Ћmh�@��:. aG!���/�t��55�6�!X�l�.u�s��Y/k)ensu)bL���eK�h��  �B\1;5g?y?�?�?D��?*rm�p�?Ktbox O2K|?0�G��C?A%ds���?1ӛ#� �TR��/� �P�4B�`�U�P�V�P"�Q�P0�U�PO��P�"�T3�U�P�f�Pk"�2}�4�T�P�f�P2�"�Q5�S�Q���R?�Ă�Q3t.�P׀al���P+OP51�7��IN0a��Q(8}g��PESTf3u�a�PB�l�ig�h�6��aq��P � sxS��`  n��0mbumpP�Q969g�69�Qq��P�0�baAp�@Q� �BOX��,>vchqe�s�>vetu㒼�=wffse�3� ��]�;u`aW��:z#ol�sm<ub�a-��]D�K�ibQ�c���p�Q<twaǂ tp�Q�҄Taror ROecov�b�O�P�642����a�0q��a⁠QErǃ�QCry�з`�P'�T�`��aar������	{'�p�ak971��71���m���>�pjo@t��PXc��C�1�adb� -�ail��na�g���b�QR629��a�Q��b�P  ?�
  �P���$$CL[q O����������$�PS_DI�GIT���"�!�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����*�璬1:PROD�UCT�Q0\PGSTK�bV,n��99�\����$FEAT_I�NDEX��~��� 搠I�LECOMP ;��)��"���SETUP2 �<��� � N !�_AP2BCK 1=�?  �)}6/"E+%,/i/��W/ �/~+/�/O/�/s/�/ ?�/>?�/b?t??�? '?�?�?]?�?�?O(O �?LO�?pO�?}O�O5O �OYO�O _�O$_�OH_ Z_�O~__�_�_C_�_ g_�_�_	o2o�_Vo�_ zo�oo�o?o�o�ouo 
�o.@�od�o� ��M�q�� �<��`�r����%� ��̏[�������!� J�ُn�������3�ȟ W������"���F�X� �|����/���֯e� �����0���T��x� �����=�ҿ�s�π��,ϻ�9�b�� P�/ 2) *.cVRiϳ�!�*�����������PC��7�!�FR6:D"�c��χ��T� �߽�Lը��ܮx���*.F��>� �	N�,�k��ߏ��STM �����Q������!�iPe�ndant Pa'nel���H��F����4������GIF�������u����JPG&P��<�����	PAN?EL1.DT�́������2 �Y�G��
3w�����//�
4�a/�O///��/�
TPEIN�S.XML�/����\�/�/�!Cus�tom Tool�bar?�PA?SSWORD/�?FRS:\R??� %Passw�ord Config�?��?k?�?O H�6O�?ZOlO�?�OO �O�OUO�OyO_�O�O D_�Oh_�Oa_�_-_�_ Q_�_�_�_o�_@oRo �_voo�o)o;o�o_o �o�o�o*�oN�or ��7��m� �&���\����� y���E�ڏi������ 4�ÏX�j�������� A�S��w�����B� џf�������+���O� ��������>�ͯ߯ t����'���ο]�� ���(Ϸ�L�ۿpς� Ϧ�5���Y�k� ߏ� $߳��Z���~�ߢ� ��C���g�����2� ��V����ߌ���?� ����u�
���.�@��� d������)���M��� q�����<��5r �%��[� &�J�n� �3�W���"/ �F/X/�|//�/�/ A/�/e/�/�/�/0?�/ T?�/M?�??�?=?�? �?s?O�?,O>O�?bO �?�OO'O�OKO�OoO �O_�O:_�O^_p_�O �_#_�_�_Y_�_}_o�_�_Ho)f�$FI�LE_DGBCK� 1=��5`��� (� �)
SUMM?ARY.DGRo�\OMD:�o�o
`�Diag Su�mmary�o�Z
CONSLOG�o��o�a
J�aCo�nsole lo�gK�[�`MEMCHECK@'�o��^qMemor?y Data��W߁)�qHADOW���P��s�Shadow ChangesS��-c-��)	F�TP=��9����w�`qmment T�BD׏�W0<�)�ETHERNE�T̏�^�q�Z��a�Ethernet� bpfigura�tion[��P��DCSVRFˏ��Ï�ܟ�q%�� v�erify alylߟ-c1PY���DIFFԟ��̟a���p%��dif!fc���q��1X�?�Q�� ����{X��CHGD��¯ԯi��px��� �¤�2`�G�Y�� 1��� �GD��ʿ�ܿq��p���Ϥ�F�Y3h�O�a��� 1��(�GD���ψ��y��p�ϡ�0��UPDATES.��Ц��[FRS:�\�����aUpd�ates Lis�t���kPSRBW�LD.CM.��\���B��_pPS_R?OBOWEL���_ ����o��,o!�3��� W���{�
�t���@��� d�����/��Se �����N�r � =�a�r �&�J���/ �9/K/�o/��/"/ �/�/X/�/|/�/#?�/ G?�/k?}??�?0?�? �?f?�?�?O�?OUO �?yOO�O�O>O�ObO �O	_�O-_�OQ_c_�O �__�_:_�_�_p_o �_o;o�__o�_�o�o $o�oHo�o�o~o�o 7�o0m�o� � �V�z�!��E� �i�{�
���.�ÏR� ���������.�S�� w������<�џ`��� ���+���O�ޟH��� ���8���߯n����$FILE_��{PR��������� ��MDONLY 1�=4�� 
 ���w�į��诨�ѿ �������+Ϻ�O�޿ sυ�ϩ�8�����n� ߒ�'߶�4�]��ρ� ߥ߷�F���j���� ��5���Y�k��ߏ�� ��B�����x����1� C���g������,��� P���������?���Lu�VISBC�KR�<�a�*.V�D|�4 FR:�\��4 Vi�sion VD file� :L bpZ�#��Y �}/$/�H/�l/ �/�/1/�/�/�/�/ �/ ?�/1?V?�/z?	? �?�???�?c?�?�?�? .O�?ROdOO�OO�O ;O�O�OqO_�O*_<_ �O`_�O�__%_�_��MR_GRP 1�>4�L�UC4�  B�P	 �]�ol`�*u����RHB� ��2 ���� ��� ��� He�Y�Q`orkbIh�o�Jd�o�Sc�o�oK��C{LXkJ��F�5U�a�R��+�o�o �E|�D����DU�?-i��
8�k=�u�c}?�\$?��))lr$��?��xq0~�� F�@ �r�d�a}J���NJk�H�9�Hu��F!��IP�sX~��`�.9�<9��896�C'6<,6�\b�}A���A�MB����B�OA�#��B�� �+~��A|�BYK��Amy�A�7A�����,.��PA�����|�ݏx����%���p�A6Β@U��{ �v�a�������П�� ��ߟ��<�'�hz;BH�P �a`�<Q��QA>�K����ï�T
6�P=��PI�`˯�o�o�B��P5���@�3�3@���4�m�,�@�UUU��U�~w�>u.�?!x��^��ֿ���3��=�[z�=�̽=�V6<�=�=�=$q��~���@8�i7�G��8�D�8@9!�7���@Ϣ���cD�@ D�� Cϫof��C��Po�C'� 6��_V� m�o��To�� xo�ߜo������A� ,�e�P�b����� ��������=�(�a� L���p���������.� ������*��N9r ]������� �8#\nY� }�������/ ԭ//A/�e/P/�/p/ �/�/�/�/�/?�/+? ?;?a?L?�?p?�?�? �?�?�?�?�?'OOKO 6OoO�OHߢOl��ߐ� ���O�� _��G_bOk_ V_�_z_�_�_�_�_�_ o�_1ooUo@oyodo vo�o�o�o�o�o�o Nu�� �������;� &�_�J���n������� ݏȏ��%�7�I�[� "/�描�����ٟ�� �����3��W�B�{� f�������կ����� ��A�,�e�P�b��� �����O�O�O��O �OL�_p�:_������ ���������'��7� ]�H߁�lߥߐ��ߴ� ������#��G�2�k� 2��Vw�������� ���1��U�@�R��� v������������� -Q�u��� r��6��) M4q\n��� ���/�#/I/4/ m/X/�/|/�/�/�/�/ �/?ֿ�B?�f?0� BϜ?f��?���/�?�? �?/OOSO>OwObO�O �O�O�O�O�O�O__ =_(_a_L_^_�_�_�_ ���_��o�_o9o$o ]oHo�olo�o�o�o�o �o�o�o#G2k V{�h���� ���C�.�g�y�`� ���������Џ�� �?�*�c�N���r��� �����̟��)�� M�_�&?H?���?���? �?�?����?@�I�4� m�X�j�����ǿ��� ֿ����E�0�i�T� ��xϱϜ�������� �_,��_S���w�b߇� �ߘ��߼������� =�(�:�s�^���� �������'�9� � ]�o����~������� ������5 YD V�z����� �1U@yd ��v�����/Я */��
/�u/��/�/ �/�/�/�/�/??;? &?_?J?�?n?�?�?�? �?�?O�?%OOIO4O "�|OBO�O>O�O�O�O �O�O!__E_0_i_T_ �_x_�_�_�_�_�_o �_/o��?oeowo�oP� �oo�o�o�o�o+ =$aL�p�� �����'��K� 6�o�Z������ɏ�� 폴� ��D�/ / z�D/��h/ş���ԟ ���1��U�@�R��� v�����ӯ������ -��Q�<�u�`���`O �O�O���޿��;� &�_�J�oϕπϹϤ� �������%��"�[� F��Fo�ߵ����ߠo ��d�!���W�>�{� b������������ ��A�,�>�w�b��� �������������=��$FNO ����\��
F0�l q  FLAG�>�(RRM_C�HKTYP  r] ��d �] ���OM� _MI�N� 	���� ��  XT SSB_CFG ?\ �����OTP�_DEF_OW � 	��,IR�COM� >�$G�ENOVRD_D�O��<�lTH�R� d�dq_�ENB] qR�AVC_GRP s1@�I X( / %/7//[/B// �/x/�/�/�/�/�/? �/3??C?i?P?�?t? �?�?�?�?�?OOO�AO(OeOLO^O�OoR�OU�F\� ��,�B,�8�?���O�O�O	_|_���  DE_��Hy_�\@@m_B��=�vR/��I�O�SMT�G�SUoo|&oRHOSTC�s1H�I� ���zMSM�l[�bo�	127�.0�`1�o  e�o�o�o#z�o�FXj|�l60s	�anonymou�s������Qao�&�&��o �x��o������ҏ� 3��,�>�a�O�� ��������Ο�U%�7� I��]����f�x��� �����ү����+� i�{�P�b�t������ ������S�(�:� L�^ϭ�oϔϦϸ��� ���=��$�6�H�Z� ����Ϳs�������� ��� �2���V�h�z� ��߰���������
� �k�}ߏߡߣ���� ����������C�* <Nq�_���� ��-�?�Q�c�eJ ��n����� ��/"/E�X/j/ |/�/�/�%'/ ?[0?B?T?f?x?� �?�?�?�?�??E/W/�,O>OPObO�KDaEN�T 1I�K P�!�?�O  �P �O�O�O�O�O#_�OG_ 
_S_._|_�_d_�_�_ �_�_o�_1o�_ogo *o�oNo�oro�o�o�o 	�o-�oQu8 n������� �#��L�q�4���X� ��|�ݏ���ď֏7����[���B�QUICC0��h�z�۟���1ܟ��ʟ+���2�,���{�!ROUTER|�X�j�˯!PCJOG̯���!192.�168.0.10���}GNAME �!�J!ROBO�T�vNS_CFG� 1H�I ��Auto-started�$/FTP�/���/ �?޿#?��&�8�J� �?nπϒϤ�ǿ��[� �����"�4ߵ&���� ������濜������� ���'�9�K�]�o�� �����������/ �/�/G���k��ߏ��� ����������1 T���Py���� �"�4�	H-|�Q cu�VD��� �/�;/M/_/q/ �/����/
/�/> ?%?7?I?[?*/?�? �?�?�/�?l?�?O!O 3OEO�/�/�/�/�?�O  ?�O�O�O__�?A_ S_e_w_�O4_._�_�_ �_�_oVOhOzO�O�_ so�O�o�o�o�o�o�_ '9Kno�o� ����o*o<oNo P5��oY�k�}����� pŏ׏����0����C�U�g�y���_�T_?ERR J;������PDUSIZ � ��^P�����>ٕWRD ?�z���  ?guest����+�=�O�a�s�*�SC�DMNGRP 2�Kz�Ð���۠\��K�� �	P01.14� 8�q   �y��B  _  ;����{� �����������������������~� �ǟI�4�m�X�|���  i  ��  
����� ����+��������
����l�.x����"B�l�ڲ۰s�d��������_GROuU��L�� ���	��۠07K�QU�PD  ����PČ�TYg������TTP_AUT�H 1M�� <�!iPenda�n���<�_�!�KAREL:*8�����KC%�5��G��VISION SETZ���|��Ҽߪ������ ���
�W�.�@��d��v���CTRL �N�������
�FFF9E3����FRS:DE�FAULT��FANUC We�b Server�
������q��������������WR_�CONFIG �O�� ���I�DL_CPU_P5C"��B��= w�BH#MIN.��BGNR_IO಑� ���% NPT_SIM_DOs�}TPMODN�TOLs �_P�RTY�=!OL_NK 1P��� '9K]o�MASTEr ���>��O_CFG���UO����CYC�LE���_AS�G 1Q���
 q2/D/V/h/z/�/ �/�/�/�/�/�/
??\y"NUM���<Q�IPCH�����RTRY_CN�"�u���SCRN(������ ����R����?���$J23_DSP_EN�����0?OBPROC�3�n�JOGV�1S_��@��8�?��';ZO'??0CPOS�REO�KANJI_�Ϡu�A#��3�T ���E�O�EC�L_LM B2e?�@EYLOGGIN��������LANGUAGE _��=� }Q��LeG�2U����� ��x�����PC �V �'0������MC:\RSC�H\00\˝LN�_DISP V��������TOC��4Dz\A�SO�GBOOK W�+��o���o�o���Xi�o�o�o�o�o~b}	x(y��	ne�i�ekElG_B�UFF 1X���}2����Ӣ� �����'�T�K� ]�����������ɏۏ����#�P��ËqD�CS Zxm =���%|d1h`����ʟܟ�g�IO 1[+ �?'����'�7�I�[�o���� ����ǯٯ����!� 3�G�W�i�{��������ÿ׿�El TM  ��d��#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y�p�ߝ߈t�SEV�0�m�TYP��� ��$�}�ARS�"�(_�s�2FL 1\��0����������������5�TP�<P���DmNG�NAM�4�U�f�UPS`GI�5�A�5}s�_LOAD@oG %j%@�_MOV�u����MAXUALRMB7��P8��y���3�0(]&q��Ca]s�3��~�� 8@=@^+k طv	��V0�+�P�A5d�r���U���� ��E(iT y������� / /A/,/Q/w/b/�/ ~/�/�/�/�/�/?? )?O?:?s?V?�?�?�? �?�?�?�?O'OOKO .OoOZOlO�O�O�O�O �O�O�O#__G_2_D_ }_`_�_�_�_�_�_�_ �_o
ooUo8oyodo �o�o�o�o�o�o�o�o�-��D_LDXD�ISA^�� �ME�MO_APX�E {?��
 � 0y�����������ISC 1_�� �O���� W�i�����Ə��� ��}��ߏD�/�h�z� a������������ ��@���O�a�5��� ���������u��ׯ <�'�`�r�Y������ y�޿�ۿ���8Ϲ� G�Y�-ϒ�}϶ϝ��� ��m�����4��X�j��#�_MSTR �`��}�SCD 1as}�R���N����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{?�?�?�?n�MKCF/G b���?�ҿLTARM_�2c�RuB ��3WpTNBpMETP�UOp�2����N�DSP_CMNT�nE@F�E�� d���N�2A�O�D�E_POSCF�G�N�PSTOL 1e�-�4@�<#�
 ;Q�1;UK_YW7_Y_[_ m_�_�_�_�_�_�_o �_oQo3oEo�oio{o��o�a�ASING_?CHK  �MAq/ODAQ2CfO�7�J�eDEV 	�Rz	MC:'|HOSIZEn@����eTASK %<z�%$123456�789 ��u�gT�RIG 1g�� l<u%���3�0��>svvYPaq���kEM_INF �1h9G �`)AT&F�V0E0(���)���E0V1&A3�&B1&D2&S0&C1S0=��)ATZ���ڄ�H������G�ֈA�O�w�2�������џ  ��������͏ߏP�� t�������]�ί��� ��(�۟�^��#� 5�����k�ܿ� ϻ� ů6��Z�A�~ϐ�C� ��g�y��������2� i�C�h�ό�G߰��� ���ߙϫ�������� d�v�)ߚ��߾�y�� ������<�N��r� %�7�I�[������ 9�&��J[�g���>ONITOR�@G ?;{   �	EXEC1T�3�2�3�4�Q5��p�7�8�9�3�n�R�R �RRRR (R4R@RLRU2Y2e2q2}U2�2�2�2�U2�2�3Y3e�3��aR_GRP?_SV 1it��q�(�a?�ڿ{
��5��۵MO~q_DCd~�1�PL_NAME �!<u� �!�Default �Personal�ity (fro�m FD) �4R�R2k! 1j)T?EX)TH��!�AX d�?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O�Ox2-?�O�O�O_�_0_B_T_f_x_�b< �O�_�_�_�_�_�_o@ o2oDoVoho&xRj"g 1o�)&0\�bO, �9��b�a� @D�  �a?���c�a?�`�a�aA�'�6�ew;��	l�b	 �xJp���`�`	p �<� �(p� ��.r� K�K ���K=*�J����J���JV���kq`q�P��x�|5p@j�@wT;f�r�f�qx�acrs�I�� ��p���p�r� h}��3��´  ��>��ph�`z��꜖"g�Jm�q� H��N��ac���dw�� � �  P� Q� �� |  �а�m�Əi}	'�� � �I�� �  �����:�È���=���(�ts�a�	���I  �n @H�i~�ab��Ӌ�b�w��urN<0��  'Ж�q��p@2��@�����r�q5�C�pC>0C�@ C��z��`
�A1�q   @�B�V~X�
nwBD0h�A��p�ӊ�p�`���aDz���֏࿯�Я	�pv�(� �� -���I��-�=��A�a���e_q�`�p �??�ff ��m�|�� �����Ƽuq@ݿ�>1�  P�apv(�`ţ�� �=�qst��?˙��`x`�5p<
�6b<߈;����<�ê<�? <�&P�ς��AO��c1��ƍ�?offf?O�?&���qt@�.�J<?�`��wi4� ���dly�e߾g;ߪ� t��p�[ߔ�߸ߣ� ���� ����6�wh�F0%�r�!�����1ى����E��� E�O�G+� F�!���/���?�e�`P���t���lyBL�cB��Enw4������� +��R��s���������h�yÔ�>���I�mXj���A�y�weC��������#/*/c/�N/wi�����v/C�`� CHs/`
=$��p�<!�!��ܼ�'��3A�A�AR�1AO�^?��$�?��5p���
=ç>�����3�W
=�s#�]�;e�׬a�@����{�����<�>�(�B�u���=B0�������	R��zH��F�G���G���H�U`E����C�+��}I�#�I��H�D�F��E��RC�j=�>�
I��@H��!H�( E?<YD0w/O *OONO9OrO]O�O�O �O�O�O�O�O_�O8_ #_\_G_�_�_}_�_�_ �_�_�_�_"oooXo Co|ogo�o�o�o�o�o �o�o	B-fQ �u������ �,��P�b�M���q� ����Ώ���ݏ�(� �L�7�p�[������ ʟ���ٟ���6�!��Z�E�W���#1($1�3�9�K���ĥ%�����ƯS�3ǭ8���S�4M�gs��,�IB+�8�J��a���{�d�d�����ȿ��(�ڼ%P8�P�=:GϚ�S�6�h�z���R�Ϯ�������,���  %�� �� h�Vߌ�z߰�&�g�/ 9�$�������7�����A�S�e�w�  ������������~�2 F�$�&'Gb������,��!C���@����8�����F� D�zN�� F�P D�������)#B�'9K]o#�?���@@v
J$�8�8��8�.
 v�� �!3EWi{�����:� ���ۨ�1��$�MSKCFMAP�  ��� ���(.��ONREL  ��!9��EX_CFENBE'
#�7%^!FNCe/W$JOGOVLIME'�dO S"d�KEY�E'�%�RUN�,�%�SFSPDTY0g&P%9#�SIGNE/W$T1�MOT�/T!�_�CE_GRP 1-p��#\x��? p��?�?�?�?�?O �?OBO�?fOO[O�O SO�O�O�O�O�O_,_ �OP__I_�_=_�_�_ �_�_�_oo�_:o��TCOM_CF/G 1q	-�vo�o�o
Va_ARC�_b"�p)UAP�_CPL�ot$NO�CHECK ?	+ �x� %7I[m�� ������!�.+�NO_WAIT_�L 7%S2NT^a�r	+�s�_ER�R_12s	)9�� A,ȍޏ��x��x�&��dT_MO��}t��, �*o|q�9�PARAM��u	+��a�ß�'g{�� =?�345678901� �,��K�]�9�i��������ɯۯ��&g������C��cUM_?RSPACE/��|����$ODRD�SP�c#6p(OFF�SET_CART��o��DISƿ��PEN_FILE��!�ai��`OPTI�ON_IO�/��PWORK ve7s# ��V�ؤ����<�p�4�p�	 ���p��<�� C��_DSBL  Đ�P#��ϸ�RI_ENTTOD ?��C�� !l�UT�_SIM_D$��"���V��LCT w}�h�iĜa[�>1�_PEXE�j�RATvШ&p%� ���2^3j)TEX)�TH�)�X d3�������%�7� I�[�m������� �������!�3�E���2��u����������� ����c�<d�A Sew���������Ǎ�^0OU�a0o(��(�����u2, ���O H @D7�  [?�aG1?��cc�D][<�Z�;�	ls���xJƵ�������_< ���s���ڐH(��H3�k7HSM5G��22G���Gpc
͜�'f�/,-,ڐCR�>�D!��M#{Z/��3�����4y H "��c/u/�/0B_�����jc��t3�!�/ �/�"�t32����/6 W ��P%�Q%��%�|T��S62�q?�'e	'� � ��2I� � � ��+==�̡ͳ?�;	�h	�0��I  �n �@�2�.��Ov;���ٟ?&gN�]O  �''�uD@!� C�C��@F#H!�/�O�O Nsb
���@�@E��@�e0@B��QA�0Yv: �13Uwz$oV_�/z_�e_�_�_	��( �� -�2@�1�1ta�Ua�c����:A����.  �?�ff���[o"o�_!U�`oX�0A8���o:�j>�1  Po�V(���eF0�f�Y����L�?����x�b0@<
6b<�߈;܍�<��ê<� <�#&�,/aA�;r��@Ov0P?fff?��0?&ip�T@�.�{r�J<?�`�u#	�Bdqt�Yc �a�Mw�Bo�� 7�"�[�F��j����� ��ُ����3�����,���(�E��� E��3G+� F��a��ҟ������,��P�;���B�pAZ�>��B��6�<O ίD���P��t�=����a�s�����6j�h�y�7o��>�S���O�����Fϑ�A�a�_��C3Ϙ�/�<%?��?������(���#	Ę��P �N�||CH���Ŀx������@I�_��'�3A�A�A�R1AO�^??�$�?������±
=ç>�����3�W
=�#� U��e����B��@��{�����<����(�B�u���=B0�������	�b�H��F�G���G���H�U`E����C�+��I�#�I��H�D�F��E��RC�j=[��
I��@H��!H�( E?<YD0߻� �������� �9�$� ]�H�Z���~������� ������#5 YD }h������ �
C.gR� ������	/� -//*/c/N/�/r/�/ �/�/�/�/?�/)?? M?8?q?\?�?�?�?�? �?�?�?O�?7O"O[O mOXO�O|O�O�O�O�O��O�O�O3_Q(���3���b��gUU���W_i_2�3ǭ8��_�_2�4M�gs�_�_�RIB+��_�_�a���{�miGo5okoYo(�o}l��P'rP�nܡݯ�o=_�o�_�[R?Q�u�,��  �p���o ��/��S��z
uү ܠ�������ڱ������������  /�M�w�e�������~�l2 F�$��'Gb��t��a�`�,p�S�C�y�@p�5��G�Y�۠F� D�z�� F�P D��]����پ��ʯܯ� ��~ÿ?���@@�J?�K�K���K���
 �|��� ����Ŀֿ������0�B�T�fϽ�V� ����{��1��$�PARAM_ME�NU ?3���  �DEFPULS�Er�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L��	�OPT���PTB4�.�C��R_DECSN ���e��ߑߣ����� ������!�3�\�W��i�{���USE_PROG %��q%�����CCR����e����_HOSoT !��!��:���T�`�V��/��X����_TIMqE��^��  ��?GDEBUG\�����GINP_FL'MSK����Tfp�����PGA  ��̹�)CH����TY+PE������� ����� - ?hcu���� ���//@/;/M/ _/�/�/�/�/�/�/�/��/??%?7?`?��W�ORD ?	=�	RSfu	P�NSUԜ2JO�K�DRTEy�]T�RACECTL �1x3��� }�`� &�`��`�>�6DT Q�y3�%@�0D �� �c��a:@V�@BR�2ODOVOhOzO�O�O �O�O�O�O�O
__.Z<TDT,Sb_t_@�_�Z]_�SM �R._T@_RXN\L�
o �["cP_�_�VJ�PbF�T�WJ`Nd	Nd
NdNdNd5of@oRo dovo�o�o�o�o�o�o (:L^p�����r�t^��r*�t�t�t�Yb� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�.Iv����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t������� ��������(: L^p��j��� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o��o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*���$PGTRACELEN  )��  ���(��>�_UP �z���m��u�Y�n�>�_C�FG {m�W�(�n���PЬ�� ��DEFSPD� |��'�P���>�IN��TRLW }��(�8���IPE_CONF�I��~m���mњ��Ԛ�>�L�ID����=�G�RP 1��W���)�A ����&ff(�A+33�D�� D]� ?CÀ A@1����(�d�Ԭ��0�0�?� 	 1��1��� ´�����B�9����O�9��s�(�>�T?��
5�������� =��=#�
�� ��P;t_��������  #Dz (�
H �X~i���� ��/�/D///h/�S/�/��
V7.10beta1���  A�E}�"ӻ�A (��� ?!G��!>˙��"����!̽��!BQ��!AA\� �!���!2p����Ț/8?J?\?n?B};� ���/��/ �?}/�?�?OO:O%O 7OpO[O�OO�O�O�O �O�O_�O6_!_Z_E_ ~_i_�_�_�_�_�_�_ 'o2o�_VoAoSo�o wo�o�o�o�o�o�o .R=v1�/�#F@ �y�}��{ m��y=��1�'�O� a��?�?�?������ߏ ʏ��'��K�6�H� ��l�����ɟ���؟ �#��G�2�k�V��� z��������o�� ίC�.�g�R�d����� �����п	���-�?� *�cώ���Ϯ�� ����B�;�f�x� ������DϹ��߶��� �����7�"�[�F�X� ��|����������� !�3��W�B�{�f��� ������ �����/ S>wbt�� ����=O zόϾψ����ϼ � /.�'/R�d�v߈� �/0�/�/�/�/�/�/ �/#??G?2?k?V?h? �?�?�?�?�?�?O�? 1OCO.OgORO�OvO�O �O���O�O�O__?_ *_c_N_�_r_�_�_�_ �_�_o�_)oTfx �to���/�o/ >/P/b/t/mo �|������ �3��W�B�{�f�x� ����Տ������� A�S�>�w�b����O�� џ������+��O� :�s�^�������ͯ�� �ܯ�@oRodo�o`� �o�o�o��ƿ�o��� *<N�Y��}�h� �ό��ϰ�������� 
�C�.�g�Rߋ�v߈� �߬�����	���-�� Q�c�N�ﲟ���l� �������;�&�_� J���n����������� ,�>�P�:L���� ��������(� :�3��0iT�x �����/�// /S/>/w/b/�/�/�/ �/�/�/�/??=?(? a?s?��?�?X?�?�? �?�?O'OOKO6OoO ZO�O~O�O�O�O�O *\&_8_r���_��_��$PLID�_KNOW_M � ��� Q�TSV �v��P��?o"o4o�OXoCo�Uo�o R�SM_G�RP 1��Z'0*{`�@�`uf�e�`
�5� �gpk 'Pe]o �����������SMR�c��mT�EyQ}? yR���� ������폯���ӏ� G�!��-��������� ��韫���ϟ�C�� �)������������ا���QST�a1 �1��)���P0� A 4��E2� D�V�h�������߿¿ Կ���9��.�o�R� d�vψ��ϬϾ�����2�0� Q�<3��3�/�A�S��A4l�~ߐߢ��5���������6
��.�@��7Y�k�}����8��������MA/D  )���PARNUM � !�}o+��S+CHE� S�
��f�8���S��UPDf�x���_CMPa_�`H�� �'�U~ER_CHK-����ZE*<RqSr��_�Q_MOG���_�X�_RES_G��!���D� >1bU�y �����/�	/����+/�k� H/g/l/��Ї/�/�/ �	��/�/�/�X�? $?)?���D?c?h?�����?�?�?�V 1�U�ax�@c]��@t@(@c\��@�@D@c[��*@��THR_ICNRr�J�b�Ud2FoMASS?O ZSG�MN>OqCMON_�QUEUE ���U�V P~P X�N�$ UhN�FV�@E�ND�A��IEXE�O�E��BE�@�O�COPTIO�G��@�PROGRAM %�J%�@�?��~�BTASK_IG��6^OCFG ��Oz��_�PDATA��c��[@Ц2 =�DoVohozo�j2o�o �o�o�o�o);�M jINFO[��m��D���� ����1�C�U�g� y���������ӏ���h	�dwpt�l )��QE DIT ���_i��^WERFL�X	C�RGADJ7 �tZA������?נʕFA��IOR�ITY�GW���M�PDSPNQ����U�GD��OTOE�@1�X� (!AF:@E� c�Ч?!tcpn����!ud����!�icm���?<�X�Y_�Q�X���Q)� *�1�5��P��]�@�L��� p��������ʿ�+�=�$�a�Hυϗ�*���PORT)QH���P�E��_CARTREPPX�ПSKSTA�H�
S�SAV�@�tZ	�2500H863����_x�
�'��X�
@�swPtS�ߕ߼����URGE�@Bl��x	WF��DO�F�"[W\�������W�RUP_DELA�Y �X���R_'HOTqX	B%�c����R_NORMA�Lq^R��v�SEM�I�����9�QSKkIP'��tUr�x 	7�1�1��X� j�|�?�tU�������� ������$J\ n4������ ��4FX| j������� /0/B//R/x/f/�/��/�/tU�$RCV�TM$��D�� DkCR'���Ў!�A���Bz�C9˫?�<�W\:�.��:���C���'����5���n:�o?�� <�
6b<߈;�܍�>u.�?!<�&�? h?�?�?�@>��?O O 2ODOVOhOzO�O�O�O �O�O�?�O�O__@_ +_=_v_Y_�_�_�?�_ �_�_oo*o<oNo`o ro�o�o�o�_�o�o�o �o�o8J-n� �_������� "�4�F�X�j�U���� ��ď���ӏ��� B�T��x��������� ҟ�����,�>�)� b�M������������ ïկ�Y�:�L�^�p� ��������ʿܿ� � ���6�!�Z�E�~ϐ� {ϴϗ�����-�� � 2�D�V�h�zߌߞ߰� ��������
���.�� R�=�v��k���� ������*�<�N�`� r�������������� ��&J\?� ������� "4FXj|��!�GN_ATC 1��	; AT&FV0E0��ATDP/6�/9/2/9��ATA�,�AT%G1%B9�60�+++��,�H/,�!I�O_TYPE  ��%�#t�RE�FPOS1 1�>V+ x�u/�n�/j�/
=�/�/ �/Q?<?u??�?4?�?�X?�?�?�+2 1�V+�/�?�?\O�?�O<�?�!3 1�O*O�<OvO�O�O_�OS4 1��O�O�O_�_�t_�_+_S5 1� B_T_f_�_o	oBo�_S6 1��_�_�_�5o�o�o�oUoS7 1�lo~o�o�oH3|l�oS8 1��%_���SMASK 1�V/�  
?�M��XN	OS/�r������!?MOTE  n��$���_CFG ���q���"PL_R�ANG�����PO�WER ������SM_DRY�PRG %o�%��P��TART ���^�UME_�PRO-�?����$_�EXEC_ENB�  ���GSP�D��Րݘ��TD�B��
�RM�
�MKT_'�T�����OBOT_NAM/E o�����OB_ORD_N_UM ?�b!�H863 � �կ����PC_TIME�OUT�� x�S�232Ă1��� LTEAC�H PENDAN��w��-���Mainten�ance Con�s���s�"���KCL/Cm��

��t�ҿ No Use-�����0�NPO�򁋁���.�CH�_L������q	���s�MAVAI�L�����糅��S�PACE1 2��, j�߂�DɈ�s�߂� �{S�8�?�k�v�k� Z߬��ߤ��ߚ� � 2�D���hߊ�|��`� ��������� � 2�D��h��|���`�@��������y���2����0�B���f��� ��{���3);M_� �����/� /44FXj|*/ ���/�/�/?(??=?5Q/c/u/�/�/ G?�/�/�?O�?$OEO,OZO6n?�?�?�? �?dO�?�?_,_�OA_b_I_w_7�O�O�O �O�O�_�O_(oIoo ^oofo�o8�_�_ �_�_�_�oo6oEf�){���G ;�o� ���
M� ���*� <�N�`�r�������w����o�収���d .��%�S�e�w����� ������Ǐَ���Θ 8�+�=�k�}������� ůׯ͟����%�'� X�K�]���������ӿ ������#�E�W�w `� @��������x�����\� e�����������R� d߂�8�j߬߾߈ߒ� �����������0�r� ���X�������� ����8����
�ύ��_MODE  y�{��S ��{|�2�0������3�	S|)CW�ORK_AD���7��+R  ��{�`� �� _I�NTVAL���d����R_OPTIO�N� ��H V�AT_GRP 2ݭ�up(N�k|� �_�����/ 0/B/��h�u/T� }/ �/�/�/�/�/�/?!? �/E?W?i?{?�?�?5? �?�?�?�?�?O/OAO OeOwO�O�O�O�OUO �O�O__�O=_O_a_ s_5_�_�_�_�_�_�_ �_o'o9o�_Iooo�o �oUo�o�o�o�o�o �o5GYk-�� �u�����1� C��g�y���M����� ӏ叧�	��-�?�Q� c������������� ��ǟ�;�M�_�����$SCAN_T�IM��_%}�R� �(�#((��<04�d d 
! D�ʣ��u�/������U��2H5���@�d5�P�g��]	����������dd�x�  P����� ��  �8� ҿ�!���D��$�M�_�qσϕ� �Ϲ��������ƿv��F�X��</� ;�ob���pm��t��_DiQ̡  � l�|�̡ĥ�� �����!�3�E�W�i� {������������ ��/�A�S�e�]�� �������������� );M_q�� �����r� ��j�Tfx��� ����//,/>/ P/b/t/�/�/�/�/�/�%�/  0��6�� !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O*�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo�O�O J�o�o�o�o�o�o�o  2DVhz� ������
�7?  ;�>�P�b�t� ��������Ǐُ��� �!�3�E�W�i�{���8����ß �ş3� ܟ��&�8�J�\�n� �����������ɯ�����,� ��+�	1234�5678�� 	� =5���f�x������������� 
��.�@�R�d�vψ� ��៾��������� *�<�N�`�r߄߳Ϩ� ����������&�8� J�\�n�ߒ����� �������"�4�F�u� j�|������������� ��0_�Tfx ������� I>Pbt�� �����!/(/ :/L/^/p/�/�/�/�/�/�/�2�/?�#�/9?K?]?�iCz�  Bp˚   ���h2��*�$�SCR_GRP �1�(�U8(ӿ\xd��@ � ��'�	 �3�1�2�4 (1*�&�I3�F1OO�XO}m��D�@�0ʛ)���HUK�L�M-10iAo 890?�90;���F;�M61C �D�:�CP��1
\&V�1	�6F��CW�9)A7Y	(R�_�_�_h�_�_�\���0 i^�oOUO>oPo#G �/���o'o�o�o�o.�oB�0�r�tAA�0*  @�Bu&Xw?��ju�b�H0{UzAF@ F�`�r��o� ����+��O�:� s��mBqrr����������B�͏b����7� "�[�F�X���|����� ٟğ���N���AO�0�B�CU
L���E�jq�Bq>g�#H@��@pϯ B����G�I
E�0EL_D�EFAULT  ��T���E��MIPOWERFL  
Ex*��7�WFDO�� *��1ERVE�NT 1����`(�� L!D?UM_EIP��>���j!AF_I�NE�¿C�!FIT������!o�:� ��a�!�RPC_MAIN�b�DȺPϭ�t�VI�S}�Cɻ����!�TP��PU�ϫ�d���E�!
PMON?_PROXYF߮�Ae4ߑ��_ߧ�f�����!RDM_S�RV�߫�g��)�!#R�Iﰴh�u�K!
v�M�ߨ�id����!RLSYN�C��>�8���!�ROS��4��4 ��Y�(�}���J�\��� ����������7�� ["4F�j|� ���!�Ei�o�ICE_KL �?%� (%SVCPRG1n >���3��3��"�4//�5./3/"�6V/[/�7~/�/���D�/�9�/�+ �@��/��#?�� K?��s?� /�?� H/�?�p/�?��/O ��/;O��/cO�? �O�9?�O�a?�O� �?_��?+_��?S_ �O{_�)O�_�QO �_�yO�_��Os� ���>o�o}1�o�o �o�o�o�o�o; M8q\���� �����7�"�[� F��j�������ُď ���!��E�0�W�{� f�����ß���ҟ� ��A�,�e�P���t���������ί�y_�DEV ���MC:��_!�OUT���2��REC 1q�`e�j� �	 �����˿��p�ڿ��
 �`e ���6�N�<�r�`ϖ� �Ϧ��Ϯ�������&� �J�8�n߀�bߤߒ� �߶�������"��2� X�F�|�j������� ��������.�T�B� x�Z�l����������� ��,P>`b t������ (L:\�d� ���� /�$/6/ /Z/H/~/l/�/�/�/ �/.��/?�/2? ?V? D?f?�?n?�?�?�?�? �?
O�?.O@O"OdORO �OvO�O�O�O�O�O�O __<_*_`_N_�_�_ x_�_�_�_�_�_oo 8oo,ono\o�o�o�o �o�o�o�o�o " 4jX����� �����B�$�f� T�v������������ ؏��>�,�b�P�r����p�V 1�}� �P
�	!��^�� ����TYP�E\��HELL_?CFG �.�F��  	�����RSR������ӯ �������?�*�<� u�`�����������~��  ��%�3�E��Q�\�bҰM�o�p��d���2Ұd]�K�:�H�K 1�H�  u�������A�<�N� `߉߄ߖߨ������߀����&�8��=�OMM �H���9��FTOV_ENB�&�1�OW_RE�G_UI���IM/WAIT��a���OUT������T�IM�����V�AL����_UNI�T��K�1�MON_�ALIAS ?e~w� ( he�# ����������Ҵ�� );M��q��� �d��%� I[m�<�� ����!/3/E/W/ /{/�/�/�/�/n/�/ �/??/?�/S?e?w? �?�?F?�?�?�?�?�? O+O=OOOaOO�O�O �O�O�OxO�O__'_ 9_�O]_o_�_�_>_�_ �_�_�_�_�_#o5oGo Yokoo�o�o�o�o�o �o�o1C�og y��H���� 	��-�?�Q�c�u� � ������ϏᏌ��� )�;��L�q������� R�˟ݟ�����7� I�[�m��*�����ǯ ٯ믖��!�3�E�� i�{�������\�տ� ����ȿA�S�e�w� ��4ϭϿ����ώ��� �+�=�O���s߅ߗ� �߻�f�������'� ��K�]�o���>�� ��������#�5�G� Y��}���������n���$SMON_D�EFPRO ������� *SYS�TEM*  d=���RECALL� ?}�� ( ��}2copy �frs:orde�rfil.dat� virt:\t�mpback\=�>inspiron:992��q��n�}).mdb:*.*CU	X����
-x.:\ �8R�m��e..a6H2 ] � //�-?Qb/ t/�/�/�F/��/�/ ??)�M�/p?�? �?�8?J?]?�? OO��%
xyzrate 61 �?�?�?�nO�O�O�%.GR(1844 HOZO�O�O_�(3./@/�Ma_s_�_�_� *�/I_�DY_ �_�_o�?3?FO�C�_no�o�o�%/�??o�I ^o�o&O8O�o�o�m��O�J620 �OX��� 2t����n�������I5512G�Y����� !_3_�_��a�s����� �_E���Y�����!o 3oFݟn������o 6�H�Z�_����'� 9�]�n��������� ɟ[�����#�5�ȯ Y�j�|ώϡ���D�ׯ ������1���U�f� xߊߝ���J�ӿ���� ��-���Q�b�t�� ���<��Ϛ����� )������p������� ��D�V������0�@����ew�����A10E I[��#�4.�@߸bt�� }+��I� Z��/��4�G�� �o/�/�/&�0��?/ �
_/�/??'9� �n?�?�?��/�[?��?�?O#��$SN�PX_ASG 1߸���9A�� P 0 �'%R[1�]@1.1O �?�#�%dO�OsO�O�O �O�O�O�O __D_'_ 9_z_]_�_�_�_�_�_ �_
o�_o@o#odoGo Yo�o}o�o�o�o�o�o �o*4`C�g y������� 	�J�-�T���c����� ��ڏ�����4�� )�j�M�t�����ğ�� ����ݟ�0��T�7� I���m��������ǯ ٯ���$�P�3�t�W� i��������ÿ�� ��:��D�p�Sϔ�w� ���ϭ��� ���$�� �Z�=�dߐ�sߴߗ� �������� ��D�'� 9�z�]������� ��
����@�#�d�G� Y���}����������� ��*4`C�g y������ 	J-T�c�� ����/�4// )/j/M/t/�/�/�/�/��/�/�/?0?4,DPARAM �9E�CA �	���:P�4�0$HO�FT_KB_CF�G  p3?E�4P�IN_SIM  9K�6�?�?�?�0�,@RVQSTP_DSB�>�21On8�J0SR ��;�� & MULT�IROBOTTA�SK=Op3�6T�OP_ON_ER�R  �F�8�AP_TN �5�@�A�BRIN�G_PRM�O �J0VDT_GRP� 1�Y9�@  	�7n8_(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o  2Dkhz�� �����
�1�.� @�R�d�v��������� Џ�����*�<�N� `�r���������̟ޟ ���&�8�J�\��� ��������ȯگ��� �"�I�F�X�j�|��� ����Ŀֿ���� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�tߛߘߪ߼��� ������(�:�a�^� p�����������  �'�$�6�H�Z�l�~���������������3V�PRG_COUN�T�6��A�5ENB�OM=�4J_UPD 1��;8  
p2� ����� )$ 6Hql~��� ��/�/ /I/D/ V/h/�/�/�/�/�/�/ �/�/!??.?@?i?d? v?�?�?�?�?�?�?�? OOAO<ONO`O�O�O �O�O�O�O�O�O__ &_8_a_\_n_�_�_�_�YSDEBUG�" � �Pdk	�PS�P_PASS"�B?�[LOG ���m�P��X�_  �g�Q
MC:\d�_b_MPCm��o�o��Qa�o �vfS_AV �m:dlUb�U\gSV�\�TEM_TIMEw 1�� (�P孳T��o	T1S�VGUNS} #'�k�spASK_?OPTION" ��gospBCCF�G ��| 8�b�{�}`��� �a&��#�\�G���k� ����ȏ������"� �F�1�j�U���y��� ğ���ӟ���0��T�f��UR���S��� ƯA������ ��D� �nd��t9�l������� ��ڿȿ�����"� X�F�|�jϠώ��ϲ� ��������B�0�f� T�v�xߊ��ߦؑ��� ����(��L�:�\� ��p���������� � �6�$�F�H�Z��� ~������������� 2 VDzh�� �������4 Fdv���� ��//*/�N/</ r/`/�/�/�/�/�/�/ �/??8?&?\?J?l? �?�?�?�?�?�?�?�? OO"OXOFO|O2�O �O�O�O�OfO_�O_ B_0_f_x_�_X_�_�_ �_�_�_�_oooPo >otobo�o�o�o�o�o �o�o:(^L np�����O� �$�6�H��l�Z�|� ����Ə؏ꏸ���� 2� �V�D�f�h�z��� ��ԟ����
�,� R�@�v�d��������� ίЯ���<��T� f�������&�̿��ܿ ��&�8�J��n�\� �π϶Ϥ�������� ��4�"�X�F�|�jߌ� �ߠ����������� .�0�B�x�f��R��� ���������,��<� b�P�������x����� ����&(:p ^�������  6$ZH~l ��������/ &/D/V/h/��/z/�/��/�/�/�&0�$T�BCSG_GRP� 2��%��  �1 
? ?�  /?A? +?e?O?�?s?�?�?�?��?�;23�<d�, �$A?1	� HC���6>�@E�5CL  �B�'2^OjH4Jݸ�B\)LFY g A�jO�MB��?F�IBl�O�O�@�JG|_�@�  D	�15_ __$YC-P{_F_$`_j\��_�]@0�> �X�Uo�_�_6oSoo�0o~o�o�k�h�0	V3.00'2�	m61c�c	�*�`�d2�o�e>əJC0(�a�i �,p�m-  �0�����omvu1JC�FG ��%� 1 #0vz��rrBrv�x�� ��z� �%��I�4� m�X���|�������� ֏���3��W�B�g� ��x�����՟����� ���S�>�w�b��� ��'2A ��ʯܯ��� ���E�0�i�T���x� ��ÿտ翢����/� �?�e�1�/���/�� �Ϯ��������,�� P�>�`߆�tߪߘ��� ���������L�:� p�^��������� ��� �6�H�>/`�r� ���������������  0Vhz8� �����
. �R@vd��� ����//</*/ L/r/`/�/�/�/�/�/ �/�/�/?8?&?\?J? �?n?�?�?�?�?���? OO�?FO4OVOXOjO �O�O�O�O�O�O__ �OB_0_f_T_v_�_�_ �_z_�_�_�_oo>o ,oboPoroto�o�o�o �o�o�o(8^ L�p����� ��$��H�6�l�~� (O����f�d��؏� ��2� �B�D�V����� ��n����ԟ
���.� @�R�d����v����� ���Я���*��N� <�^�`�r�����̿�� �޿��$�J�8�n� \ϒπ϶Ϥ������� ߊ�(�:�L���|�j� �߲ߠ���������� 0�B�T��x�f��� �����������,�� P�>�t�b��������� ������:(J L^������  �6$ZH~ l��^���dߚ  //D/2/h/V/x/�/ �/�/�/�/�/�/?
? @?.?d?v?�?�?T?�? �?�?�?�?OO<O*O `ONO�OrO�O�O�O�O �O_�O&__6_8_J_ �_n_�_�_�_�_�_�_ �_"ooFo��po�o ,oZo�o�o�o�o�o 0Tfx�H� ������,�>� �b�P���t������� ��Ώ��(��L�:� p�^�������ʟ��� ܟ� �"�$�6�l�Z� ��~�����دꯔo� �&�ЯV�D�z�h��� ����Կ¿��
��.π�R�@�v�dϚτ� s ���� ��������$TBJO�P_GRP 2����� O ?������������x/JBЌ��9�� �< �zX���� @����	 �C�� >t�b  C����>��͘Րդ��>̚йѳ33=��CLj�ff�f?��?�ffB@G��ь�����t�ц��>�(�\)��ߖ�E噙�;���hCYj��  �@h��B�  A�����f��C� � Dhъ�1���O�4�N����
�:���Bl^���j�i�l�l����A�ϙ�A�"��D��֊=qH������p�h�Q�;��A�j�ٙ7�@L��D	2��������$�6�>B�\p��T���Q�tsx�@33@���C����y�1����>G��Dh�������<���<{�h�@i� ��t� �	���K&� j�n|���p��/�/:/k/�ԇ����!��	V3�.00J�m61cI�*� IԿ��/��' Eo��E��E���E�F���F!�F8���FT�Fqe\�F�NaF����F�^lF����F�:
F�)�F��3G��G��G���G,I�!CH`��C�dTDU��?D��D���DE(!/E\��E��E�h��E�ME���sF`F+'�\FD��F`�=F}'�F���F�[
F����F��M;��;WQ�T,8�4` *Q�ϴ?�2���3�\�X/O��ESTP?ARS  ��	����HR@ABLE� 1����0��D
H�7 8��9
G
H�
H����
G	
H
�
H
HYE��
H�
H
H6FRDIAO�XOjO|O�O�O�ETO"_4[>_P_b_Ht_�^:BS _� �J GoYoko}o�o�o�o�o �o�o�o1CU gy����`#oRL �y�_�_�_�_�O�O�O��O�OX:B�rNUM�  ����P��� V@P:B_?CFG ˭�Z��h�@��IMEBF_TT%AU��2@�GVERS�q���R 1���
 (I�/����b� �� ��J�\���j�|���ǟ ��ȟ֟�����0� B�T���x�������2��_���@�
��M�I_CHAN�� �� ��DBGLV����������ET�HERAD ?*��O�������xh�����ROUT�!��!������?SNMASKD��>U�255.���#������OOLOF/S_DI%@�u.��ORQCTRL �����}ϛ3rϧ� ����������%�7� I�[�:���h�z߯�A�PE_DETAI�"�G�PON_SV�OFF=���P_M�ON �֍�2���STRTCHK� �^�����VTCOMPAT���O�����FPROG� %^�%MU�LTIROBOT�Tݱ���9�PLA�Y&H��_INST+_Mް �������US�q��LCK����QUICKM�E�=���SCRE�Z�G�tps� ���u�z�����_��@@n�.�SR_�GRP 1�^�/ �O���� 
��+O=sa�쀚�
m���� ��L/C1g U�y����� 	/�-//Q/?/a/�/�	123456�7�0�/�/@Xt�1����
 �}i�pnl/� gen.htm�? ?2?�D?V?`Pan�el setupZ<}P�?�?�?�?�?�? �??,O>OPO bOtO�O�?�O!O�O�O �O__(_�O�O^_p_ �_�_�_�_/_]_S_ o o$o6oHoZo�_~o�_ �o�o�o�o�o�oso�o 2DVhz�1 '���
��.�� R��v���������Џ|G���UALRM��oG ?9� � 1�#�5�f�Y���}��� ����џן���,���P��SEV  �����ECFG ��롽�}A��   BȽ�
 Q���^���� 	��-�?�Q�c�u���Й��������� P�����I��?����(%D�6� �$�]� Hρ�lϥϐ��ϴ��π����#��G���� ��߿U�I_Y�H�IST 1�� � (�� ���3/SOFTP�ART/GENL�INK?curr�ent=edit�page,��,1����!�3��� �����menu��962�߆����K�]�o�36u�
��.� @���W�i�{������� ��R�����/A ��ew����N ��+=O��s�������� f��f//'/9/K/ ]/`�/�/�/�/�/�/ j/�/?#?5?G?Y?�/ �/�?�?�?�?�?�?x? OO1OCOUOgO�?�O �O�O�O�O�OtO�O_ -_?_Q_c_u__�_�_ �_�_�_�_��)o;o Mo_oqo�o�_�o�o�o �o�o�o%7I[ m� ���� ���3�E�W�i�{� �����ÏՏ���� ���A�S�e�w����� *���џ�����o oO�a�s��������� ͯ߯���'���K� ]�o���������F�ۿ ����#�5�ĿY�k� }Ϗϡϳ�B������� ��1�C���g�yߋ� �߯���P�����	�� -�?�*�<�u���� ����������)�;� M�������������� ��l�%7I[ �������h z!3EWi� ������v/�///A/S/e/P����$UI_PANE�DATA 1������!?  	�}w/�/`�/�/�/?? )? >?��/i?{?�?�?�? �?*?�?�?OOOAO (OeOLO�O�O�O�O�O��O�O�O_&Y� b�>RQ?V_h_z_�_ �_�__�_G?�_
oo .o@oRodo�_�ooo�o �o�o�o�o�o*< #`G��}�-\�v�#�_��!�3� E�W��{��_����Ï Տ���`��/��S� :�w���p�����џ�� ����+��O�a�� �������ͯ߯�D� ���9�K�]�o����� ���ɿ���Կ�#� 
�G�.�k�}�dϡψ� ���Ͼ���n���1�C� U�g�yߋ��ϯ���4� ����	��-�?��c� J���������� �����;�M�4�q�X� ���������� %7��[���� ���@��3 WiP�t�� ���/�//A/�� ��w/�/�/�/�/�/$/ �/h?+?=?O?a?s? �?�/�?�?�?�?�?O �?'OOKO]ODO�OhO �O�O�O�ON/`/_#_ 5_G_Y_k_�O�_�_? �_�_�_�_oo�_Co *ogoyo`o�o�o�o�o �o�o�o-Q8u�O�O}��������)�>��U -�j�|�������ď+� �Ϗ���B�)�f� M���������������ݟ�&�S�K�$U�I_PANELI�NK 1�U�  � � ��}1234567890s� ��������ͯդ�Rq� ���!�3�E�W��{��������ÿտm�m�h&����Qo�  � 0�B�T�f�x��v�&� ����������ߤ�0� B�T�f�xߊ�"ߘ��� �������߲�>�P� b�t���0������ ������$�L�^�p� ����,�>������� $�0,&�[g I�m����� ��>P3t� i��Ϻ� -n� �'/9/K/]/o/�/t� /�/�/�/�/�/?�/ )?;?M?_?q?�?�U Q�=�2"��?�?�?O O%O7O��OOaOsO�O �O�O�OJO�O�O__ '_9_�O]_o_�_�_�_ �_F_�_�_�_o#o5o Go�_ko}o�o�o�o�o To�o�o1C�o gy�����B �	��-��Q�c�F� ����|�������֏ �)��M���=�?� �?/ȟڟ����"� ?F�X�j�|�����/� į֯�����0��? �?�?x���������ҿ Y����,�>�P�b� �ϘϪϼ�����o� ��(�:�L�^��ς� �ߦ߸�������}�� $�6�H�Z�l��ߐ�� ��������y�� �2� D�V�h�z����-��� ������
��.R dG��}��� �c���<��`r ��������/ /&/8/J/�n/�/�/ �/�/�/7�I�[�	�"? 4?F?X?j?|?��?�? �?�?�?�?�?O0OBO TOfOxO�OO�O�O�O �O�O_�O,_>_P_b_ t_�__�_�_�_�_�_ oo�_:oLo^opo�o �o#o�o�o�o�o  ��6H�l~a� �������2� �V�h�K������� 1�U
��.�@�R� d�W/��������П� �����*�<�N�`�r� �/�/?��̯ޯ�� �&���J�\�n����� ��3�ȿڿ����"� ��F�X�j�|ώϠϲ� A���������0߿� T�f�xߊߜ߮�=��� ������,�>���b� t�����+���� �����:�L�/�p��� e����������� ���6���ۏ���$UI_QUICKMEN  ���}���RESTORE �1٩�  �
�8m3\n�� �G����/� 4/F/X/j/|/'�/�/ �//�/�/??0?�/ T?f?x?�?�?�?Q?�? �?�?OO�/'O9OKO �?�O�O�O�O�OqO�O __(_:_�O^_p_�_ �_�_QO[_�_�_I_�_ $o6oHoZoloo�o�o �o�o�o{o�o 2 D�_Qcu�o�� �����.�@�R� d�v��������Џ�ޜSCRE� ?��u1sc�� u2�3�4��5�6�7�8<��USER���2�T���ks'���U4��5��6��7���8��� NDO_C�FG ڱ  ��  � PDAT�E h���None�SEU�FRAME  �ϖ��RTOL_ABRT�����ENB(��GRP� 1��	�Cz  A�~�|�%|� ������į֦���X�� UH�X�7�MS�K  K�S�7�N&�%uT�%������VISCAND�_MAXI�I��3���FAIL_ISMGI�z �% #S����IMREGNU�MI�
���SIZlI�� �ϔ,�?ONTMOU'�K��Ε�&����a��a��s��FR:\�� �� MC:�\(�\LOGh�B@Ԕ !{��Ϡ������z �MCV����UDM1 �EX	�z >��PO64_�Q���n6��PO�!�LI�Oڞ�e�V��N�f@`�I��w =	_�SZVm�w���`�WAIm����STAT ݄k�% @��4�F�T�$�#�x �2DWP�  ��P G<��=��͎����_JMPER�R 1ޱ
  ��p2345678901���	�:� -�?�]�c������������������$�ML�OW�ޘ�����_T�I/�˘'��MPHASE  k��ԓ� ��SHIF�T%�1 Ǚ��<z��_�� ��F/|Se �������0/ //?/x/O/a/�/�/��/�/�/����k�	�VSFT1\�	�V��M+3 �5��Ք p����Aȯ  B8[0[0�"Πpg3a1Y2�_3Y�F7ME��K�͗	6\e���&%��M��i�b��	��$��TDINEND3�4��4OH�+�G1�O�S2OIV I���]LRELEvI��4�.�@��1_ACTI�V�IT��B��A ��m��/_��BRD�BГOZ�YBOX c�ǝf_\��b��2�TI19o0.0.�P83p\;�V254p^�Ԓ	 �S�_�[�b��rob�ot84q_   �p�9o\�pc�PZoMh�]Hm�_�Jk@1�o�ZABC
d��k�,���P\�Xo }�o0);M� q�������H�>��aZ�b��_V