��   ?3�A��*SYST�EM*��V7.5�0122 8/�1/2   A �  ���M�N_MCR_TA�BLE   �� $MACRO�_NAME �%$PROG@E�PT_INDEX�  $OPE�N_IDaASSIGN_TYPD � qk$MO�N_NO}PRE�V_SUBy a �$USER_WO�RK���_L� M�S�DUMMY1�0  &S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VIRTUA�L�/�!;LDUI�MT  �������$MAOXDRI� ��5��%.1 �%� � d%�Open han�d 1����% ta?�? �"  �!��# �%Clo�seQ?d?�?�?�9>�7Relax�?�?H)OOO�9�6L82QO 2O�OVO�3 �?�O�O
_�O�4O�O�Ol__�6�Fh_�_d_�_�[�3���_o�_:o �_�_poomo�oUogo �o�o �o�o6H3 l-�Q�u� ���2���h�� ��;�M���ԏ������ ��.�ݏR�d��%��� I���m�������*� ٟ�`����3�E��� ̯��𯟯��&�կJ� ���E���A���e�w� 쿛�Ͽ�ѿ�X�� |�+�=ϲ�a����ϗ� �����B����x�'� u߮�]�o��ߓ��� ��>�P�;�t�#�5�� Y���}�������:� ����p����C�U��� ���� ����6��Z l-�Q�u� ���2��h �;M����� �./�R///M/�/ I/�/m//�/�/?�/ �/?`??�?3?E?�? i?�?�?�?�?&O�?JO �?O�O/O}O�OeOwO �O�O_�O�OF_X_C_ |_+_=_�_a_�_�_�_ �_o�_Bo�_oxo'o �oKo]o�o�o�o�o �o>�obt#5� Y�}����:� ��p����C�U�ʏ ܏Ǐ �����6��Z� 	��U���Q�Ɵu��� ���� �ϟ��h�� ��;�M�¯q������ ��.�ݯR�����7� ����m�������ǿ ٿN�`�Kτ�3�EϺ� i��ύϟ���&���J� ��߀�/ߤ�S�eߟ� �ߛ�����F���j� |�+�=��a����� ���	�B����x�'� ��K�]��������� ��>��b#]� Y�}��(� �#p�CU� y� /��6/�Z/ 	//�/?/�/�/u/�/ �/�/ ?�/�/V?h?S? �?;?M?�?q?�?�?�? �?.O�?ROOO�O7O �O[OmO�O�O�O_�O �ON_�Or_�_3_E_�_ i_�_�_�_o�_oJo �_o�o/o�oSoeo�o �o�o�o�oF�oj +e�a��� ��0���+�x�'� ��K�]�ҏ������� ɏ>��b��#���G� ��Ο}������(�ן �^�p�[���C�U�ʯ y�����6��Z� 	����?���c�u��� ���� �Ͽ�V��z� ��;�M���q��ϕϧ������R���
S�end Even�tU�5�SEND�EVNT��3��i��%	}�Da�ta�ߘ�DATA��߿���%}�S�ysVar��S�YSVY��1�%�Get��Z�G�ET����%�Request �Menu����RE�QMENU!��� ��?߀�;ߤ�_���� ��������F��j +�O���� �0��fxc �K]����� �>/�b//#/�/G/ �/k/}/�/?�/(?�/ �/^??�?�?C?U?�? y?�?�?�?$O�?!OZO 	OO�O?O�OcOuO�O �O�O _�O�OV__z_ )_;_u_�_q_�_�_�_ o�_@o�_o;o�o7o �o[omo�o�o�o �oN�or!3�W ������8�� �n���k���S�e�ڏ ����������F���j� �+���O�ğs����� ���0�ߟ�f���� ��K�]�ү�������� ,�ۯ)�b��#���G� ��k�}����(�׿ �^�ς�1�C�}��� y��ϝϯ�$���H��π	�Cߐ�?ߴ�c�u���$MACRO_M�AX:���  ����Ж��S�OPENBL �����՗��r�r�A���PDIgMSK�����Y�SUc�u�TPDSBEX  -�
q�U����n��� �