��   I�A��*SYST�EM*��V7.5�0130 3/�19/2015 A 
  ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��ETH_FLT�R.� $� �  �FT�P_CTRL.� @ $LOG�_8	�CMO>�$DNLD_FI�LTE� � SUB�DIRCAP��� HO��NT.� 4� H_NAM�E !AD�DRTYPA H_LENGTH'� �z +LS� D $R�OBOTIG P�EER^� MAS�KMRU~OM�GDEV#� R�DM*�DIS�ABL&� T�CPIG/ 3 $ARPSIZ&�_IPF'W_�MC��F_IN�� FA~LASS�s�HO_� IN{FO��TELKG PV�b�	 WORD  �$ACCESS�_LVL?TIM�EOUTuORT� � �ICEUS�= � �$#  ����!�� �� � VIRTUA�L�/�!'0 �%W
���F����ظ�"�%����+ �����$Ȱ� �-2%;�SHARED 1�)?  P!�!�?���!|?�?�?�?�? O�?%O�?1OOZOO BO�OfO�O�O�O�O_ �O�OE__i_,_�_P_ �_t_�_�_�_o�_/o �_SooLo�oxo�opo �o�o�o�o�o*O s6�Z�~� ����9��]� � ��D�V���z�ۏ���� #���Y�H�}�@����)7z _LIST� 1=x!1E.ܒ0��d�ە1�>d�255.$��&����%ړ2��@X���+�=�O�3Y���Р�������O�4 ѯ�H���	��-�O�5I����o�������O�6���8������ �$���-�  ���-�!�%�%��&!�Ò�)�0H!�� ���rj3O_tpd���! � >�!!KC� e��0ٙ��&W�!C�m ��w߉�S�!GCON� ��1�=�Osmon��W�